`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module local_controller_prefetch_module(clk, reset, init, controller_id, write_flag, glob_controller_sending, from_glob_controller_prefetch_start_addr, from_glob_controller_prefetch_stop_addr,  prefetch_data_from_sram, input_boundary_flag, prev_prefetch_dest_address, from_glob_prefetch_dest_addr, prefetch_packet_out, boundary_prev, prefetch_dest_address, scenario_end_flag, coeff_num, from_glob_prefetch_reqd);
    // parameter
    parameter N_row = 1024;
	parameter datawidth = 32;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for subscaled system
	parameter id_width = 11; // 1221 local controllers in subscaled system
	parameter row_address_width = 10; /// assuming 1024 rows and 64 columns: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	
	
	
        
    // input
    input clk; // system clock, generated by VCO
	input reset;
	input init;
	input glob_controller_sending; //not used
	input [2*datawidth - 1:0] prefetch_data_from_sram;
	input [id_width - 1:0] controller_id;
	input input_boundary_flag;
	input write_flag;
	input [address_vector_width - 1:0] prev__prefetch_dest_address;
	input [address_vector_width - 1:0] from_glob_prefetch_dest_addr;
	input [row_address_width - 1:0] from_glob_controller_prefetch_start_addr;
	input [row_address_width - 1:0] from_glob_controller_prefetch_stop_addr;
	input scenario_end_flag;
	input coeff_num;
	input from_glob_prefetch_reqd;

    // output
    output [packet_width-1:0] prefetch_packet_out; 
    output reg boundary_prev;
    output reg [address_vector_width - 1:0] prefetch_dest_address;
	
	

    // internal status regs/signals
    reg [row_address_width-1:0] prefetch_row_address;
	reg [id_width - 1:0] id; 
	reg [packet_width-1:0] prefetch_packet_out_internal;
	reg prefetch_reqd;
	reg [row_address_width-1:0] prefetch_stop_address;
    

    // logic part  
    assign prefetch_packet_out = prefetch_packet_out_internal;

	//sequential logic
    always @ (posedge clk) begin
        if (reset) begin
			prefetch_row_address <= 0;
			prefetch_packet_out_internal <= 264'bz;
			prefetch_dest_address <= 0;
			
        end
        else if (init) begin
			prefetch_packet_out_internal <= 264'bz;
			
			if (from_glob_prefetch_dest_addr[0] == 1'b1 || from_glob_prefetch_dest_addr[0] == 1'b0) begin
				prefetch_row_address <= from_glob_controller_prefetch_start_addr;
				prefetch_stop_address <= frm_glob_controller_prefetch_stop_addr;
				prefetch_dest_address <= from_glob_prefetch_dest_addr;
				prefetch_reqd <= 1;
			end
			
			else begin
				prefetch_row_address <= prefetch_row_address;
				prefetch_stop_address <= prefetch_stop_address;
				prefetch_dest_address <= prefetch_dest_addr;
				prefetch_reqd <= prefetch_reqd;

			end
			
        end
		else begin
			if (coeff_num == 0 && write_flag == 0 && prefetch_reqd == 1) begin
				prefetch_packet_out_internal <= {data_from_sram, prefetch_dest_address};
				prefetch_row_address <= prefetch_row_address + 1;
				
			end
			else if (coeff_num == 1 || write_flag == 1 || prefetch_reqd == 0) begin
				packet_out_internal <= {264'bz};
				prefetch_row_address <= prefetch_row_address;		
			end
			prefetch_dest_address <= prefetch_dest_address;
			prefetch_stop_sddress <= prefetch_stop_address;
			prefetch_dest_address <= prefetch_dest_address;
		end  
     end
	 
	 always @ (posedge clk) begin
		if (prefetch_row_address == N_row - 1) begin
			boundary_prev <= 1;
		end
		else begin
			boundary_prev <= 0;
		end
	 end
	 
	 
	 always @ (negedge clk) begin
		boundary_prev <= 0;
		if (reset) begin
			prefetch_row_address <= prefetch_row_address;
			prefetch_dest_address <= prefetch_dest_address;
		end
		else if (input_boundary_flag == 1) begin
			row_address <= N_row - 1;
			prefetch_dest_address <= prev_dest_address;
		end
		else if (input_boundary_flag == 0) begin
			if (boundary_next == 1) begin
				coeff_num <= 0;
			end
			else begin
				coeff_num <= coeff_num;
			end
			row_address <= row_address;
			dest_address <= dest_address;
			
		end
	 end
	 
	 


   
endmodule
    
