
module crossbar_one_hot_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [31:0] i_valid;
  input [1023:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [255:0] i_cmd;
  input clk, rst, i_en;
  wire   N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210,
         N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220,
         N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230,
         N1231, N1232, N1233, N1234, N1422, N1423, N1424, N1425, N1426, N1427,
         N1428, N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437,
         N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447,
         N1448, N1449, N1450, N1451, N1452, N1453, N1454, N1642, N1643, N1644,
         N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654,
         N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664,
         N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674,
         N1862, N1863, N1864, N1865, N1866, N1867, N1868, N1869, N1870, N1871,
         N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881,
         N1882, N1883, N1884, N1885, N1886, N1887, N1888, N1889, N1890, N1891,
         N1892, N1893, N1894, N2082, N2083, N2084, N2085, N2086, N2087, N2088,
         N2089, N2090, N2091, N2092, N2093, N2094, N2095, N2096, N2097, N2098,
         N2099, N2100, N2101, N2102, N2103, N2104, N2105, N2106, N2107, N2108,
         N2109, N2110, N2111, N2112, N2113, N2114, N2228, N2229, N2230, N2231,
         N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239, N2240, N2241,
         N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251,
         N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259, N2260, N2316,
         N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326,
         N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336,
         N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346,
         N2347, N2348, N2404, N2405, N2406, N2407, N2408, N2409, N2410, N2411,
         N2412, N2413, N2414, N2415, N2416, N2417, N2418, N2419, N2420, N2421,
         N2422, N2423, N2424, N2425, N2426, N2427, N2428, N2429, N2430, N2431,
         N2432, N2433, N2434, N2435, N2436, N2492, N2493, N2494, N2495, N2496,
         N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504, N2505, N2506,
         N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514, N2515, N2516,
         N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2580, N2581,
         N2582, N2583, N2584, N2585, N2586, N2587, N2588, N2589, N2590, N2591,
         N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, N2601,
         N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611,
         N2612, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676,
         N2677, N2678, N2679, N2680, N2681, N2682, N2683, N2684, N2685, N2686,
         N2687, N2688, N2689, N2690, N2691, N2692, N2693, N2694, N2695, N2696,
         N2697, N2698, N2699, N2700, N2756, N2757, N2758, N2759, N2760, N2761,
         N2762, N2763, N2764, N2765, N2766, N2767, N2768, N2769, N2770, N2771,
         N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2779, N2780, N2781,
         N2782, N2783, N2784, N2785, N2786, N2787, N2788, N2844, N2845, N2846,
         N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2856,
         N2857, N2858, N2859, N2860, N2861, N2862, N2863, N2864, N2865, N2866,
         N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876,
         N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941,
         N2942, N2943, N2944, N2945, N2946, N2947, N2948, N2949, N2950, N2951,
         N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961,
         N2962, N2963, N2964, N3078, N3079, N3080, N3081, N3082, N3083, N3084,
         N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094,
         N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104,
         N3105, N3106, N3107, N3108, N3109, N3110, N3294, N3295, N3296, N3297,
         N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307,
         N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317,
         N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3510,
         N3511, N3512, N3513, N3514, N3515, N3516, N3517, N3518, N3519, N3520,
         N3521, N3522, N3523, N3524, N3525, N3526, N3527, N3528, N3529, N3530,
         N3531, N3532, N3533, N3534, N3535, N3536, N3537, N3538, N3539, N3540,
         N3541, N3542, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3733,
         N3734, N3735, N3736, N3737, N3738, N3739, N3740, N3741, N3742, N3743,
         N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753,
         N3754, N3755, N3756, N3757, N3758, N3942, N3943, N3944, N3945, N3946,
         N3947, N3948, N3949, N3950, N3951, N3952, N3953, N3954, N3955, N3956,
         N3957, N3958, N3959, N3960, N3961, N3962, N3963, N3964, N3965, N3966,
         N3967, N3968, N3969, N3970, N3971, N3972, N3973, N3974, N4158, N4159,
         N4160, N4161, N4162, N4163, N4164, N4165, N4166, N4167, N4168, N4169,
         N4170, N4171, N4172, N4173, N4174, N4175, N4176, N4177, N4178, N4179,
         N4180, N4181, N4182, N4183, N4184, N4185, N4186, N4187, N4188, N4189,
         N4190, N4374, N4375, N4376, N4377, N4378, N4379, N4380, N4381, N4382,
         N4383, N4384, N4385, N4386, N4387, N4388, N4389, N4390, N4391, N4392,
         N4393, N4394, N4395, N4396, N4397, N4398, N4399, N4400, N4401, N4402,
         N4403, N4404, N4405, N4406, N4590, N4591, N4592, N4593, N4594, N4595,
         N4596, N4597, N4598, N4599, N4600, N4601, N4602, N4603, N4604, N4605,
         N4606, N4607, N4608, N4609, N4610, N4611, N4612, N4613, N4614, N4615,
         N4616, N4617, N4618, N4619, N4620, N4621, N4622, N4806, N4807, N4808,
         N4809, N4810, N4811, N4812, N4813, N4814, N4815, N4816, N4817, N4818,
         N4819, N4820, N4821, N4822, N4823, N4824, N4825, N4826, N4827, N4828,
         N4829, N4830, N4831, N4832, N4833, N4834, N4835, N4836, N4837, N4838,
         N4952, N4953, N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961,
         N4962, N4963, N4964, N4965, N4966, N4967, N4968, N4969, N4970, N4971,
         N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980, N4981,
         N4982, N4983, N4984, N5040, N5041, N5042, N5043, N5044, N5045, N5046,
         N5047, N5048, N5049, N5050, N5051, N5052, N5053, N5054, N5055, N5056,
         N5057, N5058, N5059, N5060, N5061, N5062, N5063, N5064, N5065, N5066,
         N5067, N5068, N5069, N5070, N5071, N5072, N5128, N5129, N5130, N5131,
         N5132, N5133, N5134, N5135, N5136, N5137, N5138, N5139, N5140, N5141,
         N5142, N5143, N5144, N5145, N5146, N5147, N5148, N5149, N5150, N5151,
         N5152, N5153, N5154, N5155, N5156, N5157, N5158, N5159, N5160, N5216,
         N5217, N5218, N5219, N5220, N5221, N5222, N5223, N5224, N5225, N5226,
         N5227, N5228, N5229, N5230, N5231, N5232, N5233, N5234, N5235, N5236,
         N5237, N5238, N5239, N5240, N5241, N5242, N5243, N5244, N5245, N5246,
         N5247, N5248, N5304, N5305, N5306, N5307, N5308, N5309, N5310, N5311,
         N5312, N5313, N5314, N5315, N5316, N5317, N5318, N5319, N5320, N5321,
         N5322, N5323, N5324, N5325, N5326, N5327, N5328, N5329, N5330, N5331,
         N5332, N5333, N5334, N5335, N5336, N5392, N5393, N5394, N5395, N5396,
         N5397, N5398, N5399, N5400, N5401, N5402, N5403, N5404, N5405, N5406,
         N5407, N5408, N5409, N5410, N5411, N5412, N5413, N5414, N5415, N5416,
         N5417, N5418, N5419, N5420, N5421, N5422, N5423, N5424, N5480, N5481,
         N5482, N5483, N5484, N5485, N5486, N5487, N5488, N5489, N5490, N5491,
         N5492, N5493, N5494, N5495, N5496, N5497, N5498, N5499, N5500, N5501,
         N5502, N5503, N5504, N5505, N5506, N5507, N5508, N5509, N5510, N5511,
         N5512, N5568, N5569, N5570, N5571, N5572, N5573, N5574, N5575, N5576,
         N5577, N5578, N5579, N5580, N5581, N5582, N5583, N5584, N5585, N5586,
         N5587, N5588, N5589, N5590, N5591, N5592, N5593, N5594, N5595, N5596,
         N5597, N5598, N5599, N5600, N5656, N5657, N5658, N5659, N5660, N5661,
         N5662, N5663, N5664, N5665, N5666, N5667, N5668, N5669, N5670, N5671,
         N5672, N5673, N5674, N5675, N5676, N5677, N5678, N5679, N5680, N5681,
         N5682, N5683, N5684, N5685, N5686, N5687, N5688, N5802, N5803, N5804,
         N5805, N5806, N5807, N5808, N5809, N5810, N5811, N5812, N5813, N5814,
         N5815, N5816, N5817, N5818, N5819, N5820, N5821, N5822, N5823, N5824,
         N5825, N5826, N5827, N5828, N5829, N5830, N5831, N5832, N5833, N5834,
         N6018, N6019, N6020, N6021, N6022, N6023, N6024, N6025, N6026, N6027,
         N6028, N6029, N6030, N6031, N6032, N6033, N6034, N6035, N6036, N6037,
         N6038, N6039, N6040, N6041, N6042, N6043, N6044, N6045, N6046, N6047,
         N6048, N6049, N6050, N6234, N6235, N6236, N6237, N6238, N6239, N6240,
         N6241, N6242, N6243, N6244, N6245, N6246, N6247, N6248, N6249, N6250,
         N6251, N6252, N6253, N6254, N6255, N6256, N6257, N6258, N6259, N6260,
         N6261, N6262, N6263, N6264, N6265, N6266, N6450, N6451, N6452, N6453,
         N6454, N6455, N6456, N6457, N6458, N6459, N6460, N6461, N6462, N6463,
         N6464, N6465, N6466, N6467, N6468, N6469, N6470, N6471, N6472, N6473,
         N6474, N6475, N6476, N6477, N6478, N6479, N6480, N6481, N6482, N6666,
         N6667, N6668, N6669, N6670, N6671, N6672, N6673, N6674, N6675, N6676,
         N6677, N6678, N6679, N6680, N6681, N6682, N6683, N6684, N6685, N6686,
         N6687, N6688, N6689, N6690, N6691, N6692, N6693, N6694, N6695, N6696,
         N6697, N6698, N6882, N6883, N6884, N6885, N6886, N6887, N6888, N6889,
         N6890, N6891, N6892, N6893, N6894, N6895, N6896, N6897, N6898, N6899,
         N6900, N6901, N6902, N6903, N6904, N6905, N6906, N6907, N6908, N6909,
         N6910, N6911, N6912, N6913, N6914, N7098, N7099, N7100, N7101, N7102,
         N7103, N7104, N7105, N7106, N7107, N7108, N7109, N7110, N7111, N7112,
         N7113, N7114, N7115, N7116, N7117, N7118, N7119, N7120, N7121, N7122,
         N7123, N7124, N7125, N7126, N7127, N7128, N7129, N7130, N7314, N7315,
         N7316, N7317, N7318, N7319, N7320, N7321, N7322, N7323, N7324, N7325,
         N7326, N7327, N7328, N7329, N7330, N7331, N7332, N7333, N7334, N7335,
         N7336, N7337, N7338, N7339, N7340, N7341, N7342, N7343, N7344, N7345,
         N7346, N7531, N7532, N7533, N7534, N7535, N7536, N7537, N7538, N7539,
         N7540, N7541, N7542, N7543, N7544, N7545, N7546, N7547, N7548, N7549,
         N7550, N7551, N7552, N7553, N7554, N7555, N7556, N7557, N7558, N7559,
         N7560, N7561, N7562, N7676, N7677, N7678, N7679, N7680, N7681, N7682,
         N7683, N7684, N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692,
         N7693, N7694, N7695, N7696, N7697, N7698, N7699, N7700, N7701, N7702,
         N7703, N7704, N7705, N7706, N7707, N7708, N7764, N7765, N7766, N7767,
         N7768, N7769, N7770, N7771, N7772, N7773, N7774, N7775, N7776, N7777,
         N7778, N7779, N7780, N7781, N7782, N7783, N7784, N7785, N7786, N7787,
         N7788, N7789, N7790, N7791, N7792, N7793, N7794, N7795, N7796, N7852,
         N7853, N7854, N7855, N7856, N7857, N7858, N7859, N7860, N7861, N7862,
         N7863, N7864, N7865, N7866, N7867, N7868, N7869, N7870, N7871, N7872,
         N7873, N7874, N7875, N7876, N7877, N7878, N7879, N7880, N7881, N7882,
         N7883, N7884, N7940, N7941, N7942, N7943, N7944, N7945, N7946, N7947,
         N7948, N7949, N7950, N7951, N7952, N7953, N7954, N7955, N7956, N7957,
         N7958, N7959, N7960, N7961, N7962, N7963, N7964, N7965, N7966, N7967,
         N7968, N7969, N7970, N7971, N7972, N8028, N8029, N8030, N8031, N8032,
         N8033, N8034, N8035, N8036, N8037, N8038, N8039, N8040, N8041, N8042,
         N8043, N8044, N8045, N8046, N8047, N8048, N8049, N8050, N8051, N8052,
         N8053, N8054, N8055, N8056, N8057, N8058, N8059, N8060, N8116, N8117,
         N8118, N8119, N8120, N8121, N8122, N8123, N8124, N8125, N8126, N8127,
         N8128, N8129, N8130, N8131, N8132, N8133, N8134, N8135, N8136, N8137,
         N8138, N8139, N8140, N8141, N8142, N8143, N8144, N8145, N8146, N8147,
         N8148, N8204, N8205, N8206, N8207, N8208, N8209, N8210, N8211, N8212,
         N8213, N8214, N8215, N8216, N8217, N8218, N8219, N8220, N8221, N8222,
         N8223, N8224, N8225, N8226, N8227, N8228, N8229, N8230, N8231, N8232,
         N8233, N8234, N8235, N8236, N8292, N8293, N8294, N8295, N8296, N8297,
         N8298, N8299, N8300, N8301, N8302, N8303, N8304, N8305, N8306, N8307,
         N8308, N8309, N8310, N8311, N8312, N8313, N8314, N8315, N8316, N8317,
         N8318, N8319, N8320, N8321, N8322, N8323, N8324, N8380, N8381, N8382,
         N8383, N8384, N8385, N8386, N8387, N8388, N8389, N8390, N8391, N8392,
         N8393, N8394, N8395, N8396, N8397, N8398, N8399, N8400, N8401, N8402,
         N8403, N8404, N8405, N8406, N8407, N8408, N8409, N8410, N8411, N8412,
         N8526, N8527, N8528, N8529, N8530, N8531, N8532, N8533, N8534, N8535,
         N8536, N8537, N8538, N8539, N8540, N8541, N8542, N8543, N8544, N8545,
         N8546, N8547, N8548, N8549, N8550, N8551, N8552, N8553, N8554, N8555,
         N8556, N8557, N8558, N8742, N8743, N8744, N8745, N8746, N8747, N8748,
         N8749, N8750, N8751, N8752, N8753, N8754, N8755, N8756, N8757, N8758,
         N8759, N8760, N8761, N8762, N8763, N8764, N8765, N8766, N8767, N8768,
         N8769, N8770, N8771, N8772, N8773, N8774, N8958, N8959, N8960, N8961,
         N8962, N8963, N8964, N8965, N8966, N8967, N8968, N8969, N8970, N8971,
         N8972, N8973, N8974, N8975, N8976, N8977, N8978, N8979, N8980, N8981,
         N8982, N8983, N8984, N8985, N8986, N8987, N8988, N8989, N8990, N9174,
         N9175, N9176, N9177, N9178, N9179, N9180, N9181, N9182, N9183, N9184,
         N9185, N9186, N9187, N9188, N9189, N9190, N9191, N9192, N9193, N9194,
         N9195, N9196, N9197, N9198, N9199, N9200, N9201, N9202, N9203, N9204,
         N9205, N9206, N9390, N9391, N9392, N9393, N9394, N9395, N9396, N9397,
         N9398, N9399, N9400, N9401, N9402, N9403, N9404, N9405, N9406, N9407,
         N9408, N9409, N9410, N9411, N9412, N9413, N9414, N9415, N9416, N9417,
         N9418, N9419, N9420, N9421, N9422, N9606, N9607, N9608, N9609, N9610,
         N9611, N9612, N9613, N9614, N9615, N9616, N9617, N9618, N9619, N9620,
         N9621, N9622, N9623, N9624, N9625, N9626, N9627, N9628, N9629, N9630,
         N9631, N9632, N9633, N9634, N9635, N9636, N9637, N9638, N9822, N9823,
         N9824, N9825, N9826, N9827, N9828, N9829, N9830, N9831, N9832, N9833,
         N9834, N9835, N9836, N9837, N9838, N9839, N9840, N9841, N9842, N9843,
         N9844, N9845, N9846, N9847, N9848, N9849, N9850, N9851, N9852, N9853,
         N9854, N10038, N10039, N10040, N10041, N10042, N10043, N10044, N10045,
         N10046, N10047, N10048, N10049, N10050, N10051, N10052, N10053,
         N10054, N10055, N10056, N10057, N10058, N10059, N10060, N10061,
         N10062, N10063, N10064, N10065, N10066, N10067, N10068, N10069,
         N10070, N10254, N10255, N10256, N10257, N10258, N10259, N10260,
         N10261, N10262, N10263, N10264, N10265, N10266, N10267, N10268,
         N10269, N10270, N10271, N10272, N10273, N10274, N10275, N10276,
         N10277, N10278, N10279, N10280, N10281, N10282, N10283, N10284,
         N10285, N10286, N10400, N10401, N10402, N10403, N10404, N10405,
         N10406, N10407, N10408, N10409, N10410, N10411, N10412, N10413,
         N10414, N10415, N10416, N10417, N10418, N10419, N10420, N10421,
         N10422, N10423, N10424, N10425, N10426, N10427, N10428, N10429,
         N10430, N10431, N10432, N10488, N10489, N10490, N10491, N10492,
         N10493, N10494, N10495, N10496, N10497, N10498, N10499, N10500,
         N10501, N10502, N10503, N10504, N10505, N10506, N10507, N10508,
         N10509, N10510, N10511, N10512, N10513, N10514, N10515, N10516,
         N10517, N10518, N10519, N10520, N10576, N10577, N10578, N10579,
         N10580, N10581, N10582, N10583, N10584, N10585, N10586, N10587,
         N10588, N10589, N10590, N10591, N10592, N10593, N10594, N10595,
         N10596, N10597, N10598, N10599, N10600, N10601, N10602, N10603,
         N10604, N10605, N10606, N10607, N10608, N10664, N10665, N10666,
         N10667, N10668, N10669, N10670, N10671, N10672, N10673, N10674,
         N10675, N10676, N10677, N10678, N10679, N10680, N10681, N10682,
         N10683, N10684, N10685, N10686, N10687, N10688, N10689, N10690,
         N10691, N10692, N10693, N10694, N10695, N10696, N10752, N10753,
         N10754, N10755, N10756, N10757, N10758, N10759, N10760, N10761,
         N10762, N10763, N10764, N10765, N10766, N10767, N10768, N10769,
         N10770, N10771, N10772, N10773, N10774, N10775, N10776, N10777,
         N10778, N10779, N10780, N10781, N10782, N10783, N10784, N10840,
         N10841, N10842, N10843, N10844, N10845, N10846, N10847, N10848,
         N10849, N10850, N10851, N10852, N10853, N10854, N10855, N10856,
         N10857, N10858, N10859, N10860, N10861, N10862, N10863, N10864,
         N10865, N10866, N10867, N10868, N10869, N10870, N10871, N10872,
         N10928, N10929, N10930, N10931, N10932, N10933, N10934, N10935,
         N10936, N10937, N10938, N10939, N10940, N10941, N10942, N10943,
         N10944, N10945, N10946, N10947, N10948, N10949, N10950, N10951,
         N10952, N10953, N10954, N10955, N10956, N10957, N10958, N10959,
         N10960, N11016, N11017, N11018, N11019, N11020, N11021, N11022,
         N11023, N11024, N11025, N11026, N11027, N11028, N11029, N11030,
         N11031, N11032, N11033, N11034, N11035, N11036, N11037, N11038,
         N11039, N11040, N11041, N11042, N11043, N11044, N11045, N11046,
         N11047, N11048, N11104, N11105, N11106, N11107, N11108, N11109,
         N11110, N11111, N11112, N11113, N11114, N11115, N11116, N11117,
         N11118, N11119, N11120, N11121, N11122, N11123, N11124, N11125,
         N11126, N11127, N11128, N11129, N11130, N11131, N11132, N11133,
         N11134, N11135, N11136, N11250, N11251, N11252, N11253, N11254,
         N11255, N11256, N11257, N11258, N11259, N11260, N11261, N11262,
         N11263, N11264, N11265, N11266, N11267, N11268, N11269, N11270,
         N11271, N11272, N11273, N11274, N11275, N11276, N11277, N11278,
         N11279, N11280, N11281, N11282, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304;
  wire   [2047:0] inner_first_stage_data_reg;
  wire   [63:0] inner_first_stage_valid_reg;

  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_0_ ( .D(N542), .CP(clk), 
        .Q(inner_first_stage_valid_reg[0]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_31_ ( .D(N574), .CP(clk), 
        .Q(inner_first_stage_data_reg[31]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_30_ ( .D(N573), .CP(clk), 
        .Q(inner_first_stage_data_reg[30]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_29_ ( .D(N572), .CP(clk), 
        .Q(inner_first_stage_data_reg[29]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_28_ ( .D(N571), .CP(clk), 
        .Q(inner_first_stage_data_reg[28]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_27_ ( .D(N570), .CP(clk), 
        .Q(inner_first_stage_data_reg[27]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_26_ ( .D(N569), .CP(clk), 
        .Q(inner_first_stage_data_reg[26]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_25_ ( .D(N568), .CP(clk), 
        .Q(inner_first_stage_data_reg[25]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_24_ ( .D(N567), .CP(clk), 
        .Q(inner_first_stage_data_reg[24]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_23_ ( .D(N566), .CP(clk), 
        .Q(inner_first_stage_data_reg[23]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_22_ ( .D(N565), .CP(clk), 
        .Q(inner_first_stage_data_reg[22]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_21_ ( .D(N564), .CP(clk), 
        .Q(inner_first_stage_data_reg[21]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_20_ ( .D(N563), .CP(clk), 
        .Q(inner_first_stage_data_reg[20]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_19_ ( .D(N562), .CP(clk), 
        .Q(inner_first_stage_data_reg[19]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_18_ ( .D(N561), .CP(clk), 
        .Q(inner_first_stage_data_reg[18]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_17_ ( .D(N560), .CP(clk), 
        .Q(inner_first_stage_data_reg[17]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_16_ ( .D(N559), .CP(clk), 
        .Q(inner_first_stage_data_reg[16]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_15_ ( .D(N558), .CP(clk), 
        .Q(inner_first_stage_data_reg[15]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_14_ ( .D(N557), .CP(clk), 
        .Q(inner_first_stage_data_reg[14]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_13_ ( .D(N556), .CP(clk), 
        .Q(inner_first_stage_data_reg[13]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_12_ ( .D(N555), .CP(clk), 
        .Q(inner_first_stage_data_reg[12]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_11_ ( .D(N554), .CP(clk), 
        .Q(inner_first_stage_data_reg[11]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_10_ ( .D(N553), .CP(clk), 
        .Q(inner_first_stage_data_reg[10]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_9_ ( .D(N552), .CP(clk), 
        .Q(inner_first_stage_data_reg[9]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_8_ ( .D(N551), .CP(clk), 
        .Q(inner_first_stage_data_reg[8]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_7_ ( .D(N550), .CP(clk), 
        .Q(inner_first_stage_data_reg[7]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_6_ ( .D(N549), .CP(clk), 
        .Q(inner_first_stage_data_reg[6]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_5_ ( .D(N548), .CP(clk), 
        .Q(inner_first_stage_data_reg[5]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_4_ ( .D(N547), .CP(clk), 
        .Q(inner_first_stage_data_reg[4]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_3_ ( .D(N546), .CP(clk), 
        .Q(inner_first_stage_data_reg[3]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2_ ( .D(N545), .CP(clk), 
        .Q(inner_first_stage_data_reg[2]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1_ ( .D(N544), .CP(clk), 
        .Q(inner_first_stage_data_reg[1]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_0_ ( .D(N543), .CP(clk), 
        .Q(inner_first_stage_data_reg[0]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_1_ ( .D(N762), .CP(clk), 
        .Q(inner_first_stage_valid_reg[1]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_63_ ( .D(N794), .CP(clk), 
        .Q(inner_first_stage_data_reg[63]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_62_ ( .D(N793), .CP(clk), 
        .Q(inner_first_stage_data_reg[62]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_61_ ( .D(N792), .CP(clk), 
        .Q(inner_first_stage_data_reg[61]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_60_ ( .D(N791), .CP(clk), 
        .Q(inner_first_stage_data_reg[60]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_59_ ( .D(N790), .CP(clk), 
        .Q(inner_first_stage_data_reg[59]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_58_ ( .D(N789), .CP(clk), 
        .Q(inner_first_stage_data_reg[58]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_57_ ( .D(N788), .CP(clk), 
        .Q(inner_first_stage_data_reg[57]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_56_ ( .D(N787), .CP(clk), 
        .Q(inner_first_stage_data_reg[56]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_55_ ( .D(N786), .CP(clk), 
        .Q(inner_first_stage_data_reg[55]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_54_ ( .D(N785), .CP(clk), 
        .Q(inner_first_stage_data_reg[54]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_53_ ( .D(N784), .CP(clk), 
        .Q(inner_first_stage_data_reg[53]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_52_ ( .D(N783), .CP(clk), 
        .Q(inner_first_stage_data_reg[52]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_51_ ( .D(N782), .CP(clk), 
        .Q(inner_first_stage_data_reg[51]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_50_ ( .D(N781), .CP(clk), 
        .Q(inner_first_stage_data_reg[50]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_49_ ( .D(N780), .CP(clk), 
        .Q(inner_first_stage_data_reg[49]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_48_ ( .D(N779), .CP(clk), 
        .Q(inner_first_stage_data_reg[48]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_47_ ( .D(N778), .CP(clk), 
        .Q(inner_first_stage_data_reg[47]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_46_ ( .D(N777), .CP(clk), 
        .Q(inner_first_stage_data_reg[46]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_45_ ( .D(N776), .CP(clk), 
        .Q(inner_first_stage_data_reg[45]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_44_ ( .D(N775), .CP(clk), 
        .Q(inner_first_stage_data_reg[44]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_43_ ( .D(N774), .CP(clk), 
        .Q(inner_first_stage_data_reg[43]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_42_ ( .D(N773), .CP(clk), 
        .Q(inner_first_stage_data_reg[42]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_41_ ( .D(N772), .CP(clk), 
        .Q(inner_first_stage_data_reg[41]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_40_ ( .D(N771), .CP(clk), 
        .Q(inner_first_stage_data_reg[40]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_39_ ( .D(N770), .CP(clk), 
        .Q(inner_first_stage_data_reg[39]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_38_ ( .D(N769), .CP(clk), 
        .Q(inner_first_stage_data_reg[38]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_37_ ( .D(N768), .CP(clk), 
        .Q(inner_first_stage_data_reg[37]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_36_ ( .D(N767), .CP(clk), 
        .Q(inner_first_stage_data_reg[36]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_35_ ( .D(N766), .CP(clk), 
        .Q(inner_first_stage_data_reg[35]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_34_ ( .D(N765), .CP(clk), 
        .Q(inner_first_stage_data_reg[34]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_33_ ( .D(N764), .CP(clk), 
        .Q(inner_first_stage_data_reg[33]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_32_ ( .D(N763), .CP(clk), 
        .Q(inner_first_stage_data_reg[32]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_2_ ( .D(N982), .CP(clk), 
        .Q(inner_first_stage_valid_reg[2]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_95_ ( .D(N1014), .CP(clk), 
        .Q(inner_first_stage_data_reg[95]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_94_ ( .D(N1013), .CP(clk), 
        .Q(inner_first_stage_data_reg[94]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_93_ ( .D(N1012), .CP(clk), 
        .Q(inner_first_stage_data_reg[93]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_92_ ( .D(N1011), .CP(clk), 
        .Q(inner_first_stage_data_reg[92]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_91_ ( .D(N1010), .CP(clk), 
        .Q(inner_first_stage_data_reg[91]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_90_ ( .D(N1009), .CP(clk), 
        .Q(inner_first_stage_data_reg[90]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_89_ ( .D(N1008), .CP(clk), 
        .Q(inner_first_stage_data_reg[89]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_88_ ( .D(N1007), .CP(clk), 
        .Q(inner_first_stage_data_reg[88]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_87_ ( .D(N1006), .CP(clk), 
        .Q(inner_first_stage_data_reg[87]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_86_ ( .D(N1005), .CP(clk), 
        .Q(inner_first_stage_data_reg[86]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_85_ ( .D(N1004), .CP(clk), 
        .Q(inner_first_stage_data_reg[85]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_84_ ( .D(N1003), .CP(clk), 
        .Q(inner_first_stage_data_reg[84]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_83_ ( .D(N1002), .CP(clk), 
        .Q(inner_first_stage_data_reg[83]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_82_ ( .D(N1001), .CP(clk), 
        .Q(inner_first_stage_data_reg[82]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_81_ ( .D(N1000), .CP(clk), 
        .Q(inner_first_stage_data_reg[81]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_80_ ( .D(N999), .CP(clk), 
        .Q(inner_first_stage_data_reg[80]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_79_ ( .D(N998), .CP(clk), 
        .Q(inner_first_stage_data_reg[79]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_78_ ( .D(N997), .CP(clk), 
        .Q(inner_first_stage_data_reg[78]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_77_ ( .D(N996), .CP(clk), 
        .Q(inner_first_stage_data_reg[77]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_76_ ( .D(N995), .CP(clk), 
        .Q(inner_first_stage_data_reg[76]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_75_ ( .D(N994), .CP(clk), 
        .Q(inner_first_stage_data_reg[75]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_74_ ( .D(N993), .CP(clk), 
        .Q(inner_first_stage_data_reg[74]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_73_ ( .D(N992), .CP(clk), 
        .Q(inner_first_stage_data_reg[73]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_72_ ( .D(N991), .CP(clk), 
        .Q(inner_first_stage_data_reg[72]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_71_ ( .D(N990), .CP(clk), 
        .Q(inner_first_stage_data_reg[71]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_70_ ( .D(N989), .CP(clk), 
        .Q(inner_first_stage_data_reg[70]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_69_ ( .D(N988), .CP(clk), 
        .Q(inner_first_stage_data_reg[69]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_68_ ( .D(N987), .CP(clk), 
        .Q(inner_first_stage_data_reg[68]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_67_ ( .D(N986), .CP(clk), 
        .Q(inner_first_stage_data_reg[67]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_66_ ( .D(N985), .CP(clk), 
        .Q(inner_first_stage_data_reg[66]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_65_ ( .D(N984), .CP(clk), 
        .Q(inner_first_stage_data_reg[65]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_64_ ( .D(N983), .CP(clk), 
        .Q(inner_first_stage_data_reg[64]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_3_ ( .D(N1202), .CP(clk), 
        .Q(inner_first_stage_valid_reg[3]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_127_ ( .D(N1234), .CP(clk), 
        .Q(inner_first_stage_data_reg[127]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_126_ ( .D(N1233), .CP(clk), 
        .Q(inner_first_stage_data_reg[126]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_125_ ( .D(N1232), .CP(clk), 
        .Q(inner_first_stage_data_reg[125]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_124_ ( .D(N1231), .CP(clk), 
        .Q(inner_first_stage_data_reg[124]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_123_ ( .D(N1230), .CP(clk), 
        .Q(inner_first_stage_data_reg[123]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_122_ ( .D(N1229), .CP(clk), 
        .Q(inner_first_stage_data_reg[122]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_121_ ( .D(N1228), .CP(clk), 
        .Q(inner_first_stage_data_reg[121]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_120_ ( .D(N1227), .CP(clk), 
        .Q(inner_first_stage_data_reg[120]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_119_ ( .D(N1226), .CP(clk), 
        .Q(inner_first_stage_data_reg[119]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_118_ ( .D(N1225), .CP(clk), 
        .Q(inner_first_stage_data_reg[118]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_117_ ( .D(N1224), .CP(clk), 
        .Q(inner_first_stage_data_reg[117]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_116_ ( .D(N1223), .CP(clk), 
        .Q(inner_first_stage_data_reg[116]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_115_ ( .D(N1222), .CP(clk), 
        .Q(inner_first_stage_data_reg[115]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_114_ ( .D(N1221), .CP(clk), 
        .Q(inner_first_stage_data_reg[114]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_113_ ( .D(N1220), .CP(clk), 
        .Q(inner_first_stage_data_reg[113]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_112_ ( .D(N1219), .CP(clk), 
        .Q(inner_first_stage_data_reg[112]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_111_ ( .D(N1218), .CP(clk), 
        .Q(inner_first_stage_data_reg[111]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_110_ ( .D(N1217), .CP(clk), 
        .Q(inner_first_stage_data_reg[110]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_109_ ( .D(N1216), .CP(clk), 
        .Q(inner_first_stage_data_reg[109]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_108_ ( .D(N1215), .CP(clk), 
        .Q(inner_first_stage_data_reg[108]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_107_ ( .D(N1214), .CP(clk), 
        .Q(inner_first_stage_data_reg[107]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_106_ ( .D(N1213), .CP(clk), 
        .Q(inner_first_stage_data_reg[106]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_105_ ( .D(N1212), .CP(clk), 
        .Q(inner_first_stage_data_reg[105]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_104_ ( .D(N1211), .CP(clk), 
        .Q(inner_first_stage_data_reg[104]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_103_ ( .D(N1210), .CP(clk), 
        .Q(inner_first_stage_data_reg[103]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_102_ ( .D(N1209), .CP(clk), 
        .Q(inner_first_stage_data_reg[102]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_101_ ( .D(N1208), .CP(clk), 
        .Q(inner_first_stage_data_reg[101]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_100_ ( .D(N1207), .CP(clk), 
        .Q(inner_first_stage_data_reg[100]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_99_ ( .D(N1206), .CP(clk), 
        .Q(inner_first_stage_data_reg[99]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_98_ ( .D(N1205), .CP(clk), 
        .Q(inner_first_stage_data_reg[98]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_97_ ( .D(N1204), .CP(clk), 
        .Q(inner_first_stage_data_reg[97]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_96_ ( .D(N1203), .CP(clk), 
        .Q(inner_first_stage_data_reg[96]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_4_ ( .D(N1422), .CP(clk), 
        .Q(inner_first_stage_valid_reg[4]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_159_ ( .D(N1454), .CP(clk), 
        .Q(inner_first_stage_data_reg[159]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_158_ ( .D(N1453), .CP(clk), 
        .Q(inner_first_stage_data_reg[158]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_157_ ( .D(N1452), .CP(clk), 
        .Q(inner_first_stage_data_reg[157]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_156_ ( .D(N1451), .CP(clk), 
        .Q(inner_first_stage_data_reg[156]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_155_ ( .D(N1450), .CP(clk), 
        .Q(inner_first_stage_data_reg[155]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_154_ ( .D(N1449), .CP(clk), 
        .Q(inner_first_stage_data_reg[154]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_153_ ( .D(N1448), .CP(clk), 
        .Q(inner_first_stage_data_reg[153]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_152_ ( .D(N1447), .CP(clk), 
        .Q(inner_first_stage_data_reg[152]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_151_ ( .D(N1446), .CP(clk), 
        .Q(inner_first_stage_data_reg[151]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_150_ ( .D(N1445), .CP(clk), 
        .Q(inner_first_stage_data_reg[150]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_149_ ( .D(N1444), .CP(clk), 
        .Q(inner_first_stage_data_reg[149]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_148_ ( .D(N1443), .CP(clk), 
        .Q(inner_first_stage_data_reg[148]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_147_ ( .D(N1442), .CP(clk), 
        .Q(inner_first_stage_data_reg[147]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_146_ ( .D(N1441), .CP(clk), 
        .Q(inner_first_stage_data_reg[146]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_145_ ( .D(N1440), .CP(clk), 
        .Q(inner_first_stage_data_reg[145]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_144_ ( .D(N1439), .CP(clk), 
        .Q(inner_first_stage_data_reg[144]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_143_ ( .D(N1438), .CP(clk), 
        .Q(inner_first_stage_data_reg[143]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_142_ ( .D(N1437), .CP(clk), 
        .Q(inner_first_stage_data_reg[142]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_141_ ( .D(N1436), .CP(clk), 
        .Q(inner_first_stage_data_reg[141]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_140_ ( .D(N1435), .CP(clk), 
        .Q(inner_first_stage_data_reg[140]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_139_ ( .D(N1434), .CP(clk), 
        .Q(inner_first_stage_data_reg[139]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_138_ ( .D(N1433), .CP(clk), 
        .Q(inner_first_stage_data_reg[138]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_137_ ( .D(N1432), .CP(clk), 
        .Q(inner_first_stage_data_reg[137]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_136_ ( .D(N1431), .CP(clk), 
        .Q(inner_first_stage_data_reg[136]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_135_ ( .D(N1430), .CP(clk), 
        .Q(inner_first_stage_data_reg[135]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_134_ ( .D(N1429), .CP(clk), 
        .Q(inner_first_stage_data_reg[134]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_133_ ( .D(N1428), .CP(clk), 
        .Q(inner_first_stage_data_reg[133]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_132_ ( .D(N1427), .CP(clk), 
        .Q(inner_first_stage_data_reg[132]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_131_ ( .D(N1426), .CP(clk), 
        .Q(inner_first_stage_data_reg[131]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_130_ ( .D(N1425), .CP(clk), 
        .Q(inner_first_stage_data_reg[130]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_129_ ( .D(N1424), .CP(clk), 
        .Q(inner_first_stage_data_reg[129]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_128_ ( .D(N1423), .CP(clk), 
        .Q(inner_first_stage_data_reg[128]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_5_ ( .D(N1642), .CP(clk), 
        .Q(inner_first_stage_valid_reg[5]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_191_ ( .D(N1674), .CP(clk), 
        .Q(inner_first_stage_data_reg[191]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_190_ ( .D(N1673), .CP(clk), 
        .Q(inner_first_stage_data_reg[190]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_189_ ( .D(N1672), .CP(clk), 
        .Q(inner_first_stage_data_reg[189]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_188_ ( .D(N1671), .CP(clk), 
        .Q(inner_first_stage_data_reg[188]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_187_ ( .D(N1670), .CP(clk), 
        .Q(inner_first_stage_data_reg[187]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_186_ ( .D(N1669), .CP(clk), 
        .Q(inner_first_stage_data_reg[186]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_185_ ( .D(N1668), .CP(clk), 
        .Q(inner_first_stage_data_reg[185]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_184_ ( .D(N1667), .CP(clk), 
        .Q(inner_first_stage_data_reg[184]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_183_ ( .D(N1666), .CP(clk), 
        .Q(inner_first_stage_data_reg[183]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_182_ ( .D(N1665), .CP(clk), 
        .Q(inner_first_stage_data_reg[182]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_181_ ( .D(N1664), .CP(clk), 
        .Q(inner_first_stage_data_reg[181]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_180_ ( .D(N1663), .CP(clk), 
        .Q(inner_first_stage_data_reg[180]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_179_ ( .D(N1662), .CP(clk), 
        .Q(inner_first_stage_data_reg[179]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_178_ ( .D(N1661), .CP(clk), 
        .Q(inner_first_stage_data_reg[178]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_177_ ( .D(N1660), .CP(clk), 
        .Q(inner_first_stage_data_reg[177]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_176_ ( .D(N1659), .CP(clk), 
        .Q(inner_first_stage_data_reg[176]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_175_ ( .D(N1658), .CP(clk), 
        .Q(inner_first_stage_data_reg[175]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_174_ ( .D(N1657), .CP(clk), 
        .Q(inner_first_stage_data_reg[174]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_173_ ( .D(N1656), .CP(clk), 
        .Q(inner_first_stage_data_reg[173]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_172_ ( .D(N1655), .CP(clk), 
        .Q(inner_first_stage_data_reg[172]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_171_ ( .D(N1654), .CP(clk), 
        .Q(inner_first_stage_data_reg[171]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_170_ ( .D(N1653), .CP(clk), 
        .Q(inner_first_stage_data_reg[170]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_169_ ( .D(N1652), .CP(clk), 
        .Q(inner_first_stage_data_reg[169]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_168_ ( .D(N1651), .CP(clk), 
        .Q(inner_first_stage_data_reg[168]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_167_ ( .D(N1650), .CP(clk), 
        .Q(inner_first_stage_data_reg[167]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_166_ ( .D(N1649), .CP(clk), 
        .Q(inner_first_stage_data_reg[166]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_165_ ( .D(N1648), .CP(clk), 
        .Q(inner_first_stage_data_reg[165]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_164_ ( .D(N1647), .CP(clk), 
        .Q(inner_first_stage_data_reg[164]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_163_ ( .D(N1646), .CP(clk), 
        .Q(inner_first_stage_data_reg[163]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_162_ ( .D(N1645), .CP(clk), 
        .Q(inner_first_stage_data_reg[162]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_161_ ( .D(N1644), .CP(clk), 
        .Q(inner_first_stage_data_reg[161]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_160_ ( .D(N1643), .CP(clk), 
        .Q(inner_first_stage_data_reg[160]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_6_ ( .D(N1862), .CP(clk), 
        .Q(inner_first_stage_valid_reg[6]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_223_ ( .D(N1894), .CP(clk), 
        .Q(inner_first_stage_data_reg[223]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_222_ ( .D(N1893), .CP(clk), 
        .Q(inner_first_stage_data_reg[222]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_221_ ( .D(N1892), .CP(clk), 
        .Q(inner_first_stage_data_reg[221]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_220_ ( .D(N1891), .CP(clk), 
        .Q(inner_first_stage_data_reg[220]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_219_ ( .D(N1890), .CP(clk), 
        .Q(inner_first_stage_data_reg[219]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_218_ ( .D(N1889), .CP(clk), 
        .Q(inner_first_stage_data_reg[218]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_217_ ( .D(N1888), .CP(clk), 
        .Q(inner_first_stage_data_reg[217]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_216_ ( .D(N1887), .CP(clk), 
        .Q(inner_first_stage_data_reg[216]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_215_ ( .D(N1886), .CP(clk), 
        .Q(inner_first_stage_data_reg[215]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_214_ ( .D(N1885), .CP(clk), 
        .Q(inner_first_stage_data_reg[214]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_213_ ( .D(N1884), .CP(clk), 
        .Q(inner_first_stage_data_reg[213]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_212_ ( .D(N1883), .CP(clk), 
        .Q(inner_first_stage_data_reg[212]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_211_ ( .D(N1882), .CP(clk), 
        .Q(inner_first_stage_data_reg[211]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_210_ ( .D(N1881), .CP(clk), 
        .Q(inner_first_stage_data_reg[210]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_209_ ( .D(N1880), .CP(clk), 
        .Q(inner_first_stage_data_reg[209]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_208_ ( .D(N1879), .CP(clk), 
        .Q(inner_first_stage_data_reg[208]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_207_ ( .D(N1878), .CP(clk), 
        .Q(inner_first_stage_data_reg[207]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_206_ ( .D(N1877), .CP(clk), 
        .Q(inner_first_stage_data_reg[206]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_205_ ( .D(N1876), .CP(clk), 
        .Q(inner_first_stage_data_reg[205]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_204_ ( .D(N1875), .CP(clk), 
        .Q(inner_first_stage_data_reg[204]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_203_ ( .D(N1874), .CP(clk), 
        .Q(inner_first_stage_data_reg[203]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_202_ ( .D(N1873), .CP(clk), 
        .Q(inner_first_stage_data_reg[202]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_201_ ( .D(N1872), .CP(clk), 
        .Q(inner_first_stage_data_reg[201]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_200_ ( .D(N1871), .CP(clk), 
        .Q(inner_first_stage_data_reg[200]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_199_ ( .D(N1870), .CP(clk), 
        .Q(inner_first_stage_data_reg[199]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_198_ ( .D(N1869), .CP(clk), 
        .Q(inner_first_stage_data_reg[198]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_197_ ( .D(N1868), .CP(clk), 
        .Q(inner_first_stage_data_reg[197]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_196_ ( .D(N1867), .CP(clk), 
        .Q(inner_first_stage_data_reg[196]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_195_ ( .D(N1866), .CP(clk), 
        .Q(inner_first_stage_data_reg[195]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_194_ ( .D(N1865), .CP(clk), 
        .Q(inner_first_stage_data_reg[194]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_193_ ( .D(N1864), .CP(clk), 
        .Q(inner_first_stage_data_reg[193]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_192_ ( .D(N1863), .CP(clk), 
        .Q(inner_first_stage_data_reg[192]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_7_ ( .D(N2082), .CP(clk), 
        .Q(inner_first_stage_valid_reg[7]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_255_ ( .D(N2114), .CP(clk), 
        .Q(inner_first_stage_data_reg[255]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_254_ ( .D(N2113), .CP(clk), 
        .Q(inner_first_stage_data_reg[254]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_253_ ( .D(N2112), .CP(clk), 
        .Q(inner_first_stage_data_reg[253]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_252_ ( .D(N2111), .CP(clk), 
        .Q(inner_first_stage_data_reg[252]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_251_ ( .D(N2110), .CP(clk), 
        .Q(inner_first_stage_data_reg[251]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_250_ ( .D(N2109), .CP(clk), 
        .Q(inner_first_stage_data_reg[250]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_249_ ( .D(N2108), .CP(clk), 
        .Q(inner_first_stage_data_reg[249]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_248_ ( .D(N2107), .CP(clk), 
        .Q(inner_first_stage_data_reg[248]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_247_ ( .D(N2106), .CP(clk), 
        .Q(inner_first_stage_data_reg[247]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_246_ ( .D(N2105), .CP(clk), 
        .Q(inner_first_stage_data_reg[246]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_245_ ( .D(N2104), .CP(clk), 
        .Q(inner_first_stage_data_reg[245]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_244_ ( .D(N2103), .CP(clk), 
        .Q(inner_first_stage_data_reg[244]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_243_ ( .D(N2102), .CP(clk), 
        .Q(inner_first_stage_data_reg[243]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_242_ ( .D(N2101), .CP(clk), 
        .Q(inner_first_stage_data_reg[242]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_241_ ( .D(N2100), .CP(clk), 
        .Q(inner_first_stage_data_reg[241]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_240_ ( .D(N2099), .CP(clk), 
        .Q(inner_first_stage_data_reg[240]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_239_ ( .D(N2098), .CP(clk), 
        .Q(inner_first_stage_data_reg[239]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_238_ ( .D(N2097), .CP(clk), 
        .Q(inner_first_stage_data_reg[238]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_237_ ( .D(N2096), .CP(clk), 
        .Q(inner_first_stage_data_reg[237]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_236_ ( .D(N2095), .CP(clk), 
        .Q(inner_first_stage_data_reg[236]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_235_ ( .D(N2094), .CP(clk), 
        .Q(inner_first_stage_data_reg[235]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_234_ ( .D(N2093), .CP(clk), 
        .Q(inner_first_stage_data_reg[234]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_233_ ( .D(N2092), .CP(clk), 
        .Q(inner_first_stage_data_reg[233]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_232_ ( .D(N2091), .CP(clk), 
        .Q(inner_first_stage_data_reg[232]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_231_ ( .D(N2090), .CP(clk), 
        .Q(inner_first_stage_data_reg[231]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_230_ ( .D(N2089), .CP(clk), 
        .Q(inner_first_stage_data_reg[230]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_229_ ( .D(N2088), .CP(clk), 
        .Q(inner_first_stage_data_reg[229]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_228_ ( .D(N2087), .CP(clk), 
        .Q(inner_first_stage_data_reg[228]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_227_ ( .D(N2086), .CP(clk), 
        .Q(inner_first_stage_data_reg[227]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_226_ ( .D(N2085), .CP(clk), 
        .Q(inner_first_stage_data_reg[226]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_225_ ( .D(N2084), .CP(clk), 
        .Q(inner_first_stage_data_reg[225]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_224_ ( .D(N2083), .CP(clk), 
        .Q(inner_first_stage_data_reg[224]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_8_ ( .D(N2316), .CP(clk), 
        .Q(inner_first_stage_valid_reg[8]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_287_ ( .D(N2348), .CP(clk), 
        .Q(inner_first_stage_data_reg[287]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_286_ ( .D(N2347), .CP(clk), 
        .Q(inner_first_stage_data_reg[286]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_285_ ( .D(N2346), .CP(clk), 
        .Q(inner_first_stage_data_reg[285]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_284_ ( .D(N2345), .CP(clk), 
        .Q(inner_first_stage_data_reg[284]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_283_ ( .D(N2344), .CP(clk), 
        .Q(inner_first_stage_data_reg[283]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_282_ ( .D(N2343), .CP(clk), 
        .Q(inner_first_stage_data_reg[282]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_281_ ( .D(N2342), .CP(clk), 
        .Q(inner_first_stage_data_reg[281]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_280_ ( .D(N2341), .CP(clk), 
        .Q(inner_first_stage_data_reg[280]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_279_ ( .D(N2340), .CP(clk), 
        .Q(inner_first_stage_data_reg[279]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_278_ ( .D(N2339), .CP(clk), 
        .Q(inner_first_stage_data_reg[278]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_277_ ( .D(N2338), .CP(clk), 
        .Q(inner_first_stage_data_reg[277]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_276_ ( .D(N2337), .CP(clk), 
        .Q(inner_first_stage_data_reg[276]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_275_ ( .D(N2336), .CP(clk), 
        .Q(inner_first_stage_data_reg[275]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_274_ ( .D(N2335), .CP(clk), 
        .Q(inner_first_stage_data_reg[274]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_273_ ( .D(N2334), .CP(clk), 
        .Q(inner_first_stage_data_reg[273]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_272_ ( .D(N2333), .CP(clk), 
        .Q(inner_first_stage_data_reg[272]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_271_ ( .D(N2332), .CP(clk), 
        .Q(inner_first_stage_data_reg[271]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_270_ ( .D(N2331), .CP(clk), 
        .Q(inner_first_stage_data_reg[270]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_269_ ( .D(N2330), .CP(clk), 
        .Q(inner_first_stage_data_reg[269]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_268_ ( .D(N2329), .CP(clk), 
        .Q(inner_first_stage_data_reg[268]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_267_ ( .D(N2328), .CP(clk), 
        .Q(inner_first_stage_data_reg[267]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_266_ ( .D(N2327), .CP(clk), 
        .Q(inner_first_stage_data_reg[266]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_265_ ( .D(N2326), .CP(clk), 
        .Q(inner_first_stage_data_reg[265]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_264_ ( .D(N2325), .CP(clk), 
        .Q(inner_first_stage_data_reg[264]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_263_ ( .D(N2324), .CP(clk), 
        .Q(inner_first_stage_data_reg[263]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_262_ ( .D(N2323), .CP(clk), 
        .Q(inner_first_stage_data_reg[262]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_261_ ( .D(N2322), .CP(clk), 
        .Q(inner_first_stage_data_reg[261]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_260_ ( .D(N2321), .CP(clk), 
        .Q(inner_first_stage_data_reg[260]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_259_ ( .D(N2320), .CP(clk), 
        .Q(inner_first_stage_data_reg[259]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_258_ ( .D(N2319), .CP(clk), 
        .Q(inner_first_stage_data_reg[258]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_257_ ( .D(N2318), .CP(clk), 
        .Q(inner_first_stage_data_reg[257]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_256_ ( .D(N2317), .CP(clk), 
        .Q(inner_first_stage_data_reg[256]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_9_ ( .D(N2404), .CP(clk), 
        .Q(inner_first_stage_valid_reg[9]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_319_ ( .D(N2436), .CP(clk), 
        .Q(inner_first_stage_data_reg[319]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_318_ ( .D(N2435), .CP(clk), 
        .Q(inner_first_stage_data_reg[318]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_317_ ( .D(N2434), .CP(clk), 
        .Q(inner_first_stage_data_reg[317]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_316_ ( .D(N2433), .CP(clk), 
        .Q(inner_first_stage_data_reg[316]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_315_ ( .D(N2432), .CP(clk), 
        .Q(inner_first_stage_data_reg[315]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_314_ ( .D(N2431), .CP(clk), 
        .Q(inner_first_stage_data_reg[314]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_313_ ( .D(N2430), .CP(clk), 
        .Q(inner_first_stage_data_reg[313]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_312_ ( .D(N2429), .CP(clk), 
        .Q(inner_first_stage_data_reg[312]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_311_ ( .D(N2428), .CP(clk), 
        .Q(inner_first_stage_data_reg[311]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_310_ ( .D(N2427), .CP(clk), 
        .Q(inner_first_stage_data_reg[310]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_309_ ( .D(N2426), .CP(clk), 
        .Q(inner_first_stage_data_reg[309]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_308_ ( .D(N2425), .CP(clk), 
        .Q(inner_first_stage_data_reg[308]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_307_ ( .D(N2424), .CP(clk), 
        .Q(inner_first_stage_data_reg[307]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_306_ ( .D(N2423), .CP(clk), 
        .Q(inner_first_stage_data_reg[306]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_305_ ( .D(N2422), .CP(clk), 
        .Q(inner_first_stage_data_reg[305]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_304_ ( .D(N2421), .CP(clk), 
        .Q(inner_first_stage_data_reg[304]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_303_ ( .D(N2420), .CP(clk), 
        .Q(inner_first_stage_data_reg[303]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_302_ ( .D(N2419), .CP(clk), 
        .Q(inner_first_stage_data_reg[302]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_301_ ( .D(N2418), .CP(clk), 
        .Q(inner_first_stage_data_reg[301]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_300_ ( .D(N2417), .CP(clk), 
        .Q(inner_first_stage_data_reg[300]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_299_ ( .D(N2416), .CP(clk), 
        .Q(inner_first_stage_data_reg[299]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_298_ ( .D(N2415), .CP(clk), 
        .Q(inner_first_stage_data_reg[298]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_297_ ( .D(N2414), .CP(clk), 
        .Q(inner_first_stage_data_reg[297]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_296_ ( .D(N2413), .CP(clk), 
        .Q(inner_first_stage_data_reg[296]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_295_ ( .D(N2412), .CP(clk), 
        .Q(inner_first_stage_data_reg[295]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_294_ ( .D(N2411), .CP(clk), 
        .Q(inner_first_stage_data_reg[294]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_293_ ( .D(N2410), .CP(clk), 
        .Q(inner_first_stage_data_reg[293]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_292_ ( .D(N2409), .CP(clk), 
        .Q(inner_first_stage_data_reg[292]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_291_ ( .D(N2408), .CP(clk), 
        .Q(inner_first_stage_data_reg[291]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_290_ ( .D(N2407), .CP(clk), 
        .Q(inner_first_stage_data_reg[290]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_289_ ( .D(N2406), .CP(clk), 
        .Q(inner_first_stage_data_reg[289]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_288_ ( .D(N2405), .CP(clk), 
        .Q(inner_first_stage_data_reg[288]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_10_ ( .D(N2492), .CP(clk), 
        .Q(inner_first_stage_valid_reg[10]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_351_ ( .D(N2524), .CP(clk), 
        .Q(inner_first_stage_data_reg[351]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_350_ ( .D(N2523), .CP(clk), 
        .Q(inner_first_stage_data_reg[350]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_349_ ( .D(N2522), .CP(clk), 
        .Q(inner_first_stage_data_reg[349]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_348_ ( .D(N2521), .CP(clk), 
        .Q(inner_first_stage_data_reg[348]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_347_ ( .D(N2520), .CP(clk), 
        .Q(inner_first_stage_data_reg[347]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_346_ ( .D(N2519), .CP(clk), 
        .Q(inner_first_stage_data_reg[346]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_345_ ( .D(N2518), .CP(clk), 
        .Q(inner_first_stage_data_reg[345]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_344_ ( .D(N2517), .CP(clk), 
        .Q(inner_first_stage_data_reg[344]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_343_ ( .D(N2516), .CP(clk), 
        .Q(inner_first_stage_data_reg[343]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_342_ ( .D(N2515), .CP(clk), 
        .Q(inner_first_stage_data_reg[342]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_341_ ( .D(N2514), .CP(clk), 
        .Q(inner_first_stage_data_reg[341]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_340_ ( .D(N2513), .CP(clk), 
        .Q(inner_first_stage_data_reg[340]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_339_ ( .D(N2512), .CP(clk), 
        .Q(inner_first_stage_data_reg[339]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_338_ ( .D(N2511), .CP(clk), 
        .Q(inner_first_stage_data_reg[338]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_337_ ( .D(N2510), .CP(clk), 
        .Q(inner_first_stage_data_reg[337]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_336_ ( .D(N2509), .CP(clk), 
        .Q(inner_first_stage_data_reg[336]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_335_ ( .D(N2508), .CP(clk), 
        .Q(inner_first_stage_data_reg[335]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_334_ ( .D(N2507), .CP(clk), 
        .Q(inner_first_stage_data_reg[334]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_333_ ( .D(N2506), .CP(clk), 
        .Q(inner_first_stage_data_reg[333]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_332_ ( .D(N2505), .CP(clk), 
        .Q(inner_first_stage_data_reg[332]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_331_ ( .D(N2504), .CP(clk), 
        .Q(inner_first_stage_data_reg[331]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_330_ ( .D(N2503), .CP(clk), 
        .Q(inner_first_stage_data_reg[330]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_329_ ( .D(N2502), .CP(clk), 
        .Q(inner_first_stage_data_reg[329]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_328_ ( .D(N2501), .CP(clk), 
        .Q(inner_first_stage_data_reg[328]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_327_ ( .D(N2500), .CP(clk), 
        .Q(inner_first_stage_data_reg[327]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_326_ ( .D(N2499), .CP(clk), 
        .Q(inner_first_stage_data_reg[326]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_325_ ( .D(N2498), .CP(clk), 
        .Q(inner_first_stage_data_reg[325]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_324_ ( .D(N2497), .CP(clk), 
        .Q(inner_first_stage_data_reg[324]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_323_ ( .D(N2496), .CP(clk), 
        .Q(inner_first_stage_data_reg[323]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_322_ ( .D(N2495), .CP(clk), 
        .Q(inner_first_stage_data_reg[322]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_321_ ( .D(N2494), .CP(clk), 
        .Q(inner_first_stage_data_reg[321]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_320_ ( .D(N2493), .CP(clk), 
        .Q(inner_first_stage_data_reg[320]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_11_ ( .D(N2580), .CP(clk), 
        .Q(inner_first_stage_valid_reg[11]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_383_ ( .D(N2612), .CP(clk), 
        .Q(inner_first_stage_data_reg[383]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_382_ ( .D(N2611), .CP(clk), 
        .Q(inner_first_stage_data_reg[382]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_381_ ( .D(N2610), .CP(clk), 
        .Q(inner_first_stage_data_reg[381]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_380_ ( .D(N2609), .CP(clk), 
        .Q(inner_first_stage_data_reg[380]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_379_ ( .D(N2608), .CP(clk), 
        .Q(inner_first_stage_data_reg[379]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_378_ ( .D(N2607), .CP(clk), 
        .Q(inner_first_stage_data_reg[378]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_377_ ( .D(N2606), .CP(clk), 
        .Q(inner_first_stage_data_reg[377]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_376_ ( .D(N2605), .CP(clk), 
        .Q(inner_first_stage_data_reg[376]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_375_ ( .D(N2604), .CP(clk), 
        .Q(inner_first_stage_data_reg[375]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_374_ ( .D(N2603), .CP(clk), 
        .Q(inner_first_stage_data_reg[374]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_373_ ( .D(N2602), .CP(clk), 
        .Q(inner_first_stage_data_reg[373]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_372_ ( .D(N2601), .CP(clk), 
        .Q(inner_first_stage_data_reg[372]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_371_ ( .D(N2600), .CP(clk), 
        .Q(inner_first_stage_data_reg[371]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_370_ ( .D(N2599), .CP(clk), 
        .Q(inner_first_stage_data_reg[370]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_369_ ( .D(N2598), .CP(clk), 
        .Q(inner_first_stage_data_reg[369]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_368_ ( .D(N2597), .CP(clk), 
        .Q(inner_first_stage_data_reg[368]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_367_ ( .D(N2596), .CP(clk), 
        .Q(inner_first_stage_data_reg[367]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_366_ ( .D(N2595), .CP(clk), 
        .Q(inner_first_stage_data_reg[366]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_365_ ( .D(N2594), .CP(clk), 
        .Q(inner_first_stage_data_reg[365]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_364_ ( .D(N2593), .CP(clk), 
        .Q(inner_first_stage_data_reg[364]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_363_ ( .D(N2592), .CP(clk), 
        .Q(inner_first_stage_data_reg[363]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_362_ ( .D(N2591), .CP(clk), 
        .Q(inner_first_stage_data_reg[362]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_361_ ( .D(N2590), .CP(clk), 
        .Q(inner_first_stage_data_reg[361]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_360_ ( .D(N2589), .CP(clk), 
        .Q(inner_first_stage_data_reg[360]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_359_ ( .D(N2588), .CP(clk), 
        .Q(inner_first_stage_data_reg[359]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_358_ ( .D(N2587), .CP(clk), 
        .Q(inner_first_stage_data_reg[358]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_357_ ( .D(N2586), .CP(clk), 
        .Q(inner_first_stage_data_reg[357]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_356_ ( .D(N2585), .CP(clk), 
        .Q(inner_first_stage_data_reg[356]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_355_ ( .D(N2584), .CP(clk), 
        .Q(inner_first_stage_data_reg[355]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_354_ ( .D(N2583), .CP(clk), 
        .Q(inner_first_stage_data_reg[354]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_353_ ( .D(N2582), .CP(clk), 
        .Q(inner_first_stage_data_reg[353]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_352_ ( .D(N2581), .CP(clk), 
        .Q(inner_first_stage_data_reg[352]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_12_ ( .D(N2668), .CP(clk), 
        .Q(inner_first_stage_valid_reg[12]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_415_ ( .D(N2700), .CP(clk), 
        .Q(inner_first_stage_data_reg[415]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_414_ ( .D(N2699), .CP(clk), 
        .Q(inner_first_stage_data_reg[414]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_413_ ( .D(N2698), .CP(clk), 
        .Q(inner_first_stage_data_reg[413]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_412_ ( .D(N2697), .CP(clk), 
        .Q(inner_first_stage_data_reg[412]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_411_ ( .D(N2696), .CP(clk), 
        .Q(inner_first_stage_data_reg[411]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_410_ ( .D(N2695), .CP(clk), 
        .Q(inner_first_stage_data_reg[410]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_409_ ( .D(N2694), .CP(clk), 
        .Q(inner_first_stage_data_reg[409]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_408_ ( .D(N2693), .CP(clk), 
        .Q(inner_first_stage_data_reg[408]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_407_ ( .D(N2692), .CP(clk), 
        .Q(inner_first_stage_data_reg[407]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_406_ ( .D(N2691), .CP(clk), 
        .Q(inner_first_stage_data_reg[406]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_405_ ( .D(N2690), .CP(clk), 
        .Q(inner_first_stage_data_reg[405]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_404_ ( .D(N2689), .CP(clk), 
        .Q(inner_first_stage_data_reg[404]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_403_ ( .D(N2688), .CP(clk), 
        .Q(inner_first_stage_data_reg[403]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_402_ ( .D(N2687), .CP(clk), 
        .Q(inner_first_stage_data_reg[402]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_401_ ( .D(N2686), .CP(clk), 
        .Q(inner_first_stage_data_reg[401]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_400_ ( .D(N2685), .CP(clk), 
        .Q(inner_first_stage_data_reg[400]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_399_ ( .D(N2684), .CP(clk), 
        .Q(inner_first_stage_data_reg[399]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_398_ ( .D(N2683), .CP(clk), 
        .Q(inner_first_stage_data_reg[398]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_397_ ( .D(N2682), .CP(clk), 
        .Q(inner_first_stage_data_reg[397]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_396_ ( .D(N2681), .CP(clk), 
        .Q(inner_first_stage_data_reg[396]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_395_ ( .D(N2680), .CP(clk), 
        .Q(inner_first_stage_data_reg[395]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_394_ ( .D(N2679), .CP(clk), 
        .Q(inner_first_stage_data_reg[394]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_393_ ( .D(N2678), .CP(clk), 
        .Q(inner_first_stage_data_reg[393]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_392_ ( .D(N2677), .CP(clk), 
        .Q(inner_first_stage_data_reg[392]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_391_ ( .D(N2676), .CP(clk), 
        .Q(inner_first_stage_data_reg[391]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_390_ ( .D(N2675), .CP(clk), 
        .Q(inner_first_stage_data_reg[390]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_389_ ( .D(N2674), .CP(clk), 
        .Q(inner_first_stage_data_reg[389]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_388_ ( .D(N2673), .CP(clk), 
        .Q(inner_first_stage_data_reg[388]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_387_ ( .D(N2672), .CP(clk), 
        .Q(inner_first_stage_data_reg[387]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_386_ ( .D(N2671), .CP(clk), 
        .Q(inner_first_stage_data_reg[386]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_385_ ( .D(N2670), .CP(clk), 
        .Q(inner_first_stage_data_reg[385]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_384_ ( .D(N2669), .CP(clk), 
        .Q(inner_first_stage_data_reg[384]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_13_ ( .D(N2756), .CP(clk), 
        .Q(inner_first_stage_valid_reg[13]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_447_ ( .D(N2788), .CP(clk), 
        .Q(inner_first_stage_data_reg[447]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_446_ ( .D(N2787), .CP(clk), 
        .Q(inner_first_stage_data_reg[446]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_445_ ( .D(N2786), .CP(clk), 
        .Q(inner_first_stage_data_reg[445]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_444_ ( .D(N2785), .CP(clk), 
        .Q(inner_first_stage_data_reg[444]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_443_ ( .D(N2784), .CP(clk), 
        .Q(inner_first_stage_data_reg[443]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_442_ ( .D(N2783), .CP(clk), 
        .Q(inner_first_stage_data_reg[442]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_441_ ( .D(N2782), .CP(clk), 
        .Q(inner_first_stage_data_reg[441]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_440_ ( .D(N2781), .CP(clk), 
        .Q(inner_first_stage_data_reg[440]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_439_ ( .D(N2780), .CP(clk), 
        .Q(inner_first_stage_data_reg[439]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_438_ ( .D(N2779), .CP(clk), 
        .Q(inner_first_stage_data_reg[438]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_437_ ( .D(N2778), .CP(clk), 
        .Q(inner_first_stage_data_reg[437]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_436_ ( .D(N2777), .CP(clk), 
        .Q(inner_first_stage_data_reg[436]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_435_ ( .D(N2776), .CP(clk), 
        .Q(inner_first_stage_data_reg[435]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_434_ ( .D(N2775), .CP(clk), 
        .Q(inner_first_stage_data_reg[434]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_433_ ( .D(N2774), .CP(clk), 
        .Q(inner_first_stage_data_reg[433]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_432_ ( .D(N2773), .CP(clk), 
        .Q(inner_first_stage_data_reg[432]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_431_ ( .D(N2772), .CP(clk), 
        .Q(inner_first_stage_data_reg[431]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_430_ ( .D(N2771), .CP(clk), 
        .Q(inner_first_stage_data_reg[430]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_429_ ( .D(N2770), .CP(clk), 
        .Q(inner_first_stage_data_reg[429]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_428_ ( .D(N2769), .CP(clk), 
        .Q(inner_first_stage_data_reg[428]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_427_ ( .D(N2768), .CP(clk), 
        .Q(inner_first_stage_data_reg[427]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_426_ ( .D(N2767), .CP(clk), 
        .Q(inner_first_stage_data_reg[426]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_425_ ( .D(N2766), .CP(clk), 
        .Q(inner_first_stage_data_reg[425]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_424_ ( .D(N2765), .CP(clk), 
        .Q(inner_first_stage_data_reg[424]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_423_ ( .D(N2764), .CP(clk), 
        .Q(inner_first_stage_data_reg[423]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_422_ ( .D(N2763), .CP(clk), 
        .Q(inner_first_stage_data_reg[422]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_421_ ( .D(N2762), .CP(clk), 
        .Q(inner_first_stage_data_reg[421]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_420_ ( .D(N2761), .CP(clk), 
        .Q(inner_first_stage_data_reg[420]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_419_ ( .D(N2760), .CP(clk), 
        .Q(inner_first_stage_data_reg[419]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_418_ ( .D(N2759), .CP(clk), 
        .Q(inner_first_stage_data_reg[418]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_417_ ( .D(N2758), .CP(clk), 
        .Q(inner_first_stage_data_reg[417]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_416_ ( .D(N2757), .CP(clk), 
        .Q(inner_first_stage_data_reg[416]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_14_ ( .D(N2844), .CP(clk), 
        .Q(inner_first_stage_valid_reg[14]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_479_ ( .D(N2876), .CP(clk), 
        .Q(inner_first_stage_data_reg[479]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_478_ ( .D(N2875), .CP(clk), 
        .Q(inner_first_stage_data_reg[478]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_477_ ( .D(N2874), .CP(clk), 
        .Q(inner_first_stage_data_reg[477]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_476_ ( .D(N2873), .CP(clk), 
        .Q(inner_first_stage_data_reg[476]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_475_ ( .D(N2872), .CP(clk), 
        .Q(inner_first_stage_data_reg[475]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_474_ ( .D(N2871), .CP(clk), 
        .Q(inner_first_stage_data_reg[474]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_473_ ( .D(N2870), .CP(clk), 
        .Q(inner_first_stage_data_reg[473]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_472_ ( .D(N2869), .CP(clk), 
        .Q(inner_first_stage_data_reg[472]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_471_ ( .D(N2868), .CP(clk), 
        .Q(inner_first_stage_data_reg[471]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_470_ ( .D(N2867), .CP(clk), 
        .Q(inner_first_stage_data_reg[470]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_469_ ( .D(N2866), .CP(clk), 
        .Q(inner_first_stage_data_reg[469]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_468_ ( .D(N2865), .CP(clk), 
        .Q(inner_first_stage_data_reg[468]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_467_ ( .D(N2864), .CP(clk), 
        .Q(inner_first_stage_data_reg[467]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_466_ ( .D(N2863), .CP(clk), 
        .Q(inner_first_stage_data_reg[466]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_465_ ( .D(N2862), .CP(clk), 
        .Q(inner_first_stage_data_reg[465]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_464_ ( .D(N2861), .CP(clk), 
        .Q(inner_first_stage_data_reg[464]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_463_ ( .D(N2860), .CP(clk), 
        .Q(inner_first_stage_data_reg[463]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_462_ ( .D(N2859), .CP(clk), 
        .Q(inner_first_stage_data_reg[462]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_461_ ( .D(N2858), .CP(clk), 
        .Q(inner_first_stage_data_reg[461]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_460_ ( .D(N2857), .CP(clk), 
        .Q(inner_first_stage_data_reg[460]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_459_ ( .D(N2856), .CP(clk), 
        .Q(inner_first_stage_data_reg[459]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_458_ ( .D(N2855), .CP(clk), 
        .Q(inner_first_stage_data_reg[458]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_457_ ( .D(N2854), .CP(clk), 
        .Q(inner_first_stage_data_reg[457]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_456_ ( .D(N2853), .CP(clk), 
        .Q(inner_first_stage_data_reg[456]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_455_ ( .D(N2852), .CP(clk), 
        .Q(inner_first_stage_data_reg[455]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_454_ ( .D(N2851), .CP(clk), 
        .Q(inner_first_stage_data_reg[454]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_453_ ( .D(N2850), .CP(clk), 
        .Q(inner_first_stage_data_reg[453]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_452_ ( .D(N2849), .CP(clk), 
        .Q(inner_first_stage_data_reg[452]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_451_ ( .D(N2848), .CP(clk), 
        .Q(inner_first_stage_data_reg[451]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_450_ ( .D(N2847), .CP(clk), 
        .Q(inner_first_stage_data_reg[450]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_449_ ( .D(N2846), .CP(clk), 
        .Q(inner_first_stage_data_reg[449]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_448_ ( .D(N2845), .CP(clk), 
        .Q(inner_first_stage_data_reg[448]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_15_ ( .D(N2932), .CP(clk), 
        .Q(inner_first_stage_valid_reg[15]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_511_ ( .D(N2964), .CP(clk), 
        .Q(inner_first_stage_data_reg[511]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_510_ ( .D(N2963), .CP(clk), 
        .Q(inner_first_stage_data_reg[510]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_509_ ( .D(N2962), .CP(clk), 
        .Q(inner_first_stage_data_reg[509]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_508_ ( .D(N2961), .CP(clk), 
        .Q(inner_first_stage_data_reg[508]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_507_ ( .D(N2960), .CP(clk), 
        .Q(inner_first_stage_data_reg[507]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_506_ ( .D(N2959), .CP(clk), 
        .Q(inner_first_stage_data_reg[506]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_505_ ( .D(N2958), .CP(clk), 
        .Q(inner_first_stage_data_reg[505]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_504_ ( .D(N2957), .CP(clk), 
        .Q(inner_first_stage_data_reg[504]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_503_ ( .D(N2956), .CP(clk), 
        .Q(inner_first_stage_data_reg[503]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_502_ ( .D(N2955), .CP(clk), 
        .Q(inner_first_stage_data_reg[502]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_501_ ( .D(N2954), .CP(clk), 
        .Q(inner_first_stage_data_reg[501]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_500_ ( .D(N2953), .CP(clk), 
        .Q(inner_first_stage_data_reg[500]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_499_ ( .D(N2952), .CP(clk), 
        .Q(inner_first_stage_data_reg[499]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_498_ ( .D(N2951), .CP(clk), 
        .Q(inner_first_stage_data_reg[498]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_497_ ( .D(N2950), .CP(clk), 
        .Q(inner_first_stage_data_reg[497]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_496_ ( .D(N2949), .CP(clk), 
        .Q(inner_first_stage_data_reg[496]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_495_ ( .D(N2948), .CP(clk), 
        .Q(inner_first_stage_data_reg[495]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_494_ ( .D(N2947), .CP(clk), 
        .Q(inner_first_stage_data_reg[494]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_493_ ( .D(N2946), .CP(clk), 
        .Q(inner_first_stage_data_reg[493]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_492_ ( .D(N2945), .CP(clk), 
        .Q(inner_first_stage_data_reg[492]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_491_ ( .D(N2944), .CP(clk), 
        .Q(inner_first_stage_data_reg[491]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_490_ ( .D(N2943), .CP(clk), 
        .Q(inner_first_stage_data_reg[490]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_489_ ( .D(N2942), .CP(clk), 
        .Q(inner_first_stage_data_reg[489]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_488_ ( .D(N2941), .CP(clk), 
        .Q(inner_first_stage_data_reg[488]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_487_ ( .D(N2940), .CP(clk), 
        .Q(inner_first_stage_data_reg[487]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_486_ ( .D(N2939), .CP(clk), 
        .Q(inner_first_stage_data_reg[486]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_485_ ( .D(N2938), .CP(clk), 
        .Q(inner_first_stage_data_reg[485]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_484_ ( .D(N2937), .CP(clk), 
        .Q(inner_first_stage_data_reg[484]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_483_ ( .D(N2936), .CP(clk), 
        .Q(inner_first_stage_data_reg[483]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_482_ ( .D(N2935), .CP(clk), 
        .Q(inner_first_stage_data_reg[482]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_481_ ( .D(N2934), .CP(clk), 
        .Q(inner_first_stage_data_reg[481]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_480_ ( .D(N2933), .CP(clk), 
        .Q(inner_first_stage_data_reg[480]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_16_ ( .D(N3294), .CP(clk), 
        .Q(inner_first_stage_valid_reg[16]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_543_ ( .D(N3326), .CP(clk), 
        .Q(inner_first_stage_data_reg[543]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_542_ ( .D(N3325), .CP(clk), 
        .Q(inner_first_stage_data_reg[542]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_541_ ( .D(N3324), .CP(clk), 
        .Q(inner_first_stage_data_reg[541]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_540_ ( .D(N3323), .CP(clk), 
        .Q(inner_first_stage_data_reg[540]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_539_ ( .D(N3322), .CP(clk), 
        .Q(inner_first_stage_data_reg[539]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_538_ ( .D(N3321), .CP(clk), 
        .Q(inner_first_stage_data_reg[538]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_537_ ( .D(N3320), .CP(clk), 
        .Q(inner_first_stage_data_reg[537]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_536_ ( .D(N3319), .CP(clk), 
        .Q(inner_first_stage_data_reg[536]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_535_ ( .D(N3318), .CP(clk), 
        .Q(inner_first_stage_data_reg[535]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_534_ ( .D(N3317), .CP(clk), 
        .Q(inner_first_stage_data_reg[534]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_533_ ( .D(N3316), .CP(clk), 
        .Q(inner_first_stage_data_reg[533]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_532_ ( .D(N3315), .CP(clk), 
        .Q(inner_first_stage_data_reg[532]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_531_ ( .D(N3314), .CP(clk), 
        .Q(inner_first_stage_data_reg[531]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_530_ ( .D(N3313), .CP(clk), 
        .Q(inner_first_stage_data_reg[530]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_529_ ( .D(N3312), .CP(clk), 
        .Q(inner_first_stage_data_reg[529]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_528_ ( .D(N3311), .CP(clk), 
        .Q(inner_first_stage_data_reg[528]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_527_ ( .D(N3310), .CP(clk), 
        .Q(inner_first_stage_data_reg[527]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_526_ ( .D(N3309), .CP(clk), 
        .Q(inner_first_stage_data_reg[526]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_525_ ( .D(N3308), .CP(clk), 
        .Q(inner_first_stage_data_reg[525]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_524_ ( .D(N3307), .CP(clk), 
        .Q(inner_first_stage_data_reg[524]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_523_ ( .D(N3306), .CP(clk), 
        .Q(inner_first_stage_data_reg[523]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_522_ ( .D(N3305), .CP(clk), 
        .Q(inner_first_stage_data_reg[522]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_521_ ( .D(N3304), .CP(clk), 
        .Q(inner_first_stage_data_reg[521]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_520_ ( .D(N3303), .CP(clk), 
        .Q(inner_first_stage_data_reg[520]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_519_ ( .D(N3302), .CP(clk), 
        .Q(inner_first_stage_data_reg[519]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_518_ ( .D(N3301), .CP(clk), 
        .Q(inner_first_stage_data_reg[518]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_517_ ( .D(N3300), .CP(clk), 
        .Q(inner_first_stage_data_reg[517]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_516_ ( .D(N3299), .CP(clk), 
        .Q(inner_first_stage_data_reg[516]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_515_ ( .D(N3298), .CP(clk), 
        .Q(inner_first_stage_data_reg[515]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_514_ ( .D(N3297), .CP(clk), 
        .Q(inner_first_stage_data_reg[514]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_513_ ( .D(N3296), .CP(clk), 
        .Q(inner_first_stage_data_reg[513]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_512_ ( .D(N3295), .CP(clk), 
        .Q(inner_first_stage_data_reg[512]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_17_ ( .D(N3510), .CP(clk), 
        .Q(inner_first_stage_valid_reg[17]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_575_ ( .D(N3542), .CP(clk), 
        .Q(inner_first_stage_data_reg[575]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_574_ ( .D(N3541), .CP(clk), 
        .Q(inner_first_stage_data_reg[574]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_573_ ( .D(N3540), .CP(clk), 
        .Q(inner_first_stage_data_reg[573]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_572_ ( .D(N3539), .CP(clk), 
        .Q(inner_first_stage_data_reg[572]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_571_ ( .D(N3538), .CP(clk), 
        .Q(inner_first_stage_data_reg[571]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_570_ ( .D(N3537), .CP(clk), 
        .Q(inner_first_stage_data_reg[570]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_569_ ( .D(N3536), .CP(clk), 
        .Q(inner_first_stage_data_reg[569]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_568_ ( .D(N3535), .CP(clk), 
        .Q(inner_first_stage_data_reg[568]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_567_ ( .D(N3534), .CP(clk), 
        .Q(inner_first_stage_data_reg[567]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_566_ ( .D(N3533), .CP(clk), 
        .Q(inner_first_stage_data_reg[566]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_565_ ( .D(N3532), .CP(clk), 
        .Q(inner_first_stage_data_reg[565]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_564_ ( .D(N3531), .CP(clk), 
        .Q(inner_first_stage_data_reg[564]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_563_ ( .D(N3530), .CP(clk), 
        .Q(inner_first_stage_data_reg[563]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_562_ ( .D(N3529), .CP(clk), 
        .Q(inner_first_stage_data_reg[562]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_561_ ( .D(N3528), .CP(clk), 
        .Q(inner_first_stage_data_reg[561]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_560_ ( .D(N3527), .CP(clk), 
        .Q(inner_first_stage_data_reg[560]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_559_ ( .D(N3526), .CP(clk), 
        .Q(inner_first_stage_data_reg[559]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_558_ ( .D(N3525), .CP(clk), 
        .Q(inner_first_stage_data_reg[558]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_557_ ( .D(N3524), .CP(clk), 
        .Q(inner_first_stage_data_reg[557]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_556_ ( .D(N3523), .CP(clk), 
        .Q(inner_first_stage_data_reg[556]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_555_ ( .D(N3522), .CP(clk), 
        .Q(inner_first_stage_data_reg[555]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_554_ ( .D(N3521), .CP(clk), 
        .Q(inner_first_stage_data_reg[554]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_553_ ( .D(N3520), .CP(clk), 
        .Q(inner_first_stage_data_reg[553]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_552_ ( .D(N3519), .CP(clk), 
        .Q(inner_first_stage_data_reg[552]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_551_ ( .D(N3518), .CP(clk), 
        .Q(inner_first_stage_data_reg[551]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_550_ ( .D(N3517), .CP(clk), 
        .Q(inner_first_stage_data_reg[550]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_549_ ( .D(N3516), .CP(clk), 
        .Q(inner_first_stage_data_reg[549]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_548_ ( .D(N3515), .CP(clk), 
        .Q(inner_first_stage_data_reg[548]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_547_ ( .D(N3514), .CP(clk), 
        .Q(inner_first_stage_data_reg[547]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_546_ ( .D(N3513), .CP(clk), 
        .Q(inner_first_stage_data_reg[546]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_545_ ( .D(N3512), .CP(clk), 
        .Q(inner_first_stage_data_reg[545]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_544_ ( .D(N3511), .CP(clk), 
        .Q(inner_first_stage_data_reg[544]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_18_ ( .D(N3726), .CP(clk), 
        .Q(inner_first_stage_valid_reg[18]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_607_ ( .D(N3758), .CP(clk), 
        .Q(inner_first_stage_data_reg[607]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_606_ ( .D(N3757), .CP(clk), 
        .Q(inner_first_stage_data_reg[606]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_605_ ( .D(N3756), .CP(clk), 
        .Q(inner_first_stage_data_reg[605]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_604_ ( .D(N3755), .CP(clk), 
        .Q(inner_first_stage_data_reg[604]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_603_ ( .D(N3754), .CP(clk), 
        .Q(inner_first_stage_data_reg[603]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_602_ ( .D(N3753), .CP(clk), 
        .Q(inner_first_stage_data_reg[602]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_601_ ( .D(N3752), .CP(clk), 
        .Q(inner_first_stage_data_reg[601]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_600_ ( .D(N3751), .CP(clk), 
        .Q(inner_first_stage_data_reg[600]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_599_ ( .D(N3750), .CP(clk), 
        .Q(inner_first_stage_data_reg[599]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_598_ ( .D(N3749), .CP(clk), 
        .Q(inner_first_stage_data_reg[598]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_597_ ( .D(N3748), .CP(clk), 
        .Q(inner_first_stage_data_reg[597]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_596_ ( .D(N3747), .CP(clk), 
        .Q(inner_first_stage_data_reg[596]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_595_ ( .D(N3746), .CP(clk), 
        .Q(inner_first_stage_data_reg[595]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_594_ ( .D(N3745), .CP(clk), 
        .Q(inner_first_stage_data_reg[594]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_593_ ( .D(N3744), .CP(clk), 
        .Q(inner_first_stage_data_reg[593]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_592_ ( .D(N3743), .CP(clk), 
        .Q(inner_first_stage_data_reg[592]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_591_ ( .D(N3742), .CP(clk), 
        .Q(inner_first_stage_data_reg[591]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_590_ ( .D(N3741), .CP(clk), 
        .Q(inner_first_stage_data_reg[590]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_589_ ( .D(N3740), .CP(clk), 
        .Q(inner_first_stage_data_reg[589]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_588_ ( .D(N3739), .CP(clk), 
        .Q(inner_first_stage_data_reg[588]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_587_ ( .D(N3738), .CP(clk), 
        .Q(inner_first_stage_data_reg[587]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_586_ ( .D(N3737), .CP(clk), 
        .Q(inner_first_stage_data_reg[586]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_585_ ( .D(N3736), .CP(clk), 
        .Q(inner_first_stage_data_reg[585]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_584_ ( .D(N3735), .CP(clk), 
        .Q(inner_first_stage_data_reg[584]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_583_ ( .D(N3734), .CP(clk), 
        .Q(inner_first_stage_data_reg[583]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_582_ ( .D(N3733), .CP(clk), 
        .Q(inner_first_stage_data_reg[582]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_581_ ( .D(N3732), .CP(clk), 
        .Q(inner_first_stage_data_reg[581]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_580_ ( .D(N3731), .CP(clk), 
        .Q(inner_first_stage_data_reg[580]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_579_ ( .D(N3730), .CP(clk), 
        .Q(inner_first_stage_data_reg[579]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_578_ ( .D(N3729), .CP(clk), 
        .Q(inner_first_stage_data_reg[578]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_577_ ( .D(N3728), .CP(clk), 
        .Q(inner_first_stage_data_reg[577]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_576_ ( .D(N3727), .CP(clk), 
        .Q(inner_first_stage_data_reg[576]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_19_ ( .D(N3942), .CP(clk), 
        .Q(inner_first_stage_valid_reg[19]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_639_ ( .D(N3974), .CP(clk), 
        .Q(inner_first_stage_data_reg[639]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_638_ ( .D(N3973), .CP(clk), 
        .Q(inner_first_stage_data_reg[638]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_637_ ( .D(N3972), .CP(clk), 
        .Q(inner_first_stage_data_reg[637]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_636_ ( .D(N3971), .CP(clk), 
        .Q(inner_first_stage_data_reg[636]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_635_ ( .D(N3970), .CP(clk), 
        .Q(inner_first_stage_data_reg[635]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_634_ ( .D(N3969), .CP(clk), 
        .Q(inner_first_stage_data_reg[634]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_633_ ( .D(N3968), .CP(clk), 
        .Q(inner_first_stage_data_reg[633]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_632_ ( .D(N3967), .CP(clk), 
        .Q(inner_first_stage_data_reg[632]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_631_ ( .D(N3966), .CP(clk), 
        .Q(inner_first_stage_data_reg[631]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_630_ ( .D(N3965), .CP(clk), 
        .Q(inner_first_stage_data_reg[630]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_629_ ( .D(N3964), .CP(clk), 
        .Q(inner_first_stage_data_reg[629]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_628_ ( .D(N3963), .CP(clk), 
        .Q(inner_first_stage_data_reg[628]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_627_ ( .D(N3962), .CP(clk), 
        .Q(inner_first_stage_data_reg[627]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_626_ ( .D(N3961), .CP(clk), 
        .Q(inner_first_stage_data_reg[626]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_625_ ( .D(N3960), .CP(clk), 
        .Q(inner_first_stage_data_reg[625]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_624_ ( .D(N3959), .CP(clk), 
        .Q(inner_first_stage_data_reg[624]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_623_ ( .D(N3958), .CP(clk), 
        .Q(inner_first_stage_data_reg[623]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_622_ ( .D(N3957), .CP(clk), 
        .Q(inner_first_stage_data_reg[622]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_621_ ( .D(N3956), .CP(clk), 
        .Q(inner_first_stage_data_reg[621]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_620_ ( .D(N3955), .CP(clk), 
        .Q(inner_first_stage_data_reg[620]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_619_ ( .D(N3954), .CP(clk), 
        .Q(inner_first_stage_data_reg[619]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_618_ ( .D(N3953), .CP(clk), 
        .Q(inner_first_stage_data_reg[618]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_617_ ( .D(N3952), .CP(clk), 
        .Q(inner_first_stage_data_reg[617]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_616_ ( .D(N3951), .CP(clk), 
        .Q(inner_first_stage_data_reg[616]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_615_ ( .D(N3950), .CP(clk), 
        .Q(inner_first_stage_data_reg[615]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_614_ ( .D(N3949), .CP(clk), 
        .Q(inner_first_stage_data_reg[614]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_613_ ( .D(N3948), .CP(clk), 
        .Q(inner_first_stage_data_reg[613]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_612_ ( .D(N3947), .CP(clk), 
        .Q(inner_first_stage_data_reg[612]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_611_ ( .D(N3946), .CP(clk), 
        .Q(inner_first_stage_data_reg[611]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_610_ ( .D(N3945), .CP(clk), 
        .Q(inner_first_stage_data_reg[610]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_609_ ( .D(N3944), .CP(clk), 
        .Q(inner_first_stage_data_reg[609]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_608_ ( .D(N3943), .CP(clk), 
        .Q(inner_first_stage_data_reg[608]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_20_ ( .D(N4158), .CP(clk), 
        .Q(inner_first_stage_valid_reg[20]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_671_ ( .D(N4190), .CP(clk), 
        .Q(inner_first_stage_data_reg[671]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_670_ ( .D(N4189), .CP(clk), 
        .Q(inner_first_stage_data_reg[670]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_669_ ( .D(N4188), .CP(clk), 
        .Q(inner_first_stage_data_reg[669]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_668_ ( .D(N4187), .CP(clk), 
        .Q(inner_first_stage_data_reg[668]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_667_ ( .D(N4186), .CP(clk), 
        .Q(inner_first_stage_data_reg[667]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_666_ ( .D(N4185), .CP(clk), 
        .Q(inner_first_stage_data_reg[666]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_665_ ( .D(N4184), .CP(clk), 
        .Q(inner_first_stage_data_reg[665]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_664_ ( .D(N4183), .CP(clk), 
        .Q(inner_first_stage_data_reg[664]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_663_ ( .D(N4182), .CP(clk), 
        .Q(inner_first_stage_data_reg[663]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_662_ ( .D(N4181), .CP(clk), 
        .Q(inner_first_stage_data_reg[662]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_661_ ( .D(N4180), .CP(clk), 
        .Q(inner_first_stage_data_reg[661]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_660_ ( .D(N4179), .CP(clk), 
        .Q(inner_first_stage_data_reg[660]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_659_ ( .D(N4178), .CP(clk), 
        .Q(inner_first_stage_data_reg[659]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_658_ ( .D(N4177), .CP(clk), 
        .Q(inner_first_stage_data_reg[658]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_657_ ( .D(N4176), .CP(clk), 
        .Q(inner_first_stage_data_reg[657]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_656_ ( .D(N4175), .CP(clk), 
        .Q(inner_first_stage_data_reg[656]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_655_ ( .D(N4174), .CP(clk), 
        .Q(inner_first_stage_data_reg[655]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_654_ ( .D(N4173), .CP(clk), 
        .Q(inner_first_stage_data_reg[654]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_653_ ( .D(N4172), .CP(clk), 
        .Q(inner_first_stage_data_reg[653]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_652_ ( .D(N4171), .CP(clk), 
        .Q(inner_first_stage_data_reg[652]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_651_ ( .D(N4170), .CP(clk), 
        .Q(inner_first_stage_data_reg[651]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_650_ ( .D(N4169), .CP(clk), 
        .Q(inner_first_stage_data_reg[650]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_649_ ( .D(N4168), .CP(clk), 
        .Q(inner_first_stage_data_reg[649]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_648_ ( .D(N4167), .CP(clk), 
        .Q(inner_first_stage_data_reg[648]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_647_ ( .D(N4166), .CP(clk), 
        .Q(inner_first_stage_data_reg[647]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_646_ ( .D(N4165), .CP(clk), 
        .Q(inner_first_stage_data_reg[646]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_645_ ( .D(N4164), .CP(clk), 
        .Q(inner_first_stage_data_reg[645]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_644_ ( .D(N4163), .CP(clk), 
        .Q(inner_first_stage_data_reg[644]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_643_ ( .D(N4162), .CP(clk), 
        .Q(inner_first_stage_data_reg[643]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_642_ ( .D(N4161), .CP(clk), 
        .Q(inner_first_stage_data_reg[642]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_641_ ( .D(N4160), .CP(clk), 
        .Q(inner_first_stage_data_reg[641]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_640_ ( .D(N4159), .CP(clk), 
        .Q(inner_first_stage_data_reg[640]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_21_ ( .D(N4374), .CP(clk), 
        .Q(inner_first_stage_valid_reg[21]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_703_ ( .D(N4406), .CP(clk), 
        .Q(inner_first_stage_data_reg[703]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_702_ ( .D(N4405), .CP(clk), 
        .Q(inner_first_stage_data_reg[702]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_701_ ( .D(N4404), .CP(clk), 
        .Q(inner_first_stage_data_reg[701]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_700_ ( .D(N4403), .CP(clk), 
        .Q(inner_first_stage_data_reg[700]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_699_ ( .D(N4402), .CP(clk), 
        .Q(inner_first_stage_data_reg[699]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_698_ ( .D(N4401), .CP(clk), 
        .Q(inner_first_stage_data_reg[698]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_697_ ( .D(N4400), .CP(clk), 
        .Q(inner_first_stage_data_reg[697]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_696_ ( .D(N4399), .CP(clk), 
        .Q(inner_first_stage_data_reg[696]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_695_ ( .D(N4398), .CP(clk), 
        .Q(inner_first_stage_data_reg[695]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_694_ ( .D(N4397), .CP(clk), 
        .Q(inner_first_stage_data_reg[694]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_693_ ( .D(N4396), .CP(clk), 
        .Q(inner_first_stage_data_reg[693]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_692_ ( .D(N4395), .CP(clk), 
        .Q(inner_first_stage_data_reg[692]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_691_ ( .D(N4394), .CP(clk), 
        .Q(inner_first_stage_data_reg[691]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_690_ ( .D(N4393), .CP(clk), 
        .Q(inner_first_stage_data_reg[690]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_689_ ( .D(N4392), .CP(clk), 
        .Q(inner_first_stage_data_reg[689]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_688_ ( .D(N4391), .CP(clk), 
        .Q(inner_first_stage_data_reg[688]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_687_ ( .D(N4390), .CP(clk), 
        .Q(inner_first_stage_data_reg[687]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_686_ ( .D(N4389), .CP(clk), 
        .Q(inner_first_stage_data_reg[686]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_685_ ( .D(N4388), .CP(clk), 
        .Q(inner_first_stage_data_reg[685]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_684_ ( .D(N4387), .CP(clk), 
        .Q(inner_first_stage_data_reg[684]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_683_ ( .D(N4386), .CP(clk), 
        .Q(inner_first_stage_data_reg[683]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_682_ ( .D(N4385), .CP(clk), 
        .Q(inner_first_stage_data_reg[682]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_681_ ( .D(N4384), .CP(clk), 
        .Q(inner_first_stage_data_reg[681]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_680_ ( .D(N4383), .CP(clk), 
        .Q(inner_first_stage_data_reg[680]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_679_ ( .D(N4382), .CP(clk), 
        .Q(inner_first_stage_data_reg[679]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_678_ ( .D(N4381), .CP(clk), 
        .Q(inner_first_stage_data_reg[678]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_677_ ( .D(N4380), .CP(clk), 
        .Q(inner_first_stage_data_reg[677]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_676_ ( .D(N4379), .CP(clk), 
        .Q(inner_first_stage_data_reg[676]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_675_ ( .D(N4378), .CP(clk), 
        .Q(inner_first_stage_data_reg[675]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_674_ ( .D(N4377), .CP(clk), 
        .Q(inner_first_stage_data_reg[674]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_673_ ( .D(N4376), .CP(clk), 
        .Q(inner_first_stage_data_reg[673]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_672_ ( .D(N4375), .CP(clk), 
        .Q(inner_first_stage_data_reg[672]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_22_ ( .D(N4590), .CP(clk), 
        .Q(inner_first_stage_valid_reg[22]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_735_ ( .D(N4622), .CP(clk), 
        .Q(inner_first_stage_data_reg[735]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_734_ ( .D(N4621), .CP(clk), 
        .Q(inner_first_stage_data_reg[734]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_733_ ( .D(N4620), .CP(clk), 
        .Q(inner_first_stage_data_reg[733]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_732_ ( .D(N4619), .CP(clk), 
        .Q(inner_first_stage_data_reg[732]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_731_ ( .D(N4618), .CP(clk), 
        .Q(inner_first_stage_data_reg[731]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_730_ ( .D(N4617), .CP(clk), 
        .Q(inner_first_stage_data_reg[730]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_729_ ( .D(N4616), .CP(clk), 
        .Q(inner_first_stage_data_reg[729]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_728_ ( .D(N4615), .CP(clk), 
        .Q(inner_first_stage_data_reg[728]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_727_ ( .D(N4614), .CP(clk), 
        .Q(inner_first_stage_data_reg[727]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_726_ ( .D(N4613), .CP(clk), 
        .Q(inner_first_stage_data_reg[726]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_725_ ( .D(N4612), .CP(clk), 
        .Q(inner_first_stage_data_reg[725]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_724_ ( .D(N4611), .CP(clk), 
        .Q(inner_first_stage_data_reg[724]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_723_ ( .D(N4610), .CP(clk), 
        .Q(inner_first_stage_data_reg[723]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_722_ ( .D(N4609), .CP(clk), 
        .Q(inner_first_stage_data_reg[722]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_721_ ( .D(N4608), .CP(clk), 
        .Q(inner_first_stage_data_reg[721]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_720_ ( .D(N4607), .CP(clk), 
        .Q(inner_first_stage_data_reg[720]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_719_ ( .D(N4606), .CP(clk), 
        .Q(inner_first_stage_data_reg[719]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_718_ ( .D(N4605), .CP(clk), 
        .Q(inner_first_stage_data_reg[718]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_717_ ( .D(N4604), .CP(clk), 
        .Q(inner_first_stage_data_reg[717]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_716_ ( .D(N4603), .CP(clk), 
        .Q(inner_first_stage_data_reg[716]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_715_ ( .D(N4602), .CP(clk), 
        .Q(inner_first_stage_data_reg[715]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_714_ ( .D(N4601), .CP(clk), 
        .Q(inner_first_stage_data_reg[714]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_713_ ( .D(N4600), .CP(clk), 
        .Q(inner_first_stage_data_reg[713]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_712_ ( .D(N4599), .CP(clk), 
        .Q(inner_first_stage_data_reg[712]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_711_ ( .D(N4598), .CP(clk), 
        .Q(inner_first_stage_data_reg[711]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_710_ ( .D(N4597), .CP(clk), 
        .Q(inner_first_stage_data_reg[710]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_709_ ( .D(N4596), .CP(clk), 
        .Q(inner_first_stage_data_reg[709]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_708_ ( .D(N4595), .CP(clk), 
        .Q(inner_first_stage_data_reg[708]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_707_ ( .D(N4594), .CP(clk), 
        .Q(inner_first_stage_data_reg[707]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_706_ ( .D(N4593), .CP(clk), 
        .Q(inner_first_stage_data_reg[706]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_705_ ( .D(N4592), .CP(clk), 
        .Q(inner_first_stage_data_reg[705]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_704_ ( .D(N4591), .CP(clk), 
        .Q(inner_first_stage_data_reg[704]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_23_ ( .D(N4806), .CP(clk), 
        .Q(inner_first_stage_valid_reg[23]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_767_ ( .D(N4838), .CP(clk), 
        .Q(inner_first_stage_data_reg[767]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_766_ ( .D(N4837), .CP(clk), 
        .Q(inner_first_stage_data_reg[766]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_765_ ( .D(N4836), .CP(clk), 
        .Q(inner_first_stage_data_reg[765]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_764_ ( .D(N4835), .CP(clk), 
        .Q(inner_first_stage_data_reg[764]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_763_ ( .D(N4834), .CP(clk), 
        .Q(inner_first_stage_data_reg[763]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_762_ ( .D(N4833), .CP(clk), 
        .Q(inner_first_stage_data_reg[762]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_761_ ( .D(N4832), .CP(clk), 
        .Q(inner_first_stage_data_reg[761]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_760_ ( .D(N4831), .CP(clk), 
        .Q(inner_first_stage_data_reg[760]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_759_ ( .D(N4830), .CP(clk), 
        .Q(inner_first_stage_data_reg[759]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_758_ ( .D(N4829), .CP(clk), 
        .Q(inner_first_stage_data_reg[758]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_757_ ( .D(N4828), .CP(clk), 
        .Q(inner_first_stage_data_reg[757]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_756_ ( .D(N4827), .CP(clk), 
        .Q(inner_first_stage_data_reg[756]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_755_ ( .D(N4826), .CP(clk), 
        .Q(inner_first_stage_data_reg[755]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_754_ ( .D(N4825), .CP(clk), 
        .Q(inner_first_stage_data_reg[754]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_753_ ( .D(N4824), .CP(clk), 
        .Q(inner_first_stage_data_reg[753]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_752_ ( .D(N4823), .CP(clk), 
        .Q(inner_first_stage_data_reg[752]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_751_ ( .D(N4822), .CP(clk), 
        .Q(inner_first_stage_data_reg[751]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_750_ ( .D(N4821), .CP(clk), 
        .Q(inner_first_stage_data_reg[750]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_749_ ( .D(N4820), .CP(clk), 
        .Q(inner_first_stage_data_reg[749]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_748_ ( .D(N4819), .CP(clk), 
        .Q(inner_first_stage_data_reg[748]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_747_ ( .D(N4818), .CP(clk), 
        .Q(inner_first_stage_data_reg[747]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_746_ ( .D(N4817), .CP(clk), 
        .Q(inner_first_stage_data_reg[746]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_745_ ( .D(N4816), .CP(clk), 
        .Q(inner_first_stage_data_reg[745]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_744_ ( .D(N4815), .CP(clk), 
        .Q(inner_first_stage_data_reg[744]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_743_ ( .D(N4814), .CP(clk), 
        .Q(inner_first_stage_data_reg[743]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_742_ ( .D(N4813), .CP(clk), 
        .Q(inner_first_stage_data_reg[742]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_741_ ( .D(N4812), .CP(clk), 
        .Q(inner_first_stage_data_reg[741]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_740_ ( .D(N4811), .CP(clk), 
        .Q(inner_first_stage_data_reg[740]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_739_ ( .D(N4810), .CP(clk), 
        .Q(inner_first_stage_data_reg[739]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_738_ ( .D(N4809), .CP(clk), 
        .Q(inner_first_stage_data_reg[738]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_737_ ( .D(N4808), .CP(clk), 
        .Q(inner_first_stage_data_reg[737]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_736_ ( .D(N4807), .CP(clk), 
        .Q(inner_first_stage_data_reg[736]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_24_ ( .D(N5040), .CP(clk), 
        .Q(inner_first_stage_valid_reg[24]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_799_ ( .D(N5072), .CP(clk), 
        .Q(inner_first_stage_data_reg[799]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_798_ ( .D(N5071), .CP(clk), 
        .Q(inner_first_stage_data_reg[798]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_797_ ( .D(N5070), .CP(clk), 
        .Q(inner_first_stage_data_reg[797]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_796_ ( .D(N5069), .CP(clk), 
        .Q(inner_first_stage_data_reg[796]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_795_ ( .D(N5068), .CP(clk), 
        .Q(inner_first_stage_data_reg[795]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_794_ ( .D(N5067), .CP(clk), 
        .Q(inner_first_stage_data_reg[794]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_793_ ( .D(N5066), .CP(clk), 
        .Q(inner_first_stage_data_reg[793]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_792_ ( .D(N5065), .CP(clk), 
        .Q(inner_first_stage_data_reg[792]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_791_ ( .D(N5064), .CP(clk), 
        .Q(inner_first_stage_data_reg[791]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_790_ ( .D(N5063), .CP(clk), 
        .Q(inner_first_stage_data_reg[790]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_789_ ( .D(N5062), .CP(clk), 
        .Q(inner_first_stage_data_reg[789]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_788_ ( .D(N5061), .CP(clk), 
        .Q(inner_first_stage_data_reg[788]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_787_ ( .D(N5060), .CP(clk), 
        .Q(inner_first_stage_data_reg[787]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_786_ ( .D(N5059), .CP(clk), 
        .Q(inner_first_stage_data_reg[786]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_785_ ( .D(N5058), .CP(clk), 
        .Q(inner_first_stage_data_reg[785]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_784_ ( .D(N5057), .CP(clk), 
        .Q(inner_first_stage_data_reg[784]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_783_ ( .D(N5056), .CP(clk), 
        .Q(inner_first_stage_data_reg[783]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_782_ ( .D(N5055), .CP(clk), 
        .Q(inner_first_stage_data_reg[782]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_781_ ( .D(N5054), .CP(clk), 
        .Q(inner_first_stage_data_reg[781]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_780_ ( .D(N5053), .CP(clk), 
        .Q(inner_first_stage_data_reg[780]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_779_ ( .D(N5052), .CP(clk), 
        .Q(inner_first_stage_data_reg[779]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_778_ ( .D(N5051), .CP(clk), 
        .Q(inner_first_stage_data_reg[778]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_777_ ( .D(N5050), .CP(clk), 
        .Q(inner_first_stage_data_reg[777]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_776_ ( .D(N5049), .CP(clk), 
        .Q(inner_first_stage_data_reg[776]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_775_ ( .D(N5048), .CP(clk), 
        .Q(inner_first_stage_data_reg[775]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_774_ ( .D(N5047), .CP(clk), 
        .Q(inner_first_stage_data_reg[774]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_773_ ( .D(N5046), .CP(clk), 
        .Q(inner_first_stage_data_reg[773]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_772_ ( .D(N5045), .CP(clk), 
        .Q(inner_first_stage_data_reg[772]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_771_ ( .D(N5044), .CP(clk), 
        .Q(inner_first_stage_data_reg[771]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_770_ ( .D(N5043), .CP(clk), 
        .Q(inner_first_stage_data_reg[770]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_769_ ( .D(N5042), .CP(clk), 
        .Q(inner_first_stage_data_reg[769]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_768_ ( .D(N5041), .CP(clk), 
        .Q(inner_first_stage_data_reg[768]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_25_ ( .D(N5128), .CP(clk), 
        .Q(inner_first_stage_valid_reg[25]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_831_ ( .D(N5160), .CP(clk), 
        .Q(inner_first_stage_data_reg[831]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_830_ ( .D(N5159), .CP(clk), 
        .Q(inner_first_stage_data_reg[830]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_829_ ( .D(N5158), .CP(clk), 
        .Q(inner_first_stage_data_reg[829]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_828_ ( .D(N5157), .CP(clk), 
        .Q(inner_first_stage_data_reg[828]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_827_ ( .D(N5156), .CP(clk), 
        .Q(inner_first_stage_data_reg[827]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_826_ ( .D(N5155), .CP(clk), 
        .Q(inner_first_stage_data_reg[826]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_825_ ( .D(N5154), .CP(clk), 
        .Q(inner_first_stage_data_reg[825]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_824_ ( .D(N5153), .CP(clk), 
        .Q(inner_first_stage_data_reg[824]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_823_ ( .D(N5152), .CP(clk), 
        .Q(inner_first_stage_data_reg[823]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_822_ ( .D(N5151), .CP(clk), 
        .Q(inner_first_stage_data_reg[822]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_821_ ( .D(N5150), .CP(clk), 
        .Q(inner_first_stage_data_reg[821]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_820_ ( .D(N5149), .CP(clk), 
        .Q(inner_first_stage_data_reg[820]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_819_ ( .D(N5148), .CP(clk), 
        .Q(inner_first_stage_data_reg[819]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_818_ ( .D(N5147), .CP(clk), 
        .Q(inner_first_stage_data_reg[818]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_817_ ( .D(N5146), .CP(clk), 
        .Q(inner_first_stage_data_reg[817]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_816_ ( .D(N5145), .CP(clk), 
        .Q(inner_first_stage_data_reg[816]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_815_ ( .D(N5144), .CP(clk), 
        .Q(inner_first_stage_data_reg[815]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_814_ ( .D(N5143), .CP(clk), 
        .Q(inner_first_stage_data_reg[814]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_813_ ( .D(N5142), .CP(clk), 
        .Q(inner_first_stage_data_reg[813]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_812_ ( .D(N5141), .CP(clk), 
        .Q(inner_first_stage_data_reg[812]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_811_ ( .D(N5140), .CP(clk), 
        .Q(inner_first_stage_data_reg[811]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_810_ ( .D(N5139), .CP(clk), 
        .Q(inner_first_stage_data_reg[810]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_809_ ( .D(N5138), .CP(clk), 
        .Q(inner_first_stage_data_reg[809]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_808_ ( .D(N5137), .CP(clk), 
        .Q(inner_first_stage_data_reg[808]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_807_ ( .D(N5136), .CP(clk), 
        .Q(inner_first_stage_data_reg[807]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_806_ ( .D(N5135), .CP(clk), 
        .Q(inner_first_stage_data_reg[806]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_805_ ( .D(N5134), .CP(clk), 
        .Q(inner_first_stage_data_reg[805]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_804_ ( .D(N5133), .CP(clk), 
        .Q(inner_first_stage_data_reg[804]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_803_ ( .D(N5132), .CP(clk), 
        .Q(inner_first_stage_data_reg[803]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_802_ ( .D(N5131), .CP(clk), 
        .Q(inner_first_stage_data_reg[802]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_801_ ( .D(N5130), .CP(clk), 
        .Q(inner_first_stage_data_reg[801]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_800_ ( .D(N5129), .CP(clk), 
        .Q(inner_first_stage_data_reg[800]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_26_ ( .D(N5216), .CP(clk), 
        .Q(inner_first_stage_valid_reg[26]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_863_ ( .D(N5248), .CP(clk), 
        .Q(inner_first_stage_data_reg[863]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_862_ ( .D(N5247), .CP(clk), 
        .Q(inner_first_stage_data_reg[862]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_861_ ( .D(N5246), .CP(clk), 
        .Q(inner_first_stage_data_reg[861]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_860_ ( .D(N5245), .CP(clk), 
        .Q(inner_first_stage_data_reg[860]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_859_ ( .D(N5244), .CP(clk), 
        .Q(inner_first_stage_data_reg[859]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_858_ ( .D(N5243), .CP(clk), 
        .Q(inner_first_stage_data_reg[858]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_857_ ( .D(N5242), .CP(clk), 
        .Q(inner_first_stage_data_reg[857]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_856_ ( .D(N5241), .CP(clk), 
        .Q(inner_first_stage_data_reg[856]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_855_ ( .D(N5240), .CP(clk), 
        .Q(inner_first_stage_data_reg[855]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_854_ ( .D(N5239), .CP(clk), 
        .Q(inner_first_stage_data_reg[854]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_853_ ( .D(N5238), .CP(clk), 
        .Q(inner_first_stage_data_reg[853]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_852_ ( .D(N5237), .CP(clk), 
        .Q(inner_first_stage_data_reg[852]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_851_ ( .D(N5236), .CP(clk), 
        .Q(inner_first_stage_data_reg[851]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_850_ ( .D(N5235), .CP(clk), 
        .Q(inner_first_stage_data_reg[850]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_849_ ( .D(N5234), .CP(clk), 
        .Q(inner_first_stage_data_reg[849]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_848_ ( .D(N5233), .CP(clk), 
        .Q(inner_first_stage_data_reg[848]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_847_ ( .D(N5232), .CP(clk), 
        .Q(inner_first_stage_data_reg[847]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_846_ ( .D(N5231), .CP(clk), 
        .Q(inner_first_stage_data_reg[846]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_845_ ( .D(N5230), .CP(clk), 
        .Q(inner_first_stage_data_reg[845]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_844_ ( .D(N5229), .CP(clk), 
        .Q(inner_first_stage_data_reg[844]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_843_ ( .D(N5228), .CP(clk), 
        .Q(inner_first_stage_data_reg[843]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_842_ ( .D(N5227), .CP(clk), 
        .Q(inner_first_stage_data_reg[842]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_841_ ( .D(N5226), .CP(clk), 
        .Q(inner_first_stage_data_reg[841]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_840_ ( .D(N5225), .CP(clk), 
        .Q(inner_first_stage_data_reg[840]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_839_ ( .D(N5224), .CP(clk), 
        .Q(inner_first_stage_data_reg[839]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_838_ ( .D(N5223), .CP(clk), 
        .Q(inner_first_stage_data_reg[838]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_837_ ( .D(N5222), .CP(clk), 
        .Q(inner_first_stage_data_reg[837]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_836_ ( .D(N5221), .CP(clk), 
        .Q(inner_first_stage_data_reg[836]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_835_ ( .D(N5220), .CP(clk), 
        .Q(inner_first_stage_data_reg[835]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_834_ ( .D(N5219), .CP(clk), 
        .Q(inner_first_stage_data_reg[834]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_833_ ( .D(N5218), .CP(clk), 
        .Q(inner_first_stage_data_reg[833]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_832_ ( .D(N5217), .CP(clk), 
        .Q(inner_first_stage_data_reg[832]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_27_ ( .D(N5304), .CP(clk), 
        .Q(inner_first_stage_valid_reg[27]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_895_ ( .D(N5336), .CP(clk), 
        .Q(inner_first_stage_data_reg[895]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_894_ ( .D(N5335), .CP(clk), 
        .Q(inner_first_stage_data_reg[894]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_893_ ( .D(N5334), .CP(clk), 
        .Q(inner_first_stage_data_reg[893]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_892_ ( .D(N5333), .CP(clk), 
        .Q(inner_first_stage_data_reg[892]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_891_ ( .D(N5332), .CP(clk), 
        .Q(inner_first_stage_data_reg[891]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_890_ ( .D(N5331), .CP(clk), 
        .Q(inner_first_stage_data_reg[890]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_889_ ( .D(N5330), .CP(clk), 
        .Q(inner_first_stage_data_reg[889]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_888_ ( .D(N5329), .CP(clk), 
        .Q(inner_first_stage_data_reg[888]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_887_ ( .D(N5328), .CP(clk), 
        .Q(inner_first_stage_data_reg[887]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_886_ ( .D(N5327), .CP(clk), 
        .Q(inner_first_stage_data_reg[886]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_885_ ( .D(N5326), .CP(clk), 
        .Q(inner_first_stage_data_reg[885]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_884_ ( .D(N5325), .CP(clk), 
        .Q(inner_first_stage_data_reg[884]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_883_ ( .D(N5324), .CP(clk), 
        .Q(inner_first_stage_data_reg[883]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_882_ ( .D(N5323), .CP(clk), 
        .Q(inner_first_stage_data_reg[882]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_881_ ( .D(N5322), .CP(clk), 
        .Q(inner_first_stage_data_reg[881]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_880_ ( .D(N5321), .CP(clk), 
        .Q(inner_first_stage_data_reg[880]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_879_ ( .D(N5320), .CP(clk), 
        .Q(inner_first_stage_data_reg[879]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_878_ ( .D(N5319), .CP(clk), 
        .Q(inner_first_stage_data_reg[878]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_877_ ( .D(N5318), .CP(clk), 
        .Q(inner_first_stage_data_reg[877]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_876_ ( .D(N5317), .CP(clk), 
        .Q(inner_first_stage_data_reg[876]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_875_ ( .D(N5316), .CP(clk), 
        .Q(inner_first_stage_data_reg[875]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_874_ ( .D(N5315), .CP(clk), 
        .Q(inner_first_stage_data_reg[874]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_873_ ( .D(N5314), .CP(clk), 
        .Q(inner_first_stage_data_reg[873]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_872_ ( .D(N5313), .CP(clk), 
        .Q(inner_first_stage_data_reg[872]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_871_ ( .D(N5312), .CP(clk), 
        .Q(inner_first_stage_data_reg[871]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_870_ ( .D(N5311), .CP(clk), 
        .Q(inner_first_stage_data_reg[870]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_869_ ( .D(N5310), .CP(clk), 
        .Q(inner_first_stage_data_reg[869]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_868_ ( .D(N5309), .CP(clk), 
        .Q(inner_first_stage_data_reg[868]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_867_ ( .D(N5308), .CP(clk), 
        .Q(inner_first_stage_data_reg[867]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_866_ ( .D(N5307), .CP(clk), 
        .Q(inner_first_stage_data_reg[866]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_865_ ( .D(N5306), .CP(clk), 
        .Q(inner_first_stage_data_reg[865]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_864_ ( .D(N5305), .CP(clk), 
        .Q(inner_first_stage_data_reg[864]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_28_ ( .D(N5392), .CP(clk), 
        .Q(inner_first_stage_valid_reg[28]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_927_ ( .D(N5424), .CP(clk), 
        .Q(inner_first_stage_data_reg[927]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_926_ ( .D(N5423), .CP(clk), 
        .Q(inner_first_stage_data_reg[926]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_925_ ( .D(N5422), .CP(clk), 
        .Q(inner_first_stage_data_reg[925]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_924_ ( .D(N5421), .CP(clk), 
        .Q(inner_first_stage_data_reg[924]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_923_ ( .D(N5420), .CP(clk), 
        .Q(inner_first_stage_data_reg[923]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_922_ ( .D(N5419), .CP(clk), 
        .Q(inner_first_stage_data_reg[922]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_921_ ( .D(N5418), .CP(clk), 
        .Q(inner_first_stage_data_reg[921]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_920_ ( .D(N5417), .CP(clk), 
        .Q(inner_first_stage_data_reg[920]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_919_ ( .D(N5416), .CP(clk), 
        .Q(inner_first_stage_data_reg[919]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_918_ ( .D(N5415), .CP(clk), 
        .Q(inner_first_stage_data_reg[918]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_917_ ( .D(N5414), .CP(clk), 
        .Q(inner_first_stage_data_reg[917]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_916_ ( .D(N5413), .CP(clk), 
        .Q(inner_first_stage_data_reg[916]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_915_ ( .D(N5412), .CP(clk), 
        .Q(inner_first_stage_data_reg[915]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_914_ ( .D(N5411), .CP(clk), 
        .Q(inner_first_stage_data_reg[914]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_913_ ( .D(N5410), .CP(clk), 
        .Q(inner_first_stage_data_reg[913]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_912_ ( .D(N5409), .CP(clk), 
        .Q(inner_first_stage_data_reg[912]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_911_ ( .D(N5408), .CP(clk), 
        .Q(inner_first_stage_data_reg[911]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_910_ ( .D(N5407), .CP(clk), 
        .Q(inner_first_stage_data_reg[910]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_909_ ( .D(N5406), .CP(clk), 
        .Q(inner_first_stage_data_reg[909]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_908_ ( .D(N5405), .CP(clk), 
        .Q(inner_first_stage_data_reg[908]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_907_ ( .D(N5404), .CP(clk), 
        .Q(inner_first_stage_data_reg[907]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_906_ ( .D(N5403), .CP(clk), 
        .Q(inner_first_stage_data_reg[906]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_905_ ( .D(N5402), .CP(clk), 
        .Q(inner_first_stage_data_reg[905]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_904_ ( .D(N5401), .CP(clk), 
        .Q(inner_first_stage_data_reg[904]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_903_ ( .D(N5400), .CP(clk), 
        .Q(inner_first_stage_data_reg[903]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_902_ ( .D(N5399), .CP(clk), 
        .Q(inner_first_stage_data_reg[902]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_901_ ( .D(N5398), .CP(clk), 
        .Q(inner_first_stage_data_reg[901]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_900_ ( .D(N5397), .CP(clk), 
        .Q(inner_first_stage_data_reg[900]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_899_ ( .D(N5396), .CP(clk), 
        .Q(inner_first_stage_data_reg[899]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_898_ ( .D(N5395), .CP(clk), 
        .Q(inner_first_stage_data_reg[898]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_897_ ( .D(N5394), .CP(clk), 
        .Q(inner_first_stage_data_reg[897]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_896_ ( .D(N5393), .CP(clk), 
        .Q(inner_first_stage_data_reg[896]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_29_ ( .D(N5480), .CP(clk), 
        .Q(inner_first_stage_valid_reg[29]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_959_ ( .D(N5512), .CP(clk), 
        .Q(inner_first_stage_data_reg[959]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_958_ ( .D(N5511), .CP(clk), 
        .Q(inner_first_stage_data_reg[958]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_957_ ( .D(N5510), .CP(clk), 
        .Q(inner_first_stage_data_reg[957]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_956_ ( .D(N5509), .CP(clk), 
        .Q(inner_first_stage_data_reg[956]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_955_ ( .D(N5508), .CP(clk), 
        .Q(inner_first_stage_data_reg[955]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_954_ ( .D(N5507), .CP(clk), 
        .Q(inner_first_stage_data_reg[954]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_953_ ( .D(N5506), .CP(clk), 
        .Q(inner_first_stage_data_reg[953]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_952_ ( .D(N5505), .CP(clk), 
        .Q(inner_first_stage_data_reg[952]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_951_ ( .D(N5504), .CP(clk), 
        .Q(inner_first_stage_data_reg[951]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_950_ ( .D(N5503), .CP(clk), 
        .Q(inner_first_stage_data_reg[950]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_949_ ( .D(N5502), .CP(clk), 
        .Q(inner_first_stage_data_reg[949]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_948_ ( .D(N5501), .CP(clk), 
        .Q(inner_first_stage_data_reg[948]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_947_ ( .D(N5500), .CP(clk), 
        .Q(inner_first_stage_data_reg[947]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_946_ ( .D(N5499), .CP(clk), 
        .Q(inner_first_stage_data_reg[946]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_945_ ( .D(N5498), .CP(clk), 
        .Q(inner_first_stage_data_reg[945]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_944_ ( .D(N5497), .CP(clk), 
        .Q(inner_first_stage_data_reg[944]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_943_ ( .D(N5496), .CP(clk), 
        .Q(inner_first_stage_data_reg[943]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_942_ ( .D(N5495), .CP(clk), 
        .Q(inner_first_stage_data_reg[942]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_941_ ( .D(N5494), .CP(clk), 
        .Q(inner_first_stage_data_reg[941]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_940_ ( .D(N5493), .CP(clk), 
        .Q(inner_first_stage_data_reg[940]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_939_ ( .D(N5492), .CP(clk), 
        .Q(inner_first_stage_data_reg[939]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_938_ ( .D(N5491), .CP(clk), 
        .Q(inner_first_stage_data_reg[938]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_937_ ( .D(N5490), .CP(clk), 
        .Q(inner_first_stage_data_reg[937]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_936_ ( .D(N5489), .CP(clk), 
        .Q(inner_first_stage_data_reg[936]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_935_ ( .D(N5488), .CP(clk), 
        .Q(inner_first_stage_data_reg[935]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_934_ ( .D(N5487), .CP(clk), 
        .Q(inner_first_stage_data_reg[934]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_933_ ( .D(N5486), .CP(clk), 
        .Q(inner_first_stage_data_reg[933]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_932_ ( .D(N5485), .CP(clk), 
        .Q(inner_first_stage_data_reg[932]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_931_ ( .D(N5484), .CP(clk), 
        .Q(inner_first_stage_data_reg[931]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_930_ ( .D(N5483), .CP(clk), 
        .Q(inner_first_stage_data_reg[930]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_929_ ( .D(N5482), .CP(clk), 
        .Q(inner_first_stage_data_reg[929]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_928_ ( .D(N5481), .CP(clk), 
        .Q(inner_first_stage_data_reg[928]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_30_ ( .D(N5568), .CP(clk), 
        .Q(inner_first_stage_valid_reg[30]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_991_ ( .D(N5600), .CP(clk), 
        .Q(inner_first_stage_data_reg[991]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_990_ ( .D(N5599), .CP(clk), 
        .Q(inner_first_stage_data_reg[990]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_989_ ( .D(N5598), .CP(clk), 
        .Q(inner_first_stage_data_reg[989]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_988_ ( .D(N5597), .CP(clk), 
        .Q(inner_first_stage_data_reg[988]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_987_ ( .D(N5596), .CP(clk), 
        .Q(inner_first_stage_data_reg[987]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_986_ ( .D(N5595), .CP(clk), 
        .Q(inner_first_stage_data_reg[986]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_985_ ( .D(N5594), .CP(clk), 
        .Q(inner_first_stage_data_reg[985]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_984_ ( .D(N5593), .CP(clk), 
        .Q(inner_first_stage_data_reg[984]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_983_ ( .D(N5592), .CP(clk), 
        .Q(inner_first_stage_data_reg[983]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_982_ ( .D(N5591), .CP(clk), 
        .Q(inner_first_stage_data_reg[982]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_981_ ( .D(N5590), .CP(clk), 
        .Q(inner_first_stage_data_reg[981]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_980_ ( .D(N5589), .CP(clk), 
        .Q(inner_first_stage_data_reg[980]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_979_ ( .D(N5588), .CP(clk), 
        .Q(inner_first_stage_data_reg[979]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_978_ ( .D(N5587), .CP(clk), 
        .Q(inner_first_stage_data_reg[978]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_977_ ( .D(N5586), .CP(clk), 
        .Q(inner_first_stage_data_reg[977]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_976_ ( .D(N5585), .CP(clk), 
        .Q(inner_first_stage_data_reg[976]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_975_ ( .D(N5584), .CP(clk), 
        .Q(inner_first_stage_data_reg[975]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_974_ ( .D(N5583), .CP(clk), 
        .Q(inner_first_stage_data_reg[974]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_973_ ( .D(N5582), .CP(clk), 
        .Q(inner_first_stage_data_reg[973]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_972_ ( .D(N5581), .CP(clk), 
        .Q(inner_first_stage_data_reg[972]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_971_ ( .D(N5580), .CP(clk), 
        .Q(inner_first_stage_data_reg[971]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_970_ ( .D(N5579), .CP(clk), 
        .Q(inner_first_stage_data_reg[970]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_969_ ( .D(N5578), .CP(clk), 
        .Q(inner_first_stage_data_reg[969]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_968_ ( .D(N5577), .CP(clk), 
        .Q(inner_first_stage_data_reg[968]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_967_ ( .D(N5576), .CP(clk), 
        .Q(inner_first_stage_data_reg[967]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_966_ ( .D(N5575), .CP(clk), 
        .Q(inner_first_stage_data_reg[966]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_965_ ( .D(N5574), .CP(clk), 
        .Q(inner_first_stage_data_reg[965]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_964_ ( .D(N5573), .CP(clk), 
        .Q(inner_first_stage_data_reg[964]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_963_ ( .D(N5572), .CP(clk), 
        .Q(inner_first_stage_data_reg[963]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_962_ ( .D(N5571), .CP(clk), 
        .Q(inner_first_stage_data_reg[962]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_961_ ( .D(N5570), .CP(clk), 
        .Q(inner_first_stage_data_reg[961]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_960_ ( .D(N5569), .CP(clk), 
        .Q(inner_first_stage_data_reg[960]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_31_ ( .D(N5656), .CP(clk), 
        .Q(inner_first_stage_valid_reg[31]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1023_ ( .D(N5688), .CP(clk), 
        .Q(inner_first_stage_data_reg[1023]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1022_ ( .D(N5687), .CP(clk), 
        .Q(inner_first_stage_data_reg[1022]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1021_ ( .D(N5686), .CP(clk), 
        .Q(inner_first_stage_data_reg[1021]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1020_ ( .D(N5685), .CP(clk), 
        .Q(inner_first_stage_data_reg[1020]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1019_ ( .D(N5684), .CP(clk), 
        .Q(inner_first_stage_data_reg[1019]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1018_ ( .D(N5683), .CP(clk), 
        .Q(inner_first_stage_data_reg[1018]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1017_ ( .D(N5682), .CP(clk), 
        .Q(inner_first_stage_data_reg[1017]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1016_ ( .D(N5681), .CP(clk), 
        .Q(inner_first_stage_data_reg[1016]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1015_ ( .D(N5680), .CP(clk), 
        .Q(inner_first_stage_data_reg[1015]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1014_ ( .D(N5679), .CP(clk), 
        .Q(inner_first_stage_data_reg[1014]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1013_ ( .D(N5678), .CP(clk), 
        .Q(inner_first_stage_data_reg[1013]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1012_ ( .D(N5677), .CP(clk), 
        .Q(inner_first_stage_data_reg[1012]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1011_ ( .D(N5676), .CP(clk), 
        .Q(inner_first_stage_data_reg[1011]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1010_ ( .D(N5675), .CP(clk), 
        .Q(inner_first_stage_data_reg[1010]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1009_ ( .D(N5674), .CP(clk), 
        .Q(inner_first_stage_data_reg[1009]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1008_ ( .D(N5673), .CP(clk), 
        .Q(inner_first_stage_data_reg[1008]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1007_ ( .D(N5672), .CP(clk), 
        .Q(inner_first_stage_data_reg[1007]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1006_ ( .D(N5671), .CP(clk), 
        .Q(inner_first_stage_data_reg[1006]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1005_ ( .D(N5670), .CP(clk), 
        .Q(inner_first_stage_data_reg[1005]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1004_ ( .D(N5669), .CP(clk), 
        .Q(inner_first_stage_data_reg[1004]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1003_ ( .D(N5668), .CP(clk), 
        .Q(inner_first_stage_data_reg[1003]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1002_ ( .D(N5667), .CP(clk), 
        .Q(inner_first_stage_data_reg[1002]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1001_ ( .D(N5666), .CP(clk), 
        .Q(inner_first_stage_data_reg[1001]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1000_ ( .D(N5665), .CP(clk), 
        .Q(inner_first_stage_data_reg[1000]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_999_ ( .D(N5664), .CP(clk), 
        .Q(inner_first_stage_data_reg[999]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_998_ ( .D(N5663), .CP(clk), 
        .Q(inner_first_stage_data_reg[998]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_997_ ( .D(N5662), .CP(clk), 
        .Q(inner_first_stage_data_reg[997]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_996_ ( .D(N5661), .CP(clk), 
        .Q(inner_first_stage_data_reg[996]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_995_ ( .D(N5660), .CP(clk), 
        .Q(inner_first_stage_data_reg[995]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_994_ ( .D(N5659), .CP(clk), 
        .Q(inner_first_stage_data_reg[994]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_993_ ( .D(N5658), .CP(clk), 
        .Q(inner_first_stage_data_reg[993]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_992_ ( .D(N5657), .CP(clk), 
        .Q(inner_first_stage_data_reg[992]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_32_ ( .D(N6018), .CP(clk), 
        .Q(inner_first_stage_valid_reg[32]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1055_ ( .D(N6050), .CP(clk), 
        .Q(inner_first_stage_data_reg[1055]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1054_ ( .D(N6049), .CP(clk), 
        .Q(inner_first_stage_data_reg[1054]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1053_ ( .D(N6048), .CP(clk), 
        .Q(inner_first_stage_data_reg[1053]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1052_ ( .D(N6047), .CP(clk), 
        .Q(inner_first_stage_data_reg[1052]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1051_ ( .D(N6046), .CP(clk), 
        .Q(inner_first_stage_data_reg[1051]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1050_ ( .D(N6045), .CP(clk), 
        .Q(inner_first_stage_data_reg[1050]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1049_ ( .D(N6044), .CP(clk), 
        .Q(inner_first_stage_data_reg[1049]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1048_ ( .D(N6043), .CP(clk), 
        .Q(inner_first_stage_data_reg[1048]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1047_ ( .D(N6042), .CP(clk), 
        .Q(inner_first_stage_data_reg[1047]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1046_ ( .D(N6041), .CP(clk), 
        .Q(inner_first_stage_data_reg[1046]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1045_ ( .D(N6040), .CP(clk), 
        .Q(inner_first_stage_data_reg[1045]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1044_ ( .D(N6039), .CP(clk), 
        .Q(inner_first_stage_data_reg[1044]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1043_ ( .D(N6038), .CP(clk), 
        .Q(inner_first_stage_data_reg[1043]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1042_ ( .D(N6037), .CP(clk), 
        .Q(inner_first_stage_data_reg[1042]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1041_ ( .D(N6036), .CP(clk), 
        .Q(inner_first_stage_data_reg[1041]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1040_ ( .D(N6035), .CP(clk), 
        .Q(inner_first_stage_data_reg[1040]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1039_ ( .D(N6034), .CP(clk), 
        .Q(inner_first_stage_data_reg[1039]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1038_ ( .D(N6033), .CP(clk), 
        .Q(inner_first_stage_data_reg[1038]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1037_ ( .D(N6032), .CP(clk), 
        .Q(inner_first_stage_data_reg[1037]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1036_ ( .D(N6031), .CP(clk), 
        .Q(inner_first_stage_data_reg[1036]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1035_ ( .D(N6030), .CP(clk), 
        .Q(inner_first_stage_data_reg[1035]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1034_ ( .D(N6029), .CP(clk), 
        .Q(inner_first_stage_data_reg[1034]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1033_ ( .D(N6028), .CP(clk), 
        .Q(inner_first_stage_data_reg[1033]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1032_ ( .D(N6027), .CP(clk), 
        .Q(inner_first_stage_data_reg[1032]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1031_ ( .D(N6026), .CP(clk), 
        .Q(inner_first_stage_data_reg[1031]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1030_ ( .D(N6025), .CP(clk), 
        .Q(inner_first_stage_data_reg[1030]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1029_ ( .D(N6024), .CP(clk), 
        .Q(inner_first_stage_data_reg[1029]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1028_ ( .D(N6023), .CP(clk), 
        .Q(inner_first_stage_data_reg[1028]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1027_ ( .D(N6022), .CP(clk), 
        .Q(inner_first_stage_data_reg[1027]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1026_ ( .D(N6021), .CP(clk), 
        .Q(inner_first_stage_data_reg[1026]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1025_ ( .D(N6020), .CP(clk), 
        .Q(inner_first_stage_data_reg[1025]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1024_ ( .D(N6019), .CP(clk), 
        .Q(inner_first_stage_data_reg[1024]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_33_ ( .D(N6234), .CP(clk), 
        .Q(inner_first_stage_valid_reg[33]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1087_ ( .D(N6266), .CP(clk), 
        .Q(inner_first_stage_data_reg[1087]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1086_ ( .D(N6265), .CP(clk), 
        .Q(inner_first_stage_data_reg[1086]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1085_ ( .D(N6264), .CP(clk), 
        .Q(inner_first_stage_data_reg[1085]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1084_ ( .D(N6263), .CP(clk), 
        .Q(inner_first_stage_data_reg[1084]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1083_ ( .D(N6262), .CP(clk), 
        .Q(inner_first_stage_data_reg[1083]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1082_ ( .D(N6261), .CP(clk), 
        .Q(inner_first_stage_data_reg[1082]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1081_ ( .D(N6260), .CP(clk), 
        .Q(inner_first_stage_data_reg[1081]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1080_ ( .D(N6259), .CP(clk), 
        .Q(inner_first_stage_data_reg[1080]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1079_ ( .D(N6258), .CP(clk), 
        .Q(inner_first_stage_data_reg[1079]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1078_ ( .D(N6257), .CP(clk), 
        .Q(inner_first_stage_data_reg[1078]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1077_ ( .D(N6256), .CP(clk), 
        .Q(inner_first_stage_data_reg[1077]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1076_ ( .D(N6255), .CP(clk), 
        .Q(inner_first_stage_data_reg[1076]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1075_ ( .D(N6254), .CP(clk), 
        .Q(inner_first_stage_data_reg[1075]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1074_ ( .D(N6253), .CP(clk), 
        .Q(inner_first_stage_data_reg[1074]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1073_ ( .D(N6252), .CP(clk), 
        .Q(inner_first_stage_data_reg[1073]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1072_ ( .D(N6251), .CP(clk), 
        .Q(inner_first_stage_data_reg[1072]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1071_ ( .D(N6250), .CP(clk), 
        .Q(inner_first_stage_data_reg[1071]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1070_ ( .D(N6249), .CP(clk), 
        .Q(inner_first_stage_data_reg[1070]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1069_ ( .D(N6248), .CP(clk), 
        .Q(inner_first_stage_data_reg[1069]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1068_ ( .D(N6247), .CP(clk), 
        .Q(inner_first_stage_data_reg[1068]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1067_ ( .D(N6246), .CP(clk), 
        .Q(inner_first_stage_data_reg[1067]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1066_ ( .D(N6245), .CP(clk), 
        .Q(inner_first_stage_data_reg[1066]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1065_ ( .D(N6244), .CP(clk), 
        .Q(inner_first_stage_data_reg[1065]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1064_ ( .D(N6243), .CP(clk), 
        .Q(inner_first_stage_data_reg[1064]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1063_ ( .D(N6242), .CP(clk), 
        .Q(inner_first_stage_data_reg[1063]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1062_ ( .D(N6241), .CP(clk), 
        .Q(inner_first_stage_data_reg[1062]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1061_ ( .D(N6240), .CP(clk), 
        .Q(inner_first_stage_data_reg[1061]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1060_ ( .D(N6239), .CP(clk), 
        .Q(inner_first_stage_data_reg[1060]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1059_ ( .D(N6238), .CP(clk), 
        .Q(inner_first_stage_data_reg[1059]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1058_ ( .D(N6237), .CP(clk), 
        .Q(inner_first_stage_data_reg[1058]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1057_ ( .D(N6236), .CP(clk), 
        .Q(inner_first_stage_data_reg[1057]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1056_ ( .D(N6235), .CP(clk), 
        .Q(inner_first_stage_data_reg[1056]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_34_ ( .D(N6450), .CP(clk), 
        .Q(inner_first_stage_valid_reg[34]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1119_ ( .D(N6482), .CP(clk), 
        .Q(inner_first_stage_data_reg[1119]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1118_ ( .D(N6481), .CP(clk), 
        .Q(inner_first_stage_data_reg[1118]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1117_ ( .D(N6480), .CP(clk), 
        .Q(inner_first_stage_data_reg[1117]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1116_ ( .D(N6479), .CP(clk), 
        .Q(inner_first_stage_data_reg[1116]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1115_ ( .D(N6478), .CP(clk), 
        .Q(inner_first_stage_data_reg[1115]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1114_ ( .D(N6477), .CP(clk), 
        .Q(inner_first_stage_data_reg[1114]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1113_ ( .D(N6476), .CP(clk), 
        .Q(inner_first_stage_data_reg[1113]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1112_ ( .D(N6475), .CP(clk), 
        .Q(inner_first_stage_data_reg[1112]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1111_ ( .D(N6474), .CP(clk), 
        .Q(inner_first_stage_data_reg[1111]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1110_ ( .D(N6473), .CP(clk), 
        .Q(inner_first_stage_data_reg[1110]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1109_ ( .D(N6472), .CP(clk), 
        .Q(inner_first_stage_data_reg[1109]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1108_ ( .D(N6471), .CP(clk), 
        .Q(inner_first_stage_data_reg[1108]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1107_ ( .D(N6470), .CP(clk), 
        .Q(inner_first_stage_data_reg[1107]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1106_ ( .D(N6469), .CP(clk), 
        .Q(inner_first_stage_data_reg[1106]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1105_ ( .D(N6468), .CP(clk), 
        .Q(inner_first_stage_data_reg[1105]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1104_ ( .D(N6467), .CP(clk), 
        .Q(inner_first_stage_data_reg[1104]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1103_ ( .D(N6466), .CP(clk), 
        .Q(inner_first_stage_data_reg[1103]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1102_ ( .D(N6465), .CP(clk), 
        .Q(inner_first_stage_data_reg[1102]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1101_ ( .D(N6464), .CP(clk), 
        .Q(inner_first_stage_data_reg[1101]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1100_ ( .D(N6463), .CP(clk), 
        .Q(inner_first_stage_data_reg[1100]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1099_ ( .D(N6462), .CP(clk), 
        .Q(inner_first_stage_data_reg[1099]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1098_ ( .D(N6461), .CP(clk), 
        .Q(inner_first_stage_data_reg[1098]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1097_ ( .D(N6460), .CP(clk), 
        .Q(inner_first_stage_data_reg[1097]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1096_ ( .D(N6459), .CP(clk), 
        .Q(inner_first_stage_data_reg[1096]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1095_ ( .D(N6458), .CP(clk), 
        .Q(inner_first_stage_data_reg[1095]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1094_ ( .D(N6457), .CP(clk), 
        .Q(inner_first_stage_data_reg[1094]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1093_ ( .D(N6456), .CP(clk), 
        .Q(inner_first_stage_data_reg[1093]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1092_ ( .D(N6455), .CP(clk), 
        .Q(inner_first_stage_data_reg[1092]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1091_ ( .D(N6454), .CP(clk), 
        .Q(inner_first_stage_data_reg[1091]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1090_ ( .D(N6453), .CP(clk), 
        .Q(inner_first_stage_data_reg[1090]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1089_ ( .D(N6452), .CP(clk), 
        .Q(inner_first_stage_data_reg[1089]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1088_ ( .D(N6451), .CP(clk), 
        .Q(inner_first_stage_data_reg[1088]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_35_ ( .D(N6666), .CP(clk), 
        .Q(inner_first_stage_valid_reg[35]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1151_ ( .D(N6698), .CP(clk), 
        .Q(inner_first_stage_data_reg[1151]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1150_ ( .D(N6697), .CP(clk), 
        .Q(inner_first_stage_data_reg[1150]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1149_ ( .D(N6696), .CP(clk), 
        .Q(inner_first_stage_data_reg[1149]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1148_ ( .D(N6695), .CP(clk), 
        .Q(inner_first_stage_data_reg[1148]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1147_ ( .D(N6694), .CP(clk), 
        .Q(inner_first_stage_data_reg[1147]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1146_ ( .D(N6693), .CP(clk), 
        .Q(inner_first_stage_data_reg[1146]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1145_ ( .D(N6692), .CP(clk), 
        .Q(inner_first_stage_data_reg[1145]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1144_ ( .D(N6691), .CP(clk), 
        .Q(inner_first_stage_data_reg[1144]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1143_ ( .D(N6690), .CP(clk), 
        .Q(inner_first_stage_data_reg[1143]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1142_ ( .D(N6689), .CP(clk), 
        .Q(inner_first_stage_data_reg[1142]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1141_ ( .D(N6688), .CP(clk), 
        .Q(inner_first_stage_data_reg[1141]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1140_ ( .D(N6687), .CP(clk), 
        .Q(inner_first_stage_data_reg[1140]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1139_ ( .D(N6686), .CP(clk), 
        .Q(inner_first_stage_data_reg[1139]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1138_ ( .D(N6685), .CP(clk), 
        .Q(inner_first_stage_data_reg[1138]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1137_ ( .D(N6684), .CP(clk), 
        .Q(inner_first_stage_data_reg[1137]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1136_ ( .D(N6683), .CP(clk), 
        .Q(inner_first_stage_data_reg[1136]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1135_ ( .D(N6682), .CP(clk), 
        .Q(inner_first_stage_data_reg[1135]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1134_ ( .D(N6681), .CP(clk), 
        .Q(inner_first_stage_data_reg[1134]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1133_ ( .D(N6680), .CP(clk), 
        .Q(inner_first_stage_data_reg[1133]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1132_ ( .D(N6679), .CP(clk), 
        .Q(inner_first_stage_data_reg[1132]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1131_ ( .D(N6678), .CP(clk), 
        .Q(inner_first_stage_data_reg[1131]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1130_ ( .D(N6677), .CP(clk), 
        .Q(inner_first_stage_data_reg[1130]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1129_ ( .D(N6676), .CP(clk), 
        .Q(inner_first_stage_data_reg[1129]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1128_ ( .D(N6675), .CP(clk), 
        .Q(inner_first_stage_data_reg[1128]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1127_ ( .D(N6674), .CP(clk), 
        .Q(inner_first_stage_data_reg[1127]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1126_ ( .D(N6673), .CP(clk), 
        .Q(inner_first_stage_data_reg[1126]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1125_ ( .D(N6672), .CP(clk), 
        .Q(inner_first_stage_data_reg[1125]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1124_ ( .D(N6671), .CP(clk), 
        .Q(inner_first_stage_data_reg[1124]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1123_ ( .D(N6670), .CP(clk), 
        .Q(inner_first_stage_data_reg[1123]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1122_ ( .D(N6669), .CP(clk), 
        .Q(inner_first_stage_data_reg[1122]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1121_ ( .D(N6668), .CP(clk), 
        .Q(inner_first_stage_data_reg[1121]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1120_ ( .D(N6667), .CP(clk), 
        .Q(inner_first_stage_data_reg[1120]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_36_ ( .D(N6882), .CP(clk), 
        .Q(inner_first_stage_valid_reg[36]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1183_ ( .D(N6914), .CP(clk), 
        .Q(inner_first_stage_data_reg[1183]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1182_ ( .D(N6913), .CP(clk), 
        .Q(inner_first_stage_data_reg[1182]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1181_ ( .D(N6912), .CP(clk), 
        .Q(inner_first_stage_data_reg[1181]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1180_ ( .D(N6911), .CP(clk), 
        .Q(inner_first_stage_data_reg[1180]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1179_ ( .D(N6910), .CP(clk), 
        .Q(inner_first_stage_data_reg[1179]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1178_ ( .D(N6909), .CP(clk), 
        .Q(inner_first_stage_data_reg[1178]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1177_ ( .D(N6908), .CP(clk), 
        .Q(inner_first_stage_data_reg[1177]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1176_ ( .D(N6907), .CP(clk), 
        .Q(inner_first_stage_data_reg[1176]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1175_ ( .D(N6906), .CP(clk), 
        .Q(inner_first_stage_data_reg[1175]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1174_ ( .D(N6905), .CP(clk), 
        .Q(inner_first_stage_data_reg[1174]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1173_ ( .D(N6904), .CP(clk), 
        .Q(inner_first_stage_data_reg[1173]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1172_ ( .D(N6903), .CP(clk), 
        .Q(inner_first_stage_data_reg[1172]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1171_ ( .D(N6902), .CP(clk), 
        .Q(inner_first_stage_data_reg[1171]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1170_ ( .D(N6901), .CP(clk), 
        .Q(inner_first_stage_data_reg[1170]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1169_ ( .D(N6900), .CP(clk), 
        .Q(inner_first_stage_data_reg[1169]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1168_ ( .D(N6899), .CP(clk), 
        .Q(inner_first_stage_data_reg[1168]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1167_ ( .D(N6898), .CP(clk), 
        .Q(inner_first_stage_data_reg[1167]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1166_ ( .D(N6897), .CP(clk), 
        .Q(inner_first_stage_data_reg[1166]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1165_ ( .D(N6896), .CP(clk), 
        .Q(inner_first_stage_data_reg[1165]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1164_ ( .D(N6895), .CP(clk), 
        .Q(inner_first_stage_data_reg[1164]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1163_ ( .D(N6894), .CP(clk), 
        .Q(inner_first_stage_data_reg[1163]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1162_ ( .D(N6893), .CP(clk), 
        .Q(inner_first_stage_data_reg[1162]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1161_ ( .D(N6892), .CP(clk), 
        .Q(inner_first_stage_data_reg[1161]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1160_ ( .D(N6891), .CP(clk), 
        .Q(inner_first_stage_data_reg[1160]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1159_ ( .D(N6890), .CP(clk), 
        .Q(inner_first_stage_data_reg[1159]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1158_ ( .D(N6889), .CP(clk), 
        .Q(inner_first_stage_data_reg[1158]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1157_ ( .D(N6888), .CP(clk), 
        .Q(inner_first_stage_data_reg[1157]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1156_ ( .D(N6887), .CP(clk), 
        .Q(inner_first_stage_data_reg[1156]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1155_ ( .D(N6886), .CP(clk), 
        .Q(inner_first_stage_data_reg[1155]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1154_ ( .D(N6885), .CP(clk), 
        .Q(inner_first_stage_data_reg[1154]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1153_ ( .D(N6884), .CP(clk), 
        .Q(inner_first_stage_data_reg[1153]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1152_ ( .D(N6883), .CP(clk), 
        .Q(inner_first_stage_data_reg[1152]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_37_ ( .D(N7098), .CP(clk), 
        .Q(inner_first_stage_valid_reg[37]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1215_ ( .D(N7130), .CP(clk), 
        .Q(inner_first_stage_data_reg[1215]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1214_ ( .D(N7129), .CP(clk), 
        .Q(inner_first_stage_data_reg[1214]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1213_ ( .D(N7128), .CP(clk), 
        .Q(inner_first_stage_data_reg[1213]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1212_ ( .D(N7127), .CP(clk), 
        .Q(inner_first_stage_data_reg[1212]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1211_ ( .D(N7126), .CP(clk), 
        .Q(inner_first_stage_data_reg[1211]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1210_ ( .D(N7125), .CP(clk), 
        .Q(inner_first_stage_data_reg[1210]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1209_ ( .D(N7124), .CP(clk), 
        .Q(inner_first_stage_data_reg[1209]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1208_ ( .D(N7123), .CP(clk), 
        .Q(inner_first_stage_data_reg[1208]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1207_ ( .D(N7122), .CP(clk), 
        .Q(inner_first_stage_data_reg[1207]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1206_ ( .D(N7121), .CP(clk), 
        .Q(inner_first_stage_data_reg[1206]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1205_ ( .D(N7120), .CP(clk), 
        .Q(inner_first_stage_data_reg[1205]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1204_ ( .D(N7119), .CP(clk), 
        .Q(inner_first_stage_data_reg[1204]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1203_ ( .D(N7118), .CP(clk), 
        .Q(inner_first_stage_data_reg[1203]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1202_ ( .D(N7117), .CP(clk), 
        .Q(inner_first_stage_data_reg[1202]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1201_ ( .D(N7116), .CP(clk), 
        .Q(inner_first_stage_data_reg[1201]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1200_ ( .D(N7115), .CP(clk), 
        .Q(inner_first_stage_data_reg[1200]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1199_ ( .D(N7114), .CP(clk), 
        .Q(inner_first_stage_data_reg[1199]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1198_ ( .D(N7113), .CP(clk), 
        .Q(inner_first_stage_data_reg[1198]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1197_ ( .D(N7112), .CP(clk), 
        .Q(inner_first_stage_data_reg[1197]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1196_ ( .D(N7111), .CP(clk), 
        .Q(inner_first_stage_data_reg[1196]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1195_ ( .D(N7110), .CP(clk), 
        .Q(inner_first_stage_data_reg[1195]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1194_ ( .D(N7109), .CP(clk), 
        .Q(inner_first_stage_data_reg[1194]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1193_ ( .D(N7108), .CP(clk), 
        .Q(inner_first_stage_data_reg[1193]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1192_ ( .D(N7107), .CP(clk), 
        .Q(inner_first_stage_data_reg[1192]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1191_ ( .D(N7106), .CP(clk), 
        .Q(inner_first_stage_data_reg[1191]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1190_ ( .D(N7105), .CP(clk), 
        .Q(inner_first_stage_data_reg[1190]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1189_ ( .D(N7104), .CP(clk), 
        .Q(inner_first_stage_data_reg[1189]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1188_ ( .D(N7103), .CP(clk), 
        .Q(inner_first_stage_data_reg[1188]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1187_ ( .D(N7102), .CP(clk), 
        .Q(inner_first_stage_data_reg[1187]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1186_ ( .D(N7101), .CP(clk), 
        .Q(inner_first_stage_data_reg[1186]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1185_ ( .D(N7100), .CP(clk), 
        .Q(inner_first_stage_data_reg[1185]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1184_ ( .D(N7099), .CP(clk), 
        .Q(inner_first_stage_data_reg[1184]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_38_ ( .D(N7314), .CP(clk), 
        .Q(inner_first_stage_valid_reg[38]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1247_ ( .D(N7346), .CP(clk), 
        .Q(inner_first_stage_data_reg[1247]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1246_ ( .D(N7345), .CP(clk), 
        .Q(inner_first_stage_data_reg[1246]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1245_ ( .D(N7344), .CP(clk), 
        .Q(inner_first_stage_data_reg[1245]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1244_ ( .D(N7343), .CP(clk), 
        .Q(inner_first_stage_data_reg[1244]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1243_ ( .D(N7342), .CP(clk), 
        .Q(inner_first_stage_data_reg[1243]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1242_ ( .D(N7341), .CP(clk), 
        .Q(inner_first_stage_data_reg[1242]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1241_ ( .D(N7340), .CP(clk), 
        .Q(inner_first_stage_data_reg[1241]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1240_ ( .D(N7339), .CP(clk), 
        .Q(inner_first_stage_data_reg[1240]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1239_ ( .D(N7338), .CP(clk), 
        .Q(inner_first_stage_data_reg[1239]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1238_ ( .D(N7337), .CP(clk), 
        .Q(inner_first_stage_data_reg[1238]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1237_ ( .D(N7336), .CP(clk), 
        .Q(inner_first_stage_data_reg[1237]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1236_ ( .D(N7335), .CP(clk), 
        .Q(inner_first_stage_data_reg[1236]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1235_ ( .D(N7334), .CP(clk), 
        .Q(inner_first_stage_data_reg[1235]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1234_ ( .D(N7333), .CP(clk), 
        .Q(inner_first_stage_data_reg[1234]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1233_ ( .D(N7332), .CP(clk), 
        .Q(inner_first_stage_data_reg[1233]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1232_ ( .D(N7331), .CP(clk), 
        .Q(inner_first_stage_data_reg[1232]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1231_ ( .D(N7330), .CP(clk), 
        .Q(inner_first_stage_data_reg[1231]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1230_ ( .D(N7329), .CP(clk), 
        .Q(inner_first_stage_data_reg[1230]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1229_ ( .D(N7328), .CP(clk), 
        .Q(inner_first_stage_data_reg[1229]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1228_ ( .D(N7327), .CP(clk), 
        .Q(inner_first_stage_data_reg[1228]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1227_ ( .D(N7326), .CP(clk), 
        .Q(inner_first_stage_data_reg[1227]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1226_ ( .D(N7325), .CP(clk), 
        .Q(inner_first_stage_data_reg[1226]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1225_ ( .D(N7324), .CP(clk), 
        .Q(inner_first_stage_data_reg[1225]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1224_ ( .D(N7323), .CP(clk), 
        .Q(inner_first_stage_data_reg[1224]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1223_ ( .D(N7322), .CP(clk), 
        .Q(inner_first_stage_data_reg[1223]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1222_ ( .D(N7321), .CP(clk), 
        .Q(inner_first_stage_data_reg[1222]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1221_ ( .D(N7320), .CP(clk), 
        .Q(inner_first_stage_data_reg[1221]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1220_ ( .D(N7319), .CP(clk), 
        .Q(inner_first_stage_data_reg[1220]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1219_ ( .D(N7318), .CP(clk), 
        .Q(inner_first_stage_data_reg[1219]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1218_ ( .D(N7317), .CP(clk), 
        .Q(inner_first_stage_data_reg[1218]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1217_ ( .D(N7316), .CP(clk), 
        .Q(inner_first_stage_data_reg[1217]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1216_ ( .D(N7315), .CP(clk), 
        .Q(inner_first_stage_data_reg[1216]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1279_ ( .D(N7562), .CP(clk), 
        .Q(inner_first_stage_data_reg[1279]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1278_ ( .D(N7561), .CP(clk), 
        .Q(inner_first_stage_data_reg[1278]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1277_ ( .D(N7560), .CP(clk), 
        .Q(inner_first_stage_data_reg[1277]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1276_ ( .D(N7559), .CP(clk), 
        .Q(inner_first_stage_data_reg[1276]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1275_ ( .D(N7558), .CP(clk), 
        .Q(inner_first_stage_data_reg[1275]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1274_ ( .D(N7557), .CP(clk), 
        .Q(inner_first_stage_data_reg[1274]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1273_ ( .D(N7556), .CP(clk), 
        .Q(inner_first_stage_data_reg[1273]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1272_ ( .D(N7555), .CP(clk), 
        .Q(inner_first_stage_data_reg[1272]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1271_ ( .D(N7554), .CP(clk), 
        .Q(inner_first_stage_data_reg[1271]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1270_ ( .D(N7553), .CP(clk), 
        .Q(inner_first_stage_data_reg[1270]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1269_ ( .D(N7552), .CP(clk), 
        .Q(inner_first_stage_data_reg[1269]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1268_ ( .D(N7551), .CP(clk), 
        .Q(inner_first_stage_data_reg[1268]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1267_ ( .D(N7550), .CP(clk), 
        .Q(inner_first_stage_data_reg[1267]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1266_ ( .D(N7549), .CP(clk), 
        .Q(inner_first_stage_data_reg[1266]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1265_ ( .D(N7548), .CP(clk), 
        .Q(inner_first_stage_data_reg[1265]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1264_ ( .D(N7547), .CP(clk), 
        .Q(inner_first_stage_data_reg[1264]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1263_ ( .D(N7546), .CP(clk), 
        .Q(inner_first_stage_data_reg[1263]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1262_ ( .D(N7545), .CP(clk), 
        .Q(inner_first_stage_data_reg[1262]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1261_ ( .D(N7544), .CP(clk), 
        .Q(inner_first_stage_data_reg[1261]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1260_ ( .D(N7543), .CP(clk), 
        .Q(inner_first_stage_data_reg[1260]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1259_ ( .D(N7542), .CP(clk), 
        .Q(inner_first_stage_data_reg[1259]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1258_ ( .D(N7541), .CP(clk), 
        .Q(inner_first_stage_data_reg[1258]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1257_ ( .D(N7540), .CP(clk), 
        .Q(inner_first_stage_data_reg[1257]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1256_ ( .D(N7539), .CP(clk), 
        .Q(inner_first_stage_data_reg[1256]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1255_ ( .D(N7538), .CP(clk), 
        .Q(inner_first_stage_data_reg[1255]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1254_ ( .D(N7537), .CP(clk), 
        .Q(inner_first_stage_data_reg[1254]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1253_ ( .D(N7536), .CP(clk), 
        .Q(inner_first_stage_data_reg[1253]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1252_ ( .D(N7535), .CP(clk), 
        .Q(inner_first_stage_data_reg[1252]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1251_ ( .D(N7534), .CP(clk), 
        .Q(inner_first_stage_data_reg[1251]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1250_ ( .D(N7533), .CP(clk), 
        .Q(inner_first_stage_data_reg[1250]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1249_ ( .D(N7532), .CP(clk), 
        .Q(inner_first_stage_data_reg[1249]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1248_ ( .D(N7531), .CP(clk), 
        .Q(inner_first_stage_data_reg[1248]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_40_ ( .D(N7764), .CP(clk), 
        .Q(inner_first_stage_valid_reg[40]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1311_ ( .D(N7796), .CP(clk), 
        .Q(inner_first_stage_data_reg[1311]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1310_ ( .D(N7795), .CP(clk), 
        .Q(inner_first_stage_data_reg[1310]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1309_ ( .D(N7794), .CP(clk), 
        .Q(inner_first_stage_data_reg[1309]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1308_ ( .D(N7793), .CP(clk), 
        .Q(inner_first_stage_data_reg[1308]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1307_ ( .D(N7792), .CP(clk), 
        .Q(inner_first_stage_data_reg[1307]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1306_ ( .D(N7791), .CP(clk), 
        .Q(inner_first_stage_data_reg[1306]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1305_ ( .D(N7790), .CP(clk), 
        .Q(inner_first_stage_data_reg[1305]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1304_ ( .D(N7789), .CP(clk), 
        .Q(inner_first_stage_data_reg[1304]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1303_ ( .D(N7788), .CP(clk), 
        .Q(inner_first_stage_data_reg[1303]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1302_ ( .D(N7787), .CP(clk), 
        .Q(inner_first_stage_data_reg[1302]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1301_ ( .D(N7786), .CP(clk), 
        .Q(inner_first_stage_data_reg[1301]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1300_ ( .D(N7785), .CP(clk), 
        .Q(inner_first_stage_data_reg[1300]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1299_ ( .D(N7784), .CP(clk), 
        .Q(inner_first_stage_data_reg[1299]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1298_ ( .D(N7783), .CP(clk), 
        .Q(inner_first_stage_data_reg[1298]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1297_ ( .D(N7782), .CP(clk), 
        .Q(inner_first_stage_data_reg[1297]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1296_ ( .D(N7781), .CP(clk), 
        .Q(inner_first_stage_data_reg[1296]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1295_ ( .D(N7780), .CP(clk), 
        .Q(inner_first_stage_data_reg[1295]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1294_ ( .D(N7779), .CP(clk), 
        .Q(inner_first_stage_data_reg[1294]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1293_ ( .D(N7778), .CP(clk), 
        .Q(inner_first_stage_data_reg[1293]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1292_ ( .D(N7777), .CP(clk), 
        .Q(inner_first_stage_data_reg[1292]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1291_ ( .D(N7776), .CP(clk), 
        .Q(inner_first_stage_data_reg[1291]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1290_ ( .D(N7775), .CP(clk), 
        .Q(inner_first_stage_data_reg[1290]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1289_ ( .D(N7774), .CP(clk), 
        .Q(inner_first_stage_data_reg[1289]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1288_ ( .D(N7773), .CP(clk), 
        .Q(inner_first_stage_data_reg[1288]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1287_ ( .D(N7772), .CP(clk), 
        .Q(inner_first_stage_data_reg[1287]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1286_ ( .D(N7771), .CP(clk), 
        .Q(inner_first_stage_data_reg[1286]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1285_ ( .D(N7770), .CP(clk), 
        .Q(inner_first_stage_data_reg[1285]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1284_ ( .D(N7769), .CP(clk), 
        .Q(inner_first_stage_data_reg[1284]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1283_ ( .D(N7768), .CP(clk), 
        .Q(inner_first_stage_data_reg[1283]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1282_ ( .D(N7767), .CP(clk), 
        .Q(inner_first_stage_data_reg[1282]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1281_ ( .D(N7766), .CP(clk), 
        .Q(inner_first_stage_data_reg[1281]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1280_ ( .D(N7765), .CP(clk), 
        .Q(inner_first_stage_data_reg[1280]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_41_ ( .D(N7852), .CP(clk), 
        .Q(inner_first_stage_valid_reg[41]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1343_ ( .D(N7884), .CP(clk), 
        .Q(inner_first_stage_data_reg[1343]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1342_ ( .D(N7883), .CP(clk), 
        .Q(inner_first_stage_data_reg[1342]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1341_ ( .D(N7882), .CP(clk), 
        .Q(inner_first_stage_data_reg[1341]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1340_ ( .D(N7881), .CP(clk), 
        .Q(inner_first_stage_data_reg[1340]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1339_ ( .D(N7880), .CP(clk), 
        .Q(inner_first_stage_data_reg[1339]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1338_ ( .D(N7879), .CP(clk), 
        .Q(inner_first_stage_data_reg[1338]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1337_ ( .D(N7878), .CP(clk), 
        .Q(inner_first_stage_data_reg[1337]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1336_ ( .D(N7877), .CP(clk), 
        .Q(inner_first_stage_data_reg[1336]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1335_ ( .D(N7876), .CP(clk), 
        .Q(inner_first_stage_data_reg[1335]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1334_ ( .D(N7875), .CP(clk), 
        .Q(inner_first_stage_data_reg[1334]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1333_ ( .D(N7874), .CP(clk), 
        .Q(inner_first_stage_data_reg[1333]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1332_ ( .D(N7873), .CP(clk), 
        .Q(inner_first_stage_data_reg[1332]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1331_ ( .D(N7872), .CP(clk), 
        .Q(inner_first_stage_data_reg[1331]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1330_ ( .D(N7871), .CP(clk), 
        .Q(inner_first_stage_data_reg[1330]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1329_ ( .D(N7870), .CP(clk), 
        .Q(inner_first_stage_data_reg[1329]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1328_ ( .D(N7869), .CP(clk), 
        .Q(inner_first_stage_data_reg[1328]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1327_ ( .D(N7868), .CP(clk), 
        .Q(inner_first_stage_data_reg[1327]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1326_ ( .D(N7867), .CP(clk), 
        .Q(inner_first_stage_data_reg[1326]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1325_ ( .D(N7866), .CP(clk), 
        .Q(inner_first_stage_data_reg[1325]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1324_ ( .D(N7865), .CP(clk), 
        .Q(inner_first_stage_data_reg[1324]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1323_ ( .D(N7864), .CP(clk), 
        .Q(inner_first_stage_data_reg[1323]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1322_ ( .D(N7863), .CP(clk), 
        .Q(inner_first_stage_data_reg[1322]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1321_ ( .D(N7862), .CP(clk), 
        .Q(inner_first_stage_data_reg[1321]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1320_ ( .D(N7861), .CP(clk), 
        .Q(inner_first_stage_data_reg[1320]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1319_ ( .D(N7860), .CP(clk), 
        .Q(inner_first_stage_data_reg[1319]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1318_ ( .D(N7859), .CP(clk), 
        .Q(inner_first_stage_data_reg[1318]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1317_ ( .D(N7858), .CP(clk), 
        .Q(inner_first_stage_data_reg[1317]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1316_ ( .D(N7857), .CP(clk), 
        .Q(inner_first_stage_data_reg[1316]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1315_ ( .D(N7856), .CP(clk), 
        .Q(inner_first_stage_data_reg[1315]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1314_ ( .D(N7855), .CP(clk), 
        .Q(inner_first_stage_data_reg[1314]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1313_ ( .D(N7854), .CP(clk), 
        .Q(inner_first_stage_data_reg[1313]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1312_ ( .D(N7853), .CP(clk), 
        .Q(inner_first_stage_data_reg[1312]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_42_ ( .D(N7940), .CP(clk), 
        .Q(inner_first_stage_valid_reg[42]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1375_ ( .D(N7972), .CP(clk), 
        .Q(inner_first_stage_data_reg[1375]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1374_ ( .D(N7971), .CP(clk), 
        .Q(inner_first_stage_data_reg[1374]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1373_ ( .D(N7970), .CP(clk), 
        .Q(inner_first_stage_data_reg[1373]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1372_ ( .D(N7969), .CP(clk), 
        .Q(inner_first_stage_data_reg[1372]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1371_ ( .D(N7968), .CP(clk), 
        .Q(inner_first_stage_data_reg[1371]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1370_ ( .D(N7967), .CP(clk), 
        .Q(inner_first_stage_data_reg[1370]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1369_ ( .D(N7966), .CP(clk), 
        .Q(inner_first_stage_data_reg[1369]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1368_ ( .D(N7965), .CP(clk), 
        .Q(inner_first_stage_data_reg[1368]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1367_ ( .D(N7964), .CP(clk), 
        .Q(inner_first_stage_data_reg[1367]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1366_ ( .D(N7963), .CP(clk), 
        .Q(inner_first_stage_data_reg[1366]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1365_ ( .D(N7962), .CP(clk), 
        .Q(inner_first_stage_data_reg[1365]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1364_ ( .D(N7961), .CP(clk), 
        .Q(inner_first_stage_data_reg[1364]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1363_ ( .D(N7960), .CP(clk), 
        .Q(inner_first_stage_data_reg[1363]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1362_ ( .D(N7959), .CP(clk), 
        .Q(inner_first_stage_data_reg[1362]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1361_ ( .D(N7958), .CP(clk), 
        .Q(inner_first_stage_data_reg[1361]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1360_ ( .D(N7957), .CP(clk), 
        .Q(inner_first_stage_data_reg[1360]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1359_ ( .D(N7956), .CP(clk), 
        .Q(inner_first_stage_data_reg[1359]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1358_ ( .D(N7955), .CP(clk), 
        .Q(inner_first_stage_data_reg[1358]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1357_ ( .D(N7954), .CP(clk), 
        .Q(inner_first_stage_data_reg[1357]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1356_ ( .D(N7953), .CP(clk), 
        .Q(inner_first_stage_data_reg[1356]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1355_ ( .D(N7952), .CP(clk), 
        .Q(inner_first_stage_data_reg[1355]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1354_ ( .D(N7951), .CP(clk), 
        .Q(inner_first_stage_data_reg[1354]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1353_ ( .D(N7950), .CP(clk), 
        .Q(inner_first_stage_data_reg[1353]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1352_ ( .D(N7949), .CP(clk), 
        .Q(inner_first_stage_data_reg[1352]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1351_ ( .D(N7948), .CP(clk), 
        .Q(inner_first_stage_data_reg[1351]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1350_ ( .D(N7947), .CP(clk), 
        .Q(inner_first_stage_data_reg[1350]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1349_ ( .D(N7946), .CP(clk), 
        .Q(inner_first_stage_data_reg[1349]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1348_ ( .D(N7945), .CP(clk), 
        .Q(inner_first_stage_data_reg[1348]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1347_ ( .D(N7944), .CP(clk), 
        .Q(inner_first_stage_data_reg[1347]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1346_ ( .D(N7943), .CP(clk), 
        .Q(inner_first_stage_data_reg[1346]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1345_ ( .D(N7942), .CP(clk), 
        .Q(inner_first_stage_data_reg[1345]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1344_ ( .D(N7941), .CP(clk), 
        .Q(inner_first_stage_data_reg[1344]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_43_ ( .D(N8028), .CP(clk), 
        .Q(inner_first_stage_valid_reg[43]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1407_ ( .D(N8060), .CP(clk), 
        .Q(inner_first_stage_data_reg[1407]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1406_ ( .D(N8059), .CP(clk), 
        .Q(inner_first_stage_data_reg[1406]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1405_ ( .D(N8058), .CP(clk), 
        .Q(inner_first_stage_data_reg[1405]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1404_ ( .D(N8057), .CP(clk), 
        .Q(inner_first_stage_data_reg[1404]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1403_ ( .D(N8056), .CP(clk), 
        .Q(inner_first_stage_data_reg[1403]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1402_ ( .D(N8055), .CP(clk), 
        .Q(inner_first_stage_data_reg[1402]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1401_ ( .D(N8054), .CP(clk), 
        .Q(inner_first_stage_data_reg[1401]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1400_ ( .D(N8053), .CP(clk), 
        .Q(inner_first_stage_data_reg[1400]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1399_ ( .D(N8052), .CP(clk), 
        .Q(inner_first_stage_data_reg[1399]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1398_ ( .D(N8051), .CP(clk), 
        .Q(inner_first_stage_data_reg[1398]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1397_ ( .D(N8050), .CP(clk), 
        .Q(inner_first_stage_data_reg[1397]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1396_ ( .D(N8049), .CP(clk), 
        .Q(inner_first_stage_data_reg[1396]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1395_ ( .D(N8048), .CP(clk), 
        .Q(inner_first_stage_data_reg[1395]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1394_ ( .D(N8047), .CP(clk), 
        .Q(inner_first_stage_data_reg[1394]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1393_ ( .D(N8046), .CP(clk), 
        .Q(inner_first_stage_data_reg[1393]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1392_ ( .D(N8045), .CP(clk), 
        .Q(inner_first_stage_data_reg[1392]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1391_ ( .D(N8044), .CP(clk), 
        .Q(inner_first_stage_data_reg[1391]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1390_ ( .D(N8043), .CP(clk), 
        .Q(inner_first_stage_data_reg[1390]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1389_ ( .D(N8042), .CP(clk), 
        .Q(inner_first_stage_data_reg[1389]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1388_ ( .D(N8041), .CP(clk), 
        .Q(inner_first_stage_data_reg[1388]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1387_ ( .D(N8040), .CP(clk), 
        .Q(inner_first_stage_data_reg[1387]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1386_ ( .D(N8039), .CP(clk), 
        .Q(inner_first_stage_data_reg[1386]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1385_ ( .D(N8038), .CP(clk), 
        .Q(inner_first_stage_data_reg[1385]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1384_ ( .D(N8037), .CP(clk), 
        .Q(inner_first_stage_data_reg[1384]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1383_ ( .D(N8036), .CP(clk), 
        .Q(inner_first_stage_data_reg[1383]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1382_ ( .D(N8035), .CP(clk), 
        .Q(inner_first_stage_data_reg[1382]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1381_ ( .D(N8034), .CP(clk), 
        .Q(inner_first_stage_data_reg[1381]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1380_ ( .D(N8033), .CP(clk), 
        .Q(inner_first_stage_data_reg[1380]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1379_ ( .D(N8032), .CP(clk), 
        .Q(inner_first_stage_data_reg[1379]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1378_ ( .D(N8031), .CP(clk), 
        .Q(inner_first_stage_data_reg[1378]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1377_ ( .D(N8030), .CP(clk), 
        .Q(inner_first_stage_data_reg[1377]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1376_ ( .D(N8029), .CP(clk), 
        .Q(inner_first_stage_data_reg[1376]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_44_ ( .D(N8116), .CP(clk), 
        .Q(inner_first_stage_valid_reg[44]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1439_ ( .D(N8148), .CP(clk), 
        .Q(inner_first_stage_data_reg[1439]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1438_ ( .D(N8147), .CP(clk), 
        .Q(inner_first_stage_data_reg[1438]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1437_ ( .D(N8146), .CP(clk), 
        .Q(inner_first_stage_data_reg[1437]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1436_ ( .D(N8145), .CP(clk), 
        .Q(inner_first_stage_data_reg[1436]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1435_ ( .D(N8144), .CP(clk), 
        .Q(inner_first_stage_data_reg[1435]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1434_ ( .D(N8143), .CP(clk), 
        .Q(inner_first_stage_data_reg[1434]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1433_ ( .D(N8142), .CP(clk), 
        .Q(inner_first_stage_data_reg[1433]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1432_ ( .D(N8141), .CP(clk), 
        .Q(inner_first_stage_data_reg[1432]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1431_ ( .D(N8140), .CP(clk), 
        .Q(inner_first_stage_data_reg[1431]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1430_ ( .D(N8139), .CP(clk), 
        .Q(inner_first_stage_data_reg[1430]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1429_ ( .D(N8138), .CP(clk), 
        .Q(inner_first_stage_data_reg[1429]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1428_ ( .D(N8137), .CP(clk), 
        .Q(inner_first_stage_data_reg[1428]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1427_ ( .D(N8136), .CP(clk), 
        .Q(inner_first_stage_data_reg[1427]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1426_ ( .D(N8135), .CP(clk), 
        .Q(inner_first_stage_data_reg[1426]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1425_ ( .D(N8134), .CP(clk), 
        .Q(inner_first_stage_data_reg[1425]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1424_ ( .D(N8133), .CP(clk), 
        .Q(inner_first_stage_data_reg[1424]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1423_ ( .D(N8132), .CP(clk), 
        .Q(inner_first_stage_data_reg[1423]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1422_ ( .D(N8131), .CP(clk), 
        .Q(inner_first_stage_data_reg[1422]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1421_ ( .D(N8130), .CP(clk), 
        .Q(inner_first_stage_data_reg[1421]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1420_ ( .D(N8129), .CP(clk), 
        .Q(inner_first_stage_data_reg[1420]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1419_ ( .D(N8128), .CP(clk), 
        .Q(inner_first_stage_data_reg[1419]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1418_ ( .D(N8127), .CP(clk), 
        .Q(inner_first_stage_data_reg[1418]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1417_ ( .D(N8126), .CP(clk), 
        .Q(inner_first_stage_data_reg[1417]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1416_ ( .D(N8125), .CP(clk), 
        .Q(inner_first_stage_data_reg[1416]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1415_ ( .D(N8124), .CP(clk), 
        .Q(inner_first_stage_data_reg[1415]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1414_ ( .D(N8123), .CP(clk), 
        .Q(inner_first_stage_data_reg[1414]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1413_ ( .D(N8122), .CP(clk), 
        .Q(inner_first_stage_data_reg[1413]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1412_ ( .D(N8121), .CP(clk), 
        .Q(inner_first_stage_data_reg[1412]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1411_ ( .D(N8120), .CP(clk), 
        .Q(inner_first_stage_data_reg[1411]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1410_ ( .D(N8119), .CP(clk), 
        .Q(inner_first_stage_data_reg[1410]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1409_ ( .D(N8118), .CP(clk), 
        .Q(inner_first_stage_data_reg[1409]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1408_ ( .D(N8117), .CP(clk), 
        .Q(inner_first_stage_data_reg[1408]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_45_ ( .D(N8204), .CP(clk), 
        .Q(inner_first_stage_valid_reg[45]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1471_ ( .D(N8236), .CP(clk), 
        .Q(inner_first_stage_data_reg[1471]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1470_ ( .D(N8235), .CP(clk), 
        .Q(inner_first_stage_data_reg[1470]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1469_ ( .D(N8234), .CP(clk), 
        .Q(inner_first_stage_data_reg[1469]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1468_ ( .D(N8233), .CP(clk), 
        .Q(inner_first_stage_data_reg[1468]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1467_ ( .D(N8232), .CP(clk), 
        .Q(inner_first_stage_data_reg[1467]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1466_ ( .D(N8231), .CP(clk), 
        .Q(inner_first_stage_data_reg[1466]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1465_ ( .D(N8230), .CP(clk), 
        .Q(inner_first_stage_data_reg[1465]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1464_ ( .D(N8229), .CP(clk), 
        .Q(inner_first_stage_data_reg[1464]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1463_ ( .D(N8228), .CP(clk), 
        .Q(inner_first_stage_data_reg[1463]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1462_ ( .D(N8227), .CP(clk), 
        .Q(inner_first_stage_data_reg[1462]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1461_ ( .D(N8226), .CP(clk), 
        .Q(inner_first_stage_data_reg[1461]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1460_ ( .D(N8225), .CP(clk), 
        .Q(inner_first_stage_data_reg[1460]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1459_ ( .D(N8224), .CP(clk), 
        .Q(inner_first_stage_data_reg[1459]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1458_ ( .D(N8223), .CP(clk), 
        .Q(inner_first_stage_data_reg[1458]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1457_ ( .D(N8222), .CP(clk), 
        .Q(inner_first_stage_data_reg[1457]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1456_ ( .D(N8221), .CP(clk), 
        .Q(inner_first_stage_data_reg[1456]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1455_ ( .D(N8220), .CP(clk), 
        .Q(inner_first_stage_data_reg[1455]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1454_ ( .D(N8219), .CP(clk), 
        .Q(inner_first_stage_data_reg[1454]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1453_ ( .D(N8218), .CP(clk), 
        .Q(inner_first_stage_data_reg[1453]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1452_ ( .D(N8217), .CP(clk), 
        .Q(inner_first_stage_data_reg[1452]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1451_ ( .D(N8216), .CP(clk), 
        .Q(inner_first_stage_data_reg[1451]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1450_ ( .D(N8215), .CP(clk), 
        .Q(inner_first_stage_data_reg[1450]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1449_ ( .D(N8214), .CP(clk), 
        .Q(inner_first_stage_data_reg[1449]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1448_ ( .D(N8213), .CP(clk), 
        .Q(inner_first_stage_data_reg[1448]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1447_ ( .D(N8212), .CP(clk), 
        .Q(inner_first_stage_data_reg[1447]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1446_ ( .D(N8211), .CP(clk), 
        .Q(inner_first_stage_data_reg[1446]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1445_ ( .D(N8210), .CP(clk), 
        .Q(inner_first_stage_data_reg[1445]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1444_ ( .D(N8209), .CP(clk), 
        .Q(inner_first_stage_data_reg[1444]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1443_ ( .D(N8208), .CP(clk), 
        .Q(inner_first_stage_data_reg[1443]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1442_ ( .D(N8207), .CP(clk), 
        .Q(inner_first_stage_data_reg[1442]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1441_ ( .D(N8206), .CP(clk), 
        .Q(inner_first_stage_data_reg[1441]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1440_ ( .D(N8205), .CP(clk), 
        .Q(inner_first_stage_data_reg[1440]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_46_ ( .D(N8292), .CP(clk), 
        .Q(inner_first_stage_valid_reg[46]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1503_ ( .D(N8324), .CP(clk), 
        .Q(inner_first_stage_data_reg[1503]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1502_ ( .D(N8323), .CP(clk), 
        .Q(inner_first_stage_data_reg[1502]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1501_ ( .D(N8322), .CP(clk), 
        .Q(inner_first_stage_data_reg[1501]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1500_ ( .D(N8321), .CP(clk), 
        .Q(inner_first_stage_data_reg[1500]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1499_ ( .D(N8320), .CP(clk), 
        .Q(inner_first_stage_data_reg[1499]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1498_ ( .D(N8319), .CP(clk), 
        .Q(inner_first_stage_data_reg[1498]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1497_ ( .D(N8318), .CP(clk), 
        .Q(inner_first_stage_data_reg[1497]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1496_ ( .D(N8317), .CP(clk), 
        .Q(inner_first_stage_data_reg[1496]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1495_ ( .D(N8316), .CP(clk), 
        .Q(inner_first_stage_data_reg[1495]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1494_ ( .D(N8315), .CP(clk), 
        .Q(inner_first_stage_data_reg[1494]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1493_ ( .D(N8314), .CP(clk), 
        .Q(inner_first_stage_data_reg[1493]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1492_ ( .D(N8313), .CP(clk), 
        .Q(inner_first_stage_data_reg[1492]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1491_ ( .D(N8312), .CP(clk), 
        .Q(inner_first_stage_data_reg[1491]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1490_ ( .D(N8311), .CP(clk), 
        .Q(inner_first_stage_data_reg[1490]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1489_ ( .D(N8310), .CP(clk), 
        .Q(inner_first_stage_data_reg[1489]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1488_ ( .D(N8309), .CP(clk), 
        .Q(inner_first_stage_data_reg[1488]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1487_ ( .D(N8308), .CP(clk), 
        .Q(inner_first_stage_data_reg[1487]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1486_ ( .D(N8307), .CP(clk), 
        .Q(inner_first_stage_data_reg[1486]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1485_ ( .D(N8306), .CP(clk), 
        .Q(inner_first_stage_data_reg[1485]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1484_ ( .D(N8305), .CP(clk), 
        .Q(inner_first_stage_data_reg[1484]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1483_ ( .D(N8304), .CP(clk), 
        .Q(inner_first_stage_data_reg[1483]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1482_ ( .D(N8303), .CP(clk), 
        .Q(inner_first_stage_data_reg[1482]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1481_ ( .D(N8302), .CP(clk), 
        .Q(inner_first_stage_data_reg[1481]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1480_ ( .D(N8301), .CP(clk), 
        .Q(inner_first_stage_data_reg[1480]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1479_ ( .D(N8300), .CP(clk), 
        .Q(inner_first_stage_data_reg[1479]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1478_ ( .D(N8299), .CP(clk), 
        .Q(inner_first_stage_data_reg[1478]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1477_ ( .D(N8298), .CP(clk), 
        .Q(inner_first_stage_data_reg[1477]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1476_ ( .D(N8297), .CP(clk), 
        .Q(inner_first_stage_data_reg[1476]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1475_ ( .D(N8296), .CP(clk), 
        .Q(inner_first_stage_data_reg[1475]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1474_ ( .D(N8295), .CP(clk), 
        .Q(inner_first_stage_data_reg[1474]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1473_ ( .D(N8294), .CP(clk), 
        .Q(inner_first_stage_data_reg[1473]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1472_ ( .D(N8293), .CP(clk), 
        .Q(inner_first_stage_data_reg[1472]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_47_ ( .D(N8380), .CP(clk), 
        .Q(inner_first_stage_valid_reg[47]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1535_ ( .D(N8412), .CP(clk), 
        .Q(inner_first_stage_data_reg[1535]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1534_ ( .D(N8411), .CP(clk), 
        .Q(inner_first_stage_data_reg[1534]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1533_ ( .D(N8410), .CP(clk), 
        .Q(inner_first_stage_data_reg[1533]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1532_ ( .D(N8409), .CP(clk), 
        .Q(inner_first_stage_data_reg[1532]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1531_ ( .D(N8408), .CP(clk), 
        .Q(inner_first_stage_data_reg[1531]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1530_ ( .D(N8407), .CP(clk), 
        .Q(inner_first_stage_data_reg[1530]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1529_ ( .D(N8406), .CP(clk), 
        .Q(inner_first_stage_data_reg[1529]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1528_ ( .D(N8405), .CP(clk), 
        .Q(inner_first_stage_data_reg[1528]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1527_ ( .D(N8404), .CP(clk), 
        .Q(inner_first_stage_data_reg[1527]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1526_ ( .D(N8403), .CP(clk), 
        .Q(inner_first_stage_data_reg[1526]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1525_ ( .D(N8402), .CP(clk), 
        .Q(inner_first_stage_data_reg[1525]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1524_ ( .D(N8401), .CP(clk), 
        .Q(inner_first_stage_data_reg[1524]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1523_ ( .D(N8400), .CP(clk), 
        .Q(inner_first_stage_data_reg[1523]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1522_ ( .D(N8399), .CP(clk), 
        .Q(inner_first_stage_data_reg[1522]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1521_ ( .D(N8398), .CP(clk), 
        .Q(inner_first_stage_data_reg[1521]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1520_ ( .D(N8397), .CP(clk), 
        .Q(inner_first_stage_data_reg[1520]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1519_ ( .D(N8396), .CP(clk), 
        .Q(inner_first_stage_data_reg[1519]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1518_ ( .D(N8395), .CP(clk), 
        .Q(inner_first_stage_data_reg[1518]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1517_ ( .D(N8394), .CP(clk), 
        .Q(inner_first_stage_data_reg[1517]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1516_ ( .D(N8393), .CP(clk), 
        .Q(inner_first_stage_data_reg[1516]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1515_ ( .D(N8392), .CP(clk), 
        .Q(inner_first_stage_data_reg[1515]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1514_ ( .D(N8391), .CP(clk), 
        .Q(inner_first_stage_data_reg[1514]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1513_ ( .D(N8390), .CP(clk), 
        .Q(inner_first_stage_data_reg[1513]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1512_ ( .D(N8389), .CP(clk), 
        .Q(inner_first_stage_data_reg[1512]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1511_ ( .D(N8388), .CP(clk), 
        .Q(inner_first_stage_data_reg[1511]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1510_ ( .D(N8387), .CP(clk), 
        .Q(inner_first_stage_data_reg[1510]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1509_ ( .D(N8386), .CP(clk), 
        .Q(inner_first_stage_data_reg[1509]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1508_ ( .D(N8385), .CP(clk), 
        .Q(inner_first_stage_data_reg[1508]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1507_ ( .D(N8384), .CP(clk), 
        .Q(inner_first_stage_data_reg[1507]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1506_ ( .D(N8383), .CP(clk), 
        .Q(inner_first_stage_data_reg[1506]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1505_ ( .D(N8382), .CP(clk), 
        .Q(inner_first_stage_data_reg[1505]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1504_ ( .D(N8381), .CP(clk), 
        .Q(inner_first_stage_data_reg[1504]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_48_ ( .D(N8742), .CP(clk), 
        .Q(inner_first_stage_valid_reg[48]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1567_ ( .D(N8774), .CP(clk), 
        .Q(inner_first_stage_data_reg[1567]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1566_ ( .D(N8773), .CP(clk), 
        .Q(inner_first_stage_data_reg[1566]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1565_ ( .D(N8772), .CP(clk), 
        .Q(inner_first_stage_data_reg[1565]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1564_ ( .D(N8771), .CP(clk), 
        .Q(inner_first_stage_data_reg[1564]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1563_ ( .D(N8770), .CP(clk), 
        .Q(inner_first_stage_data_reg[1563]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1562_ ( .D(N8769), .CP(clk), 
        .Q(inner_first_stage_data_reg[1562]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1561_ ( .D(N8768), .CP(clk), 
        .Q(inner_first_stage_data_reg[1561]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1560_ ( .D(N8767), .CP(clk), 
        .Q(inner_first_stage_data_reg[1560]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1559_ ( .D(N8766), .CP(clk), 
        .Q(inner_first_stage_data_reg[1559]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1558_ ( .D(N8765), .CP(clk), 
        .Q(inner_first_stage_data_reg[1558]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1557_ ( .D(N8764), .CP(clk), 
        .Q(inner_first_stage_data_reg[1557]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1556_ ( .D(N8763), .CP(clk), 
        .Q(inner_first_stage_data_reg[1556]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1555_ ( .D(N8762), .CP(clk), 
        .Q(inner_first_stage_data_reg[1555]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1554_ ( .D(N8761), .CP(clk), 
        .Q(inner_first_stage_data_reg[1554]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1553_ ( .D(N8760), .CP(clk), 
        .Q(inner_first_stage_data_reg[1553]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1552_ ( .D(N8759), .CP(clk), 
        .Q(inner_first_stage_data_reg[1552]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1551_ ( .D(N8758), .CP(clk), 
        .Q(inner_first_stage_data_reg[1551]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1550_ ( .D(N8757), .CP(clk), 
        .Q(inner_first_stage_data_reg[1550]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1549_ ( .D(N8756), .CP(clk), 
        .Q(inner_first_stage_data_reg[1549]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1548_ ( .D(N8755), .CP(clk), 
        .Q(inner_first_stage_data_reg[1548]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1547_ ( .D(N8754), .CP(clk), 
        .Q(inner_first_stage_data_reg[1547]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1546_ ( .D(N8753), .CP(clk), 
        .Q(inner_first_stage_data_reg[1546]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1545_ ( .D(N8752), .CP(clk), 
        .Q(inner_first_stage_data_reg[1545]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1544_ ( .D(N8751), .CP(clk), 
        .Q(inner_first_stage_data_reg[1544]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1543_ ( .D(N8750), .CP(clk), 
        .Q(inner_first_stage_data_reg[1543]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1542_ ( .D(N8749), .CP(clk), 
        .Q(inner_first_stage_data_reg[1542]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1541_ ( .D(N8748), .CP(clk), 
        .Q(inner_first_stage_data_reg[1541]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1540_ ( .D(N8747), .CP(clk), 
        .Q(inner_first_stage_data_reg[1540]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1539_ ( .D(N8746), .CP(clk), 
        .Q(inner_first_stage_data_reg[1539]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1538_ ( .D(N8745), .CP(clk), 
        .Q(inner_first_stage_data_reg[1538]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1537_ ( .D(N8744), .CP(clk), 
        .Q(inner_first_stage_data_reg[1537]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1536_ ( .D(N8743), .CP(clk), 
        .Q(inner_first_stage_data_reg[1536]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_49_ ( .D(N8958), .CP(clk), 
        .Q(inner_first_stage_valid_reg[49]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1599_ ( .D(N8990), .CP(clk), 
        .Q(inner_first_stage_data_reg[1599]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1598_ ( .D(N8989), .CP(clk), 
        .Q(inner_first_stage_data_reg[1598]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1597_ ( .D(N8988), .CP(clk), 
        .Q(inner_first_stage_data_reg[1597]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1596_ ( .D(N8987), .CP(clk), 
        .Q(inner_first_stage_data_reg[1596]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1595_ ( .D(N8986), .CP(clk), 
        .Q(inner_first_stage_data_reg[1595]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1594_ ( .D(N8985), .CP(clk), 
        .Q(inner_first_stage_data_reg[1594]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1593_ ( .D(N8984), .CP(clk), 
        .Q(inner_first_stage_data_reg[1593]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1592_ ( .D(N8983), .CP(clk), 
        .Q(inner_first_stage_data_reg[1592]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1591_ ( .D(N8982), .CP(clk), 
        .Q(inner_first_stage_data_reg[1591]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1590_ ( .D(N8981), .CP(clk), 
        .Q(inner_first_stage_data_reg[1590]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1589_ ( .D(N8980), .CP(clk), 
        .Q(inner_first_stage_data_reg[1589]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1588_ ( .D(N8979), .CP(clk), 
        .Q(inner_first_stage_data_reg[1588]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1587_ ( .D(N8978), .CP(clk), 
        .Q(inner_first_stage_data_reg[1587]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1586_ ( .D(N8977), .CP(clk), 
        .Q(inner_first_stage_data_reg[1586]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1585_ ( .D(N8976), .CP(clk), 
        .Q(inner_first_stage_data_reg[1585]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1584_ ( .D(N8975), .CP(clk), 
        .Q(inner_first_stage_data_reg[1584]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1583_ ( .D(N8974), .CP(clk), 
        .Q(inner_first_stage_data_reg[1583]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1582_ ( .D(N8973), .CP(clk), 
        .Q(inner_first_stage_data_reg[1582]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1581_ ( .D(N8972), .CP(clk), 
        .Q(inner_first_stage_data_reg[1581]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1580_ ( .D(N8971), .CP(clk), 
        .Q(inner_first_stage_data_reg[1580]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1579_ ( .D(N8970), .CP(clk), 
        .Q(inner_first_stage_data_reg[1579]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1578_ ( .D(N8969), .CP(clk), 
        .Q(inner_first_stage_data_reg[1578]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1577_ ( .D(N8968), .CP(clk), 
        .Q(inner_first_stage_data_reg[1577]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1576_ ( .D(N8967), .CP(clk), 
        .Q(inner_first_stage_data_reg[1576]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1575_ ( .D(N8966), .CP(clk), 
        .Q(inner_first_stage_data_reg[1575]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1574_ ( .D(N8965), .CP(clk), 
        .Q(inner_first_stage_data_reg[1574]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1573_ ( .D(N8964), .CP(clk), 
        .Q(inner_first_stage_data_reg[1573]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1572_ ( .D(N8963), .CP(clk), 
        .Q(inner_first_stage_data_reg[1572]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1571_ ( .D(N8962), .CP(clk), 
        .Q(inner_first_stage_data_reg[1571]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1570_ ( .D(N8961), .CP(clk), 
        .Q(inner_first_stage_data_reg[1570]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1569_ ( .D(N8960), .CP(clk), 
        .Q(inner_first_stage_data_reg[1569]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1568_ ( .D(N8959), .CP(clk), 
        .Q(inner_first_stage_data_reg[1568]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_50_ ( .D(N9174), .CP(clk), 
        .Q(inner_first_stage_valid_reg[50]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1631_ ( .D(N9206), .CP(clk), 
        .Q(inner_first_stage_data_reg[1631]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1630_ ( .D(N9205), .CP(clk), 
        .Q(inner_first_stage_data_reg[1630]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1629_ ( .D(N9204), .CP(clk), 
        .Q(inner_first_stage_data_reg[1629]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1628_ ( .D(N9203), .CP(clk), 
        .Q(inner_first_stage_data_reg[1628]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1627_ ( .D(N9202), .CP(clk), 
        .Q(inner_first_stage_data_reg[1627]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1626_ ( .D(N9201), .CP(clk), 
        .Q(inner_first_stage_data_reg[1626]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1625_ ( .D(N9200), .CP(clk), 
        .Q(inner_first_stage_data_reg[1625]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1624_ ( .D(N9199), .CP(clk), 
        .Q(inner_first_stage_data_reg[1624]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1623_ ( .D(N9198), .CP(clk), 
        .Q(inner_first_stage_data_reg[1623]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1622_ ( .D(N9197), .CP(clk), 
        .Q(inner_first_stage_data_reg[1622]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1621_ ( .D(N9196), .CP(clk), 
        .Q(inner_first_stage_data_reg[1621]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1620_ ( .D(N9195), .CP(clk), 
        .Q(inner_first_stage_data_reg[1620]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1619_ ( .D(N9194), .CP(clk), 
        .Q(inner_first_stage_data_reg[1619]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1618_ ( .D(N9193), .CP(clk), 
        .Q(inner_first_stage_data_reg[1618]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1617_ ( .D(N9192), .CP(clk), 
        .Q(inner_first_stage_data_reg[1617]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1616_ ( .D(N9191), .CP(clk), 
        .Q(inner_first_stage_data_reg[1616]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1615_ ( .D(N9190), .CP(clk), 
        .Q(inner_first_stage_data_reg[1615]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1614_ ( .D(N9189), .CP(clk), 
        .Q(inner_first_stage_data_reg[1614]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1613_ ( .D(N9188), .CP(clk), 
        .Q(inner_first_stage_data_reg[1613]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1612_ ( .D(N9187), .CP(clk), 
        .Q(inner_first_stage_data_reg[1612]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1611_ ( .D(N9186), .CP(clk), 
        .Q(inner_first_stage_data_reg[1611]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1610_ ( .D(N9185), .CP(clk), 
        .Q(inner_first_stage_data_reg[1610]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1609_ ( .D(N9184), .CP(clk), 
        .Q(inner_first_stage_data_reg[1609]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1608_ ( .D(N9183), .CP(clk), 
        .Q(inner_first_stage_data_reg[1608]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1607_ ( .D(N9182), .CP(clk), 
        .Q(inner_first_stage_data_reg[1607]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1606_ ( .D(N9181), .CP(clk), 
        .Q(inner_first_stage_data_reg[1606]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1605_ ( .D(N9180), .CP(clk), 
        .Q(inner_first_stage_data_reg[1605]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1604_ ( .D(N9179), .CP(clk), 
        .Q(inner_first_stage_data_reg[1604]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1603_ ( .D(N9178), .CP(clk), 
        .Q(inner_first_stage_data_reg[1603]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1602_ ( .D(N9177), .CP(clk), 
        .Q(inner_first_stage_data_reg[1602]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1601_ ( .D(N9176), .CP(clk), 
        .Q(inner_first_stage_data_reg[1601]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1600_ ( .D(N9175), .CP(clk), 
        .Q(inner_first_stage_data_reg[1600]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_51_ ( .D(N9390), .CP(clk), 
        .Q(inner_first_stage_valid_reg[51]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1663_ ( .D(N9422), .CP(clk), 
        .Q(inner_first_stage_data_reg[1663]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1662_ ( .D(N9421), .CP(clk), 
        .Q(inner_first_stage_data_reg[1662]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1661_ ( .D(N9420), .CP(clk), 
        .Q(inner_first_stage_data_reg[1661]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1660_ ( .D(N9419), .CP(clk), 
        .Q(inner_first_stage_data_reg[1660]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1659_ ( .D(N9418), .CP(clk), 
        .Q(inner_first_stage_data_reg[1659]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1658_ ( .D(N9417), .CP(clk), 
        .Q(inner_first_stage_data_reg[1658]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1657_ ( .D(N9416), .CP(clk), 
        .Q(inner_first_stage_data_reg[1657]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1656_ ( .D(N9415), .CP(clk), 
        .Q(inner_first_stage_data_reg[1656]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1655_ ( .D(N9414), .CP(clk), 
        .Q(inner_first_stage_data_reg[1655]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1654_ ( .D(N9413), .CP(clk), 
        .Q(inner_first_stage_data_reg[1654]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1653_ ( .D(N9412), .CP(clk), 
        .Q(inner_first_stage_data_reg[1653]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1652_ ( .D(N9411), .CP(clk), 
        .Q(inner_first_stage_data_reg[1652]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1651_ ( .D(N9410), .CP(clk), 
        .Q(inner_first_stage_data_reg[1651]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1650_ ( .D(N9409), .CP(clk), 
        .Q(inner_first_stage_data_reg[1650]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1649_ ( .D(N9408), .CP(clk), 
        .Q(inner_first_stage_data_reg[1649]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1648_ ( .D(N9407), .CP(clk), 
        .Q(inner_first_stage_data_reg[1648]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1647_ ( .D(N9406), .CP(clk), 
        .Q(inner_first_stage_data_reg[1647]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1646_ ( .D(N9405), .CP(clk), 
        .Q(inner_first_stage_data_reg[1646]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1645_ ( .D(N9404), .CP(clk), 
        .Q(inner_first_stage_data_reg[1645]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1644_ ( .D(N9403), .CP(clk), 
        .Q(inner_first_stage_data_reg[1644]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1643_ ( .D(N9402), .CP(clk), 
        .Q(inner_first_stage_data_reg[1643]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1642_ ( .D(N9401), .CP(clk), 
        .Q(inner_first_stage_data_reg[1642]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1641_ ( .D(N9400), .CP(clk), 
        .Q(inner_first_stage_data_reg[1641]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1640_ ( .D(N9399), .CP(clk), 
        .Q(inner_first_stage_data_reg[1640]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1639_ ( .D(N9398), .CP(clk), 
        .Q(inner_first_stage_data_reg[1639]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1638_ ( .D(N9397), .CP(clk), 
        .Q(inner_first_stage_data_reg[1638]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1637_ ( .D(N9396), .CP(clk), 
        .Q(inner_first_stage_data_reg[1637]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1636_ ( .D(N9395), .CP(clk), 
        .Q(inner_first_stage_data_reg[1636]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1635_ ( .D(N9394), .CP(clk), 
        .Q(inner_first_stage_data_reg[1635]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1634_ ( .D(N9393), .CP(clk), 
        .Q(inner_first_stage_data_reg[1634]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1633_ ( .D(N9392), .CP(clk), 
        .Q(inner_first_stage_data_reg[1633]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1632_ ( .D(N9391), .CP(clk), 
        .Q(inner_first_stage_data_reg[1632]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_52_ ( .D(N9606), .CP(clk), 
        .Q(inner_first_stage_valid_reg[52]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1695_ ( .D(N9638), .CP(clk), 
        .Q(inner_first_stage_data_reg[1695]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1694_ ( .D(N9637), .CP(clk), 
        .Q(inner_first_stage_data_reg[1694]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1693_ ( .D(N9636), .CP(clk), 
        .Q(inner_first_stage_data_reg[1693]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1692_ ( .D(N9635), .CP(clk), 
        .Q(inner_first_stage_data_reg[1692]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1691_ ( .D(N9634), .CP(clk), 
        .Q(inner_first_stage_data_reg[1691]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1690_ ( .D(N9633), .CP(clk), 
        .Q(inner_first_stage_data_reg[1690]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1689_ ( .D(N9632), .CP(clk), 
        .Q(inner_first_stage_data_reg[1689]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1688_ ( .D(N9631), .CP(clk), 
        .Q(inner_first_stage_data_reg[1688]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1687_ ( .D(N9630), .CP(clk), 
        .Q(inner_first_stage_data_reg[1687]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1686_ ( .D(N9629), .CP(clk), 
        .Q(inner_first_stage_data_reg[1686]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1685_ ( .D(N9628), .CP(clk), 
        .Q(inner_first_stage_data_reg[1685]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1684_ ( .D(N9627), .CP(clk), 
        .Q(inner_first_stage_data_reg[1684]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1683_ ( .D(N9626), .CP(clk), 
        .Q(inner_first_stage_data_reg[1683]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1682_ ( .D(N9625), .CP(clk), 
        .Q(inner_first_stage_data_reg[1682]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1681_ ( .D(N9624), .CP(clk), 
        .Q(inner_first_stage_data_reg[1681]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1680_ ( .D(N9623), .CP(clk), 
        .Q(inner_first_stage_data_reg[1680]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1679_ ( .D(N9622), .CP(clk), 
        .Q(inner_first_stage_data_reg[1679]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1678_ ( .D(N9621), .CP(clk), 
        .Q(inner_first_stage_data_reg[1678]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1677_ ( .D(N9620), .CP(clk), 
        .Q(inner_first_stage_data_reg[1677]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1676_ ( .D(N9619), .CP(clk), 
        .Q(inner_first_stage_data_reg[1676]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1675_ ( .D(N9618), .CP(clk), 
        .Q(inner_first_stage_data_reg[1675]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1674_ ( .D(N9617), .CP(clk), 
        .Q(inner_first_stage_data_reg[1674]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1673_ ( .D(N9616), .CP(clk), 
        .Q(inner_first_stage_data_reg[1673]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1672_ ( .D(N9615), .CP(clk), 
        .Q(inner_first_stage_data_reg[1672]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1671_ ( .D(N9614), .CP(clk), 
        .Q(inner_first_stage_data_reg[1671]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1670_ ( .D(N9613), .CP(clk), 
        .Q(inner_first_stage_data_reg[1670]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1669_ ( .D(N9612), .CP(clk), 
        .Q(inner_first_stage_data_reg[1669]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1668_ ( .D(N9611), .CP(clk), 
        .Q(inner_first_stage_data_reg[1668]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1667_ ( .D(N9610), .CP(clk), 
        .Q(inner_first_stage_data_reg[1667]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1666_ ( .D(N9609), .CP(clk), 
        .Q(inner_first_stage_data_reg[1666]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1665_ ( .D(N9608), .CP(clk), 
        .Q(inner_first_stage_data_reg[1665]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1664_ ( .D(N9607), .CP(clk), 
        .Q(inner_first_stage_data_reg[1664]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_53_ ( .D(N9822), .CP(clk), 
        .Q(inner_first_stage_valid_reg[53]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1727_ ( .D(N9854), .CP(clk), 
        .Q(inner_first_stage_data_reg[1727]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1726_ ( .D(N9853), .CP(clk), 
        .Q(inner_first_stage_data_reg[1726]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1725_ ( .D(N9852), .CP(clk), 
        .Q(inner_first_stage_data_reg[1725]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1724_ ( .D(N9851), .CP(clk), 
        .Q(inner_first_stage_data_reg[1724]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1723_ ( .D(N9850), .CP(clk), 
        .Q(inner_first_stage_data_reg[1723]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1722_ ( .D(N9849), .CP(clk), 
        .Q(inner_first_stage_data_reg[1722]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1721_ ( .D(N9848), .CP(clk), 
        .Q(inner_first_stage_data_reg[1721]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1720_ ( .D(N9847), .CP(clk), 
        .Q(inner_first_stage_data_reg[1720]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1719_ ( .D(N9846), .CP(clk), 
        .Q(inner_first_stage_data_reg[1719]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1718_ ( .D(N9845), .CP(clk), 
        .Q(inner_first_stage_data_reg[1718]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1717_ ( .D(N9844), .CP(clk), 
        .Q(inner_first_stage_data_reg[1717]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1716_ ( .D(N9843), .CP(clk), 
        .Q(inner_first_stage_data_reg[1716]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1715_ ( .D(N9842), .CP(clk), 
        .Q(inner_first_stage_data_reg[1715]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1714_ ( .D(N9841), .CP(clk), 
        .Q(inner_first_stage_data_reg[1714]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1713_ ( .D(N9840), .CP(clk), 
        .Q(inner_first_stage_data_reg[1713]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1712_ ( .D(N9839), .CP(clk), 
        .Q(inner_first_stage_data_reg[1712]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1711_ ( .D(N9838), .CP(clk), 
        .Q(inner_first_stage_data_reg[1711]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1710_ ( .D(N9837), .CP(clk), 
        .Q(inner_first_stage_data_reg[1710]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1709_ ( .D(N9836), .CP(clk), 
        .Q(inner_first_stage_data_reg[1709]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1708_ ( .D(N9835), .CP(clk), 
        .Q(inner_first_stage_data_reg[1708]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1707_ ( .D(N9834), .CP(clk), 
        .Q(inner_first_stage_data_reg[1707]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1706_ ( .D(N9833), .CP(clk), 
        .Q(inner_first_stage_data_reg[1706]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1705_ ( .D(N9832), .CP(clk), 
        .Q(inner_first_stage_data_reg[1705]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1704_ ( .D(N9831), .CP(clk), 
        .Q(inner_first_stage_data_reg[1704]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1703_ ( .D(N9830), .CP(clk), 
        .Q(inner_first_stage_data_reg[1703]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1702_ ( .D(N9829), .CP(clk), 
        .Q(inner_first_stage_data_reg[1702]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1701_ ( .D(N9828), .CP(clk), 
        .Q(inner_first_stage_data_reg[1701]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1700_ ( .D(N9827), .CP(clk), 
        .Q(inner_first_stage_data_reg[1700]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1699_ ( .D(N9826), .CP(clk), 
        .Q(inner_first_stage_data_reg[1699]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1698_ ( .D(N9825), .CP(clk), 
        .Q(inner_first_stage_data_reg[1698]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1697_ ( .D(N9824), .CP(clk), 
        .Q(inner_first_stage_data_reg[1697]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1696_ ( .D(N9823), .CP(clk), 
        .Q(inner_first_stage_data_reg[1696]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_54_ ( .D(N10038), .CP(clk), 
        .Q(inner_first_stage_valid_reg[54]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1759_ ( .D(N10070), .CP(clk), .Q(inner_first_stage_data_reg[1759]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1758_ ( .D(N10069), .CP(clk), .Q(inner_first_stage_data_reg[1758]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1757_ ( .D(N10068), .CP(clk), .Q(inner_first_stage_data_reg[1757]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1756_ ( .D(N10067), .CP(clk), .Q(inner_first_stage_data_reg[1756]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1755_ ( .D(N10066), .CP(clk), .Q(inner_first_stage_data_reg[1755]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1754_ ( .D(N10065), .CP(clk), .Q(inner_first_stage_data_reg[1754]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1753_ ( .D(N10064), .CP(clk), .Q(inner_first_stage_data_reg[1753]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1752_ ( .D(N10063), .CP(clk), .Q(inner_first_stage_data_reg[1752]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1751_ ( .D(N10062), .CP(clk), .Q(inner_first_stage_data_reg[1751]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1750_ ( .D(N10061), .CP(clk), .Q(inner_first_stage_data_reg[1750]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1749_ ( .D(N10060), .CP(clk), .Q(inner_first_stage_data_reg[1749]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1748_ ( .D(N10059), .CP(clk), .Q(inner_first_stage_data_reg[1748]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1747_ ( .D(N10058), .CP(clk), .Q(inner_first_stage_data_reg[1747]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1746_ ( .D(N10057), .CP(clk), .Q(inner_first_stage_data_reg[1746]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1745_ ( .D(N10056), .CP(clk), .Q(inner_first_stage_data_reg[1745]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1744_ ( .D(N10055), .CP(clk), .Q(inner_first_stage_data_reg[1744]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1743_ ( .D(N10054), .CP(clk), .Q(inner_first_stage_data_reg[1743]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1742_ ( .D(N10053), .CP(clk), .Q(inner_first_stage_data_reg[1742]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1741_ ( .D(N10052), .CP(clk), .Q(inner_first_stage_data_reg[1741]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1740_ ( .D(N10051), .CP(clk), .Q(inner_first_stage_data_reg[1740]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1739_ ( .D(N10050), .CP(clk), .Q(inner_first_stage_data_reg[1739]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1738_ ( .D(N10049), .CP(clk), .Q(inner_first_stage_data_reg[1738]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1737_ ( .D(N10048), .CP(clk), .Q(inner_first_stage_data_reg[1737]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1736_ ( .D(N10047), .CP(clk), .Q(inner_first_stage_data_reg[1736]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1735_ ( .D(N10046), .CP(clk), .Q(inner_first_stage_data_reg[1735]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1734_ ( .D(N10045), .CP(clk), .Q(inner_first_stage_data_reg[1734]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1733_ ( .D(N10044), .CP(clk), .Q(inner_first_stage_data_reg[1733]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1732_ ( .D(N10043), .CP(clk), .Q(inner_first_stage_data_reg[1732]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1731_ ( .D(N10042), .CP(clk), .Q(inner_first_stage_data_reg[1731]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1730_ ( .D(N10041), .CP(clk), .Q(inner_first_stage_data_reg[1730]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1729_ ( .D(N10040), .CP(clk), .Q(inner_first_stage_data_reg[1729]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1728_ ( .D(N10039), .CP(clk), .Q(inner_first_stage_data_reg[1728]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_55_ ( .D(N10254), .CP(clk), 
        .Q(inner_first_stage_valid_reg[55]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1791_ ( .D(N10286), .CP(clk), .Q(inner_first_stage_data_reg[1791]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1790_ ( .D(N10285), .CP(clk), .Q(inner_first_stage_data_reg[1790]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1789_ ( .D(N10284), .CP(clk), .Q(inner_first_stage_data_reg[1789]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1788_ ( .D(N10283), .CP(clk), .Q(inner_first_stage_data_reg[1788]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1787_ ( .D(N10282), .CP(clk), .Q(inner_first_stage_data_reg[1787]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1786_ ( .D(N10281), .CP(clk), .Q(inner_first_stage_data_reg[1786]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1785_ ( .D(N10280), .CP(clk), .Q(inner_first_stage_data_reg[1785]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1784_ ( .D(N10279), .CP(clk), .Q(inner_first_stage_data_reg[1784]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1783_ ( .D(N10278), .CP(clk), .Q(inner_first_stage_data_reg[1783]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1782_ ( .D(N10277), .CP(clk), .Q(inner_first_stage_data_reg[1782]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1781_ ( .D(N10276), .CP(clk), .Q(inner_first_stage_data_reg[1781]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1780_ ( .D(N10275), .CP(clk), .Q(inner_first_stage_data_reg[1780]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1779_ ( .D(N10274), .CP(clk), .Q(inner_first_stage_data_reg[1779]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1778_ ( .D(N10273), .CP(clk), .Q(inner_first_stage_data_reg[1778]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1777_ ( .D(N10272), .CP(clk), .Q(inner_first_stage_data_reg[1777]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1776_ ( .D(N10271), .CP(clk), .Q(inner_first_stage_data_reg[1776]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1775_ ( .D(N10270), .CP(clk), .Q(inner_first_stage_data_reg[1775]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1774_ ( .D(N10269), .CP(clk), .Q(inner_first_stage_data_reg[1774]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1773_ ( .D(N10268), .CP(clk), .Q(inner_first_stage_data_reg[1773]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1772_ ( .D(N10267), .CP(clk), .Q(inner_first_stage_data_reg[1772]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1771_ ( .D(N10266), .CP(clk), .Q(inner_first_stage_data_reg[1771]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1770_ ( .D(N10265), .CP(clk), .Q(inner_first_stage_data_reg[1770]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1769_ ( .D(N10264), .CP(clk), .Q(inner_first_stage_data_reg[1769]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1768_ ( .D(N10263), .CP(clk), .Q(inner_first_stage_data_reg[1768]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1767_ ( .D(N10262), .CP(clk), .Q(inner_first_stage_data_reg[1767]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1766_ ( .D(N10261), .CP(clk), .Q(inner_first_stage_data_reg[1766]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1765_ ( .D(N10260), .CP(clk), .Q(inner_first_stage_data_reg[1765]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1764_ ( .D(N10259), .CP(clk), .Q(inner_first_stage_data_reg[1764]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1763_ ( .D(N10258), .CP(clk), .Q(inner_first_stage_data_reg[1763]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1762_ ( .D(N10257), .CP(clk), .Q(inner_first_stage_data_reg[1762]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1761_ ( .D(N10256), .CP(clk), .Q(inner_first_stage_data_reg[1761]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1760_ ( .D(N10255), .CP(clk), .Q(inner_first_stage_data_reg[1760]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_56_ ( .D(N10488), .CP(clk), 
        .Q(inner_first_stage_valid_reg[56]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1823_ ( .D(N10520), .CP(clk), .Q(inner_first_stage_data_reg[1823]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1822_ ( .D(N10519), .CP(clk), .Q(inner_first_stage_data_reg[1822]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1821_ ( .D(N10518), .CP(clk), .Q(inner_first_stage_data_reg[1821]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1820_ ( .D(N10517), .CP(clk), .Q(inner_first_stage_data_reg[1820]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1819_ ( .D(N10516), .CP(clk), .Q(inner_first_stage_data_reg[1819]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1818_ ( .D(N10515), .CP(clk), .Q(inner_first_stage_data_reg[1818]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1817_ ( .D(N10514), .CP(clk), .Q(inner_first_stage_data_reg[1817]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1816_ ( .D(N10513), .CP(clk), .Q(inner_first_stage_data_reg[1816]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1815_ ( .D(N10512), .CP(clk), .Q(inner_first_stage_data_reg[1815]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1814_ ( .D(N10511), .CP(clk), .Q(inner_first_stage_data_reg[1814]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1813_ ( .D(N10510), .CP(clk), .Q(inner_first_stage_data_reg[1813]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1812_ ( .D(N10509), .CP(clk), .Q(inner_first_stage_data_reg[1812]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1811_ ( .D(N10508), .CP(clk), .Q(inner_first_stage_data_reg[1811]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1810_ ( .D(N10507), .CP(clk), .Q(inner_first_stage_data_reg[1810]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1809_ ( .D(N10506), .CP(clk), .Q(inner_first_stage_data_reg[1809]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1808_ ( .D(N10505), .CP(clk), .Q(inner_first_stage_data_reg[1808]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1807_ ( .D(N10504), .CP(clk), .Q(inner_first_stage_data_reg[1807]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1806_ ( .D(N10503), .CP(clk), .Q(inner_first_stage_data_reg[1806]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1805_ ( .D(N10502), .CP(clk), .Q(inner_first_stage_data_reg[1805]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1804_ ( .D(N10501), .CP(clk), .Q(inner_first_stage_data_reg[1804]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1803_ ( .D(N10500), .CP(clk), .Q(inner_first_stage_data_reg[1803]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1802_ ( .D(N10499), .CP(clk), .Q(inner_first_stage_data_reg[1802]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1801_ ( .D(N10498), .CP(clk), .Q(inner_first_stage_data_reg[1801]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1800_ ( .D(N10497), .CP(clk), .Q(inner_first_stage_data_reg[1800]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1799_ ( .D(N10496), .CP(clk), .Q(inner_first_stage_data_reg[1799]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1798_ ( .D(N10495), .CP(clk), .Q(inner_first_stage_data_reg[1798]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1797_ ( .D(N10494), .CP(clk), .Q(inner_first_stage_data_reg[1797]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1796_ ( .D(N10493), .CP(clk), .Q(inner_first_stage_data_reg[1796]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1795_ ( .D(N10492), .CP(clk), .Q(inner_first_stage_data_reg[1795]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1794_ ( .D(N10491), .CP(clk), .Q(inner_first_stage_data_reg[1794]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1793_ ( .D(N10490), .CP(clk), .Q(inner_first_stage_data_reg[1793]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1792_ ( .D(N10489), .CP(clk), .Q(inner_first_stage_data_reg[1792]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_57_ ( .D(N10576), .CP(clk), 
        .Q(inner_first_stage_valid_reg[57]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1855_ ( .D(N10608), .CP(clk), .Q(inner_first_stage_data_reg[1855]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1854_ ( .D(N10607), .CP(clk), .Q(inner_first_stage_data_reg[1854]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1853_ ( .D(N10606), .CP(clk), .Q(inner_first_stage_data_reg[1853]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1852_ ( .D(N10605), .CP(clk), .Q(inner_first_stage_data_reg[1852]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1851_ ( .D(N10604), .CP(clk), .Q(inner_first_stage_data_reg[1851]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1850_ ( .D(N10603), .CP(clk), .Q(inner_first_stage_data_reg[1850]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1849_ ( .D(N10602), .CP(clk), .Q(inner_first_stage_data_reg[1849]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1848_ ( .D(N10601), .CP(clk), .Q(inner_first_stage_data_reg[1848]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1847_ ( .D(N10600), .CP(clk), .Q(inner_first_stage_data_reg[1847]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1846_ ( .D(N10599), .CP(clk), .Q(inner_first_stage_data_reg[1846]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1845_ ( .D(N10598), .CP(clk), .Q(inner_first_stage_data_reg[1845]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1844_ ( .D(N10597), .CP(clk), .Q(inner_first_stage_data_reg[1844]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1843_ ( .D(N10596), .CP(clk), .Q(inner_first_stage_data_reg[1843]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1842_ ( .D(N10595), .CP(clk), .Q(inner_first_stage_data_reg[1842]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1841_ ( .D(N10594), .CP(clk), .Q(inner_first_stage_data_reg[1841]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1840_ ( .D(N10593), .CP(clk), .Q(inner_first_stage_data_reg[1840]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1839_ ( .D(N10592), .CP(clk), .Q(inner_first_stage_data_reg[1839]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1838_ ( .D(N10591), .CP(clk), .Q(inner_first_stage_data_reg[1838]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1837_ ( .D(N10590), .CP(clk), .Q(inner_first_stage_data_reg[1837]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1836_ ( .D(N10589), .CP(clk), .Q(inner_first_stage_data_reg[1836]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1835_ ( .D(N10588), .CP(clk), .Q(inner_first_stage_data_reg[1835]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1834_ ( .D(N10587), .CP(clk), .Q(inner_first_stage_data_reg[1834]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1833_ ( .D(N10586), .CP(clk), .Q(inner_first_stage_data_reg[1833]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1832_ ( .D(N10585), .CP(clk), .Q(inner_first_stage_data_reg[1832]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1831_ ( .D(N10584), .CP(clk), .Q(inner_first_stage_data_reg[1831]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1830_ ( .D(N10583), .CP(clk), .Q(inner_first_stage_data_reg[1830]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1829_ ( .D(N10582), .CP(clk), .Q(inner_first_stage_data_reg[1829]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1828_ ( .D(N10581), .CP(clk), .Q(inner_first_stage_data_reg[1828]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1827_ ( .D(N10580), .CP(clk), .Q(inner_first_stage_data_reg[1827]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1826_ ( .D(N10579), .CP(clk), .Q(inner_first_stage_data_reg[1826]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1825_ ( .D(N10578), .CP(clk), .Q(inner_first_stage_data_reg[1825]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1824_ ( .D(N10577), .CP(clk), .Q(inner_first_stage_data_reg[1824]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_58_ ( .D(N10664), .CP(clk), 
        .Q(inner_first_stage_valid_reg[58]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1887_ ( .D(N10696), .CP(clk), .Q(inner_first_stage_data_reg[1887]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1886_ ( .D(N10695), .CP(clk), .Q(inner_first_stage_data_reg[1886]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1885_ ( .D(N10694), .CP(clk), .Q(inner_first_stage_data_reg[1885]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1884_ ( .D(N10693), .CP(clk), .Q(inner_first_stage_data_reg[1884]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1883_ ( .D(N10692), .CP(clk), .Q(inner_first_stage_data_reg[1883]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1882_ ( .D(N10691), .CP(clk), .Q(inner_first_stage_data_reg[1882]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1881_ ( .D(N10690), .CP(clk), .Q(inner_first_stage_data_reg[1881]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1880_ ( .D(N10689), .CP(clk), .Q(inner_first_stage_data_reg[1880]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1879_ ( .D(N10688), .CP(clk), .Q(inner_first_stage_data_reg[1879]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1878_ ( .D(N10687), .CP(clk), .Q(inner_first_stage_data_reg[1878]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1877_ ( .D(N10686), .CP(clk), .Q(inner_first_stage_data_reg[1877]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1876_ ( .D(N10685), .CP(clk), .Q(inner_first_stage_data_reg[1876]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1875_ ( .D(N10684), .CP(clk), .Q(inner_first_stage_data_reg[1875]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1874_ ( .D(N10683), .CP(clk), .Q(inner_first_stage_data_reg[1874]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1873_ ( .D(N10682), .CP(clk), .Q(inner_first_stage_data_reg[1873]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1872_ ( .D(N10681), .CP(clk), .Q(inner_first_stage_data_reg[1872]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1871_ ( .D(N10680), .CP(clk), .Q(inner_first_stage_data_reg[1871]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1870_ ( .D(N10679), .CP(clk), .Q(inner_first_stage_data_reg[1870]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1869_ ( .D(N10678), .CP(clk), .Q(inner_first_stage_data_reg[1869]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1868_ ( .D(N10677), .CP(clk), .Q(inner_first_stage_data_reg[1868]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1867_ ( .D(N10676), .CP(clk), .Q(inner_first_stage_data_reg[1867]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1866_ ( .D(N10675), .CP(clk), .Q(inner_first_stage_data_reg[1866]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1865_ ( .D(N10674), .CP(clk), .Q(inner_first_stage_data_reg[1865]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1864_ ( .D(N10673), .CP(clk), .Q(inner_first_stage_data_reg[1864]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1863_ ( .D(N10672), .CP(clk), .Q(inner_first_stage_data_reg[1863]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1862_ ( .D(N10671), .CP(clk), .Q(inner_first_stage_data_reg[1862]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1861_ ( .D(N10670), .CP(clk), .Q(inner_first_stage_data_reg[1861]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1860_ ( .D(N10669), .CP(clk), .Q(inner_first_stage_data_reg[1860]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1859_ ( .D(N10668), .CP(clk), .Q(inner_first_stage_data_reg[1859]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1858_ ( .D(N10667), .CP(clk), .Q(inner_first_stage_data_reg[1858]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1857_ ( .D(N10666), .CP(clk), .Q(inner_first_stage_data_reg[1857]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1856_ ( .D(N10665), .CP(clk), .Q(inner_first_stage_data_reg[1856]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_59_ ( .D(N10752), .CP(clk), 
        .Q(inner_first_stage_valid_reg[59]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1919_ ( .D(N10784), .CP(clk), .Q(inner_first_stage_data_reg[1919]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1918_ ( .D(N10783), .CP(clk), .Q(inner_first_stage_data_reg[1918]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1917_ ( .D(N10782), .CP(clk), .Q(inner_first_stage_data_reg[1917]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1916_ ( .D(N10781), .CP(clk), .Q(inner_first_stage_data_reg[1916]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1915_ ( .D(N10780), .CP(clk), .Q(inner_first_stage_data_reg[1915]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1914_ ( .D(N10779), .CP(clk), .Q(inner_first_stage_data_reg[1914]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1913_ ( .D(N10778), .CP(clk), .Q(inner_first_stage_data_reg[1913]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1912_ ( .D(N10777), .CP(clk), .Q(inner_first_stage_data_reg[1912]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1911_ ( .D(N10776), .CP(clk), .Q(inner_first_stage_data_reg[1911]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1910_ ( .D(N10775), .CP(clk), .Q(inner_first_stage_data_reg[1910]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1909_ ( .D(N10774), .CP(clk), .Q(inner_first_stage_data_reg[1909]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1908_ ( .D(N10773), .CP(clk), .Q(inner_first_stage_data_reg[1908]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1907_ ( .D(N10772), .CP(clk), .Q(inner_first_stage_data_reg[1907]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1906_ ( .D(N10771), .CP(clk), .Q(inner_first_stage_data_reg[1906]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1905_ ( .D(N10770), .CP(clk), .Q(inner_first_stage_data_reg[1905]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1904_ ( .D(N10769), .CP(clk), .Q(inner_first_stage_data_reg[1904]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1903_ ( .D(N10768), .CP(clk), .Q(inner_first_stage_data_reg[1903]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1902_ ( .D(N10767), .CP(clk), .Q(inner_first_stage_data_reg[1902]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1901_ ( .D(N10766), .CP(clk), .Q(inner_first_stage_data_reg[1901]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1900_ ( .D(N10765), .CP(clk), .Q(inner_first_stage_data_reg[1900]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1899_ ( .D(N10764), .CP(clk), .Q(inner_first_stage_data_reg[1899]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1898_ ( .D(N10763), .CP(clk), .Q(inner_first_stage_data_reg[1898]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1897_ ( .D(N10762), .CP(clk), .Q(inner_first_stage_data_reg[1897]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1896_ ( .D(N10761), .CP(clk), .Q(inner_first_stage_data_reg[1896]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1895_ ( .D(N10760), .CP(clk), .Q(inner_first_stage_data_reg[1895]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1894_ ( .D(N10759), .CP(clk), .Q(inner_first_stage_data_reg[1894]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1893_ ( .D(N10758), .CP(clk), .Q(inner_first_stage_data_reg[1893]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1892_ ( .D(N10757), .CP(clk), .Q(inner_first_stage_data_reg[1892]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1891_ ( .D(N10756), .CP(clk), .Q(inner_first_stage_data_reg[1891]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1890_ ( .D(N10755), .CP(clk), .Q(inner_first_stage_data_reg[1890]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1889_ ( .D(N10754), .CP(clk), .Q(inner_first_stage_data_reg[1889]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1888_ ( .D(N10753), .CP(clk), .Q(inner_first_stage_data_reg[1888]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_60_ ( .D(N10840), .CP(clk), 
        .Q(inner_first_stage_valid_reg[60]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1951_ ( .D(N10872), .CP(clk), .Q(inner_first_stage_data_reg[1951]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1950_ ( .D(N10871), .CP(clk), .Q(inner_first_stage_data_reg[1950]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1949_ ( .D(N10870), .CP(clk), .Q(inner_first_stage_data_reg[1949]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1948_ ( .D(N10869), .CP(clk), .Q(inner_first_stage_data_reg[1948]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1947_ ( .D(N10868), .CP(clk), .Q(inner_first_stage_data_reg[1947]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1946_ ( .D(N10867), .CP(clk), .Q(inner_first_stage_data_reg[1946]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1945_ ( .D(N10866), .CP(clk), .Q(inner_first_stage_data_reg[1945]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1944_ ( .D(N10865), .CP(clk), .Q(inner_first_stage_data_reg[1944]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1943_ ( .D(N10864), .CP(clk), .Q(inner_first_stage_data_reg[1943]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1942_ ( .D(N10863), .CP(clk), .Q(inner_first_stage_data_reg[1942]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1941_ ( .D(N10862), .CP(clk), .Q(inner_first_stage_data_reg[1941]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1940_ ( .D(N10861), .CP(clk), .Q(inner_first_stage_data_reg[1940]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1939_ ( .D(N10860), .CP(clk), .Q(inner_first_stage_data_reg[1939]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1938_ ( .D(N10859), .CP(clk), .Q(inner_first_stage_data_reg[1938]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1937_ ( .D(N10858), .CP(clk), .Q(inner_first_stage_data_reg[1937]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1936_ ( .D(N10857), .CP(clk), .Q(inner_first_stage_data_reg[1936]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1935_ ( .D(N10856), .CP(clk), .Q(inner_first_stage_data_reg[1935]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1934_ ( .D(N10855), .CP(clk), .Q(inner_first_stage_data_reg[1934]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1933_ ( .D(N10854), .CP(clk), .Q(inner_first_stage_data_reg[1933]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1932_ ( .D(N10853), .CP(clk), .Q(inner_first_stage_data_reg[1932]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1931_ ( .D(N10852), .CP(clk), .Q(inner_first_stage_data_reg[1931]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1930_ ( .D(N10851), .CP(clk), .Q(inner_first_stage_data_reg[1930]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1929_ ( .D(N10850), .CP(clk), .Q(inner_first_stage_data_reg[1929]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1928_ ( .D(N10849), .CP(clk), .Q(inner_first_stage_data_reg[1928]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1927_ ( .D(N10848), .CP(clk), .Q(inner_first_stage_data_reg[1927]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1926_ ( .D(N10847), .CP(clk), .Q(inner_first_stage_data_reg[1926]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1925_ ( .D(N10846), .CP(clk), .Q(inner_first_stage_data_reg[1925]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1924_ ( .D(N10845), .CP(clk), .Q(inner_first_stage_data_reg[1924]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1923_ ( .D(N10844), .CP(clk), .Q(inner_first_stage_data_reg[1923]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1922_ ( .D(N10843), .CP(clk), .Q(inner_first_stage_data_reg[1922]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1921_ ( .D(N10842), .CP(clk), .Q(inner_first_stage_data_reg[1921]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1920_ ( .D(N10841), .CP(clk), .Q(inner_first_stage_data_reg[1920]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_61_ ( .D(N10928), .CP(clk), 
        .Q(inner_first_stage_valid_reg[61]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1983_ ( .D(N10960), .CP(clk), .Q(inner_first_stage_data_reg[1983]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1982_ ( .D(N10959), .CP(clk), .Q(inner_first_stage_data_reg[1982]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1981_ ( .D(N10958), .CP(clk), .Q(inner_first_stage_data_reg[1981]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1980_ ( .D(N10957), .CP(clk), .Q(inner_first_stage_data_reg[1980]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1979_ ( .D(N10956), .CP(clk), .Q(inner_first_stage_data_reg[1979]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1978_ ( .D(N10955), .CP(clk), .Q(inner_first_stage_data_reg[1978]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1977_ ( .D(N10954), .CP(clk), .Q(inner_first_stage_data_reg[1977]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1976_ ( .D(N10953), .CP(clk), .Q(inner_first_stage_data_reg[1976]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1975_ ( .D(N10952), .CP(clk), .Q(inner_first_stage_data_reg[1975]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1974_ ( .D(N10951), .CP(clk), .Q(inner_first_stage_data_reg[1974]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1973_ ( .D(N10950), .CP(clk), .Q(inner_first_stage_data_reg[1973]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1972_ ( .D(N10949), .CP(clk), .Q(inner_first_stage_data_reg[1972]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1971_ ( .D(N10948), .CP(clk), .Q(inner_first_stage_data_reg[1971]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1970_ ( .D(N10947), .CP(clk), .Q(inner_first_stage_data_reg[1970]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1969_ ( .D(N10946), .CP(clk), .Q(inner_first_stage_data_reg[1969]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1968_ ( .D(N10945), .CP(clk), .Q(inner_first_stage_data_reg[1968]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1967_ ( .D(N10944), .CP(clk), .Q(inner_first_stage_data_reg[1967]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1966_ ( .D(N10943), .CP(clk), .Q(inner_first_stage_data_reg[1966]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1965_ ( .D(N10942), .CP(clk), .Q(inner_first_stage_data_reg[1965]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1964_ ( .D(N10941), .CP(clk), .Q(inner_first_stage_data_reg[1964]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1963_ ( .D(N10940), .CP(clk), .Q(inner_first_stage_data_reg[1963]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1962_ ( .D(N10939), .CP(clk), .Q(inner_first_stage_data_reg[1962]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1961_ ( .D(N10938), .CP(clk), .Q(inner_first_stage_data_reg[1961]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1960_ ( .D(N10937), .CP(clk), .Q(inner_first_stage_data_reg[1960]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1959_ ( .D(N10936), .CP(clk), .Q(inner_first_stage_data_reg[1959]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1958_ ( .D(N10935), .CP(clk), .Q(inner_first_stage_data_reg[1958]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1957_ ( .D(N10934), .CP(clk), .Q(inner_first_stage_data_reg[1957]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1956_ ( .D(N10933), .CP(clk), .Q(inner_first_stage_data_reg[1956]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1955_ ( .D(N10932), .CP(clk), .Q(inner_first_stage_data_reg[1955]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1954_ ( .D(N10931), .CP(clk), .Q(inner_first_stage_data_reg[1954]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1953_ ( .D(N10930), .CP(clk), .Q(inner_first_stage_data_reg[1953]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1952_ ( .D(N10929), .CP(clk), .Q(inner_first_stage_data_reg[1952]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_62_ ( .D(N11016), .CP(clk), 
        .Q(inner_first_stage_valid_reg[62]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2015_ ( .D(N11048), .CP(clk), .Q(inner_first_stage_data_reg[2015]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2014_ ( .D(N11047), .CP(clk), .Q(inner_first_stage_data_reg[2014]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2013_ ( .D(N11046), .CP(clk), .Q(inner_first_stage_data_reg[2013]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2012_ ( .D(N11045), .CP(clk), .Q(inner_first_stage_data_reg[2012]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2011_ ( .D(N11044), .CP(clk), .Q(inner_first_stage_data_reg[2011]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2010_ ( .D(N11043), .CP(clk), .Q(inner_first_stage_data_reg[2010]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2009_ ( .D(N11042), .CP(clk), .Q(inner_first_stage_data_reg[2009]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2008_ ( .D(N11041), .CP(clk), .Q(inner_first_stage_data_reg[2008]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2007_ ( .D(N11040), .CP(clk), .Q(inner_first_stage_data_reg[2007]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2006_ ( .D(N11039), .CP(clk), .Q(inner_first_stage_data_reg[2006]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2005_ ( .D(N11038), .CP(clk), .Q(inner_first_stage_data_reg[2005]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2004_ ( .D(N11037), .CP(clk), .Q(inner_first_stage_data_reg[2004]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2003_ ( .D(N11036), .CP(clk), .Q(inner_first_stage_data_reg[2003]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2002_ ( .D(N11035), .CP(clk), .Q(inner_first_stage_data_reg[2002]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2001_ ( .D(N11034), .CP(clk), .Q(inner_first_stage_data_reg[2001]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2000_ ( .D(N11033), .CP(clk), .Q(inner_first_stage_data_reg[2000]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1999_ ( .D(N11032), .CP(clk), .Q(inner_first_stage_data_reg[1999]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1998_ ( .D(N11031), .CP(clk), .Q(inner_first_stage_data_reg[1998]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1997_ ( .D(N11030), .CP(clk), .Q(inner_first_stage_data_reg[1997]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1996_ ( .D(N11029), .CP(clk), .Q(inner_first_stage_data_reg[1996]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1995_ ( .D(N11028), .CP(clk), .Q(inner_first_stage_data_reg[1995]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1994_ ( .D(N11027), .CP(clk), .Q(inner_first_stage_data_reg[1994]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1993_ ( .D(N11026), .CP(clk), .Q(inner_first_stage_data_reg[1993]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1992_ ( .D(N11025), .CP(clk), .Q(inner_first_stage_data_reg[1992]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1991_ ( .D(N11024), .CP(clk), .Q(inner_first_stage_data_reg[1991]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1990_ ( .D(N11023), .CP(clk), .Q(inner_first_stage_data_reg[1990]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1989_ ( .D(N11022), .CP(clk), .Q(inner_first_stage_data_reg[1989]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1988_ ( .D(N11021), .CP(clk), .Q(inner_first_stage_data_reg[1988]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1987_ ( .D(N11020), .CP(clk), .Q(inner_first_stage_data_reg[1987]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1986_ ( .D(N11019), .CP(clk), .Q(inner_first_stage_data_reg[1986]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1985_ ( .D(N11018), .CP(clk), .Q(inner_first_stage_data_reg[1985]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_1984_ ( .D(N11017), .CP(clk), .Q(inner_first_stage_data_reg[1984]) );
  DFQD1BWP30P140LVT inner_first_stage_valid_reg_reg_63_ ( .D(N11104), .CP(clk), 
        .Q(inner_first_stage_valid_reg[63]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2047_ ( .D(N11136), .CP(clk), .Q(inner_first_stage_data_reg[2047]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2046_ ( .D(N11135), .CP(clk), .Q(inner_first_stage_data_reg[2046]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2045_ ( .D(N11134), .CP(clk), .Q(inner_first_stage_data_reg[2045]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2044_ ( .D(N11133), .CP(clk), .Q(inner_first_stage_data_reg[2044]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2043_ ( .D(N11132), .CP(clk), .Q(inner_first_stage_data_reg[2043]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2042_ ( .D(N11131), .CP(clk), .Q(inner_first_stage_data_reg[2042]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2041_ ( .D(N11130), .CP(clk), .Q(inner_first_stage_data_reg[2041]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2040_ ( .D(N11129), .CP(clk), .Q(inner_first_stage_data_reg[2040]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2039_ ( .D(N11128), .CP(clk), .Q(inner_first_stage_data_reg[2039]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2038_ ( .D(N11127), .CP(clk), .Q(inner_first_stage_data_reg[2038]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2037_ ( .D(N11126), .CP(clk), .Q(inner_first_stage_data_reg[2037]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2036_ ( .D(N11125), .CP(clk), .Q(inner_first_stage_data_reg[2036]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2035_ ( .D(N11124), .CP(clk), .Q(inner_first_stage_data_reg[2035]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2034_ ( .D(N11123), .CP(clk), .Q(inner_first_stage_data_reg[2034]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2033_ ( .D(N11122), .CP(clk), .Q(inner_first_stage_data_reg[2033]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2032_ ( .D(N11121), .CP(clk), .Q(inner_first_stage_data_reg[2032]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2031_ ( .D(N11120), .CP(clk), .Q(inner_first_stage_data_reg[2031]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2030_ ( .D(N11119), .CP(clk), .Q(inner_first_stage_data_reg[2030]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2029_ ( .D(N11118), .CP(clk), .Q(inner_first_stage_data_reg[2029]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2028_ ( .D(N11117), .CP(clk), .Q(inner_first_stage_data_reg[2028]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2027_ ( .D(N11116), .CP(clk), .Q(inner_first_stage_data_reg[2027]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2026_ ( .D(N11115), .CP(clk), .Q(inner_first_stage_data_reg[2026]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2025_ ( .D(N11114), .CP(clk), .Q(inner_first_stage_data_reg[2025]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2024_ ( .D(N11113), .CP(clk), .Q(inner_first_stage_data_reg[2024]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2023_ ( .D(N11112), .CP(clk), .Q(inner_first_stage_data_reg[2023]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2022_ ( .D(N11111), .CP(clk), .Q(inner_first_stage_data_reg[2022]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2021_ ( .D(N11110), .CP(clk), .Q(inner_first_stage_data_reg[2021]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2020_ ( .D(N11109), .CP(clk), .Q(inner_first_stage_data_reg[2020]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2019_ ( .D(N11108), .CP(clk), .Q(inner_first_stage_data_reg[2019]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2018_ ( .D(N11107), .CP(clk), .Q(inner_first_stage_data_reg[2018]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2017_ ( .D(N11106), .CP(clk), .Q(inner_first_stage_data_reg[2017]) );
  DFQD1BWP30P140LVT inner_first_stage_data_reg_reg_2016_ ( .D(N11105), .CP(clk), .Q(inner_first_stage_data_reg[2016]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_7_ ( .D(N11250), .CP(clk), .Q(o_valid[7])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_6_ ( .D(N10400), .CP(clk), .Q(o_valid[6])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_5_ ( .D(N8526), .CP(clk), .Q(o_valid[5])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_4_ ( .D(N7676), .CP(clk), .Q(o_valid[4])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_3_ ( .D(N5802), .CP(clk), .Q(o_valid[3])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_2_ ( .D(N4952), .CP(clk), .Q(o_valid[2])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_1_ ( .D(N3078), .CP(clk), .Q(o_valid[1])
         );
  DFQD2BWP30P140LVT o_valid_reg_reg_0_ ( .D(N2228), .CP(clk), .Q(o_valid[0])
         );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N11282), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N11281), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N11280), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N11279), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N11278), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N11277), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N11276), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N11275), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N11274), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N11273), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N11272), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N11271), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N11270), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N11269), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N11268), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N11267), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N11266), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N11265), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N11264), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N11263), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N11262), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N11261), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N11260), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N11259), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N11258), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N11257), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N11256), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N11255), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N11254), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N11253), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N11252), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N11251), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N10432), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N10431), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N10430), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N10429), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N10428), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N10427), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N10426), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N10425), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N10424), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N10423), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N10422), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N10421), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N10420), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N10419), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N10418), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N10417), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N10416), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N10415), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N10414), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N10413), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N10412), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N10411), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N10410), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N10409), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N10408), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N10407), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N10406), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N10405), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N10404), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N10403), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N10402), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N10401), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N8558), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N8557), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N8556), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N8555), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N8554), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N8553), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N8552), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N8551), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N8550), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N8549), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N8548), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N8547), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N8546), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N8545), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N8544), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N8543), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N8542), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N8541), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N8540), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N8539), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N8538), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N8537), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N8536), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N8535), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N8534), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N8533), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N8532), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N8531), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N8530), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N8529), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N8528), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N8527), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N7708), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N7707), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N7706), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N7705), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N7704), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N7703), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N7702), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N7701), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N7700), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N7699), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N7698), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N7697), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N7696), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N7695), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N7694), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N7693), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N7692), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N7691), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N7690), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N7689), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N7688), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N7687), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N7686), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N7685), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N7684), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N7683), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N7682), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N7681), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N7680), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N7679), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N7678), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N7677), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N5834), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N5833), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N5832), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N5831), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N5830), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N5829), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N5828), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N5827), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N5826), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N5825), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N5824), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N5823), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N5822), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N5821), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N5820), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N5819), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N5818), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N5817), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N5816), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N5815), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N5814), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N5813), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N5812), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N5811), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N5810), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N5809), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N5808), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N5807), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N5806), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N5805), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N5804), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N5803), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N4984), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N4983), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N4982), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N4981), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N4980), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N4979), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N4978), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N4977), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N4976), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N4975), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N4974), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N4973), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N4972), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N4971), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N4970), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N4969), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N4968), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N4967), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N4966), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N4965), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N4964), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N4963), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N4962), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N4961), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N4960), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N4959), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N4958), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N4957), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N4956), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N4955), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N4954), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N4953), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N3110), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N3109), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N3108), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N3107), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N3106), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N3105), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N3104), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N3103), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N3102), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N3101), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N3100), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N3099), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N3098), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N3097), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N3096), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N3095), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N3094), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N3093), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N3092), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N3091), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N3090), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N3089), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N3088), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N3087), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N3086), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N3085), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N3084), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N3083), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N3082), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N3081), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N3080), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N3079), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N2260), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N2259), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N2258), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N2257), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N2256), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N2255), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N2254), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N2253), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N2252), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N2251), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N2250), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N2249), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N2248), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N2247), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N2246), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N2245), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N2244), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N2243), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N2242), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N2241), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N2240), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N2239), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N2238), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N2237), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N2236), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N2235), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N2234), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N2233), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N2232), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N2231), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N2230), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N2229), .CP(clk), .Q(
        o_data_bus[0]) );
  DFKSND1BWP30P140LVT inner_first_stage_valid_reg_reg_39_ ( .D(n12304), .SN(
        n12302), .CP(clk), .Q(n12303), .QN(inner_first_stage_valid_reg[39]) );
  NR3D1P5BWP30P140LVT U8589 ( .A1(inner_first_stage_valid_reg[2]), .A2(
        inner_first_stage_valid_reg[7]), .A3(n8585), .ZN(n11345) );
  INVD1BWP30P140LVT U8590 ( .I(n12302), .ZN(n11057) );
  INVD2BWP30P140LVT U8591 ( .I(n6239), .ZN(n10869) );
  INVD2BWP30P140LVT U8592 ( .I(n10869), .ZN(n11173) );
  NR3D0P7BWP30P140LVT U8593 ( .A1(inner_first_stage_valid_reg[63]), .A2(n8828), 
        .A3(n8827), .ZN(n6211) );
  ND2D1BWP30P140LVT U8594 ( .A1(n10886), .A2(n10884), .ZN(n10885) );
  ND2D1BWP30P140LVT U8595 ( .A1(n10901), .A2(n10902), .ZN(n10899) );
  ND2D1BWP30P140LVT U8596 ( .A1(n10879), .A2(n10877), .ZN(n10871) );
  ND2D1BWP30P140LVT U8597 ( .A1(n12302), .A2(n10872), .ZN(n10876) );
  INR3D1BWP30P140LVT U8598 ( .A1(n10875), .B1(n10874), .B2(n10873), .ZN(n11887) );
  NR2D1BWP30P140LVT U8599 ( .A1(n11173), .A2(inner_first_stage_valid_reg[60]), 
        .ZN(n8825) );
  ND2D1BWP30P140LVT U8600 ( .A1(n10887), .A2(n10882), .ZN(n10891) );
  ND2D1BWP30P140LVT U8601 ( .A1(n12302), .A2(i_valid[1]), .ZN(n10634) );
  ND2D1BWP30P140LVT U8602 ( .A1(n12302), .A2(i_valid[2]), .ZN(n10632) );
  ND2D1BWP30P140LVT U8603 ( .A1(n12302), .A2(i_valid[3]), .ZN(n10630) );
  ND2D1BWP30P140LVT U8604 ( .A1(n12302), .A2(i_valid[9]), .ZN(n10391) );
  ND2D1BWP30P140LVT U8605 ( .A1(n12302), .A2(i_valid[0]), .ZN(n10629) );
  ND2D1BWP30P140LVT U8606 ( .A1(n12302), .A2(i_valid[5]), .ZN(n10664) );
  ND2D1BWP30P140LVT U8607 ( .A1(n12302), .A2(i_valid[4]), .ZN(n10663) );
  ND2D1BWP30P140LVT U8608 ( .A1(n12302), .A2(i_valid[8]), .ZN(n10394) );
  ND2D1BWP30P140LVT U8609 ( .A1(n12302), .A2(i_valid[11]), .ZN(n10392) );
  ND2D1BWP30P140LVT U8610 ( .A1(n12302), .A2(i_valid[7]), .ZN(n10670) );
  ND2D1BWP30P140LVT U8611 ( .A1(n12302), .A2(i_valid[12]), .ZN(n8441) );
  ND2D1BWP30P140LVT U8612 ( .A1(n12302), .A2(i_valid[6]), .ZN(n10667) );
  ND2D1BWP30P140LVT U8613 ( .A1(n12302), .A2(i_valid[10]), .ZN(n10395) );
  ND2D1BWP30P140LVT U8614 ( .A1(n12302), .A2(i_valid[15]), .ZN(n8447) );
  ND2D1BWP30P140LVT U8615 ( .A1(n12302), .A2(i_valid[13]), .ZN(n8445) );
  ND2D1BWP30P140LVT U8616 ( .A1(n12302), .A2(i_valid[14]), .ZN(n8443) );
  ND2D1BWP30P140LVT U8617 ( .A1(n12302), .A2(i_valid[20]), .ZN(n6689) );
  ND2D1BWP30P140LVT U8618 ( .A1(n12302), .A2(i_valid[23]), .ZN(n6690) );
  ND2D1BWP30P140LVT U8619 ( .A1(n12302), .A2(i_valid[22]), .ZN(n6691) );
  ND2D1BWP30P140LVT U8620 ( .A1(n12302), .A2(i_valid[21]), .ZN(n6693) );
  ND2D1BWP30P140LVT U8621 ( .A1(n12302), .A2(i_valid[16]), .ZN(n10691) );
  ND2D1BWP30P140LVT U8622 ( .A1(n12302), .A2(i_valid[17]), .ZN(n10696) );
  ND2D1BWP30P140LVT U8623 ( .A1(n12302), .A2(i_valid[19]), .ZN(n10694) );
  ND2D1BWP30P140LVT U8624 ( .A1(n12302), .A2(i_valid[18]), .ZN(n10692) );
  ND2D1BWP30P140LVT U8625 ( .A1(n12302), .A2(i_valid[31]), .ZN(n7771) );
  ND2D1BWP30P140LVT U8626 ( .A1(n12302), .A2(i_valid[30]), .ZN(n7765) );
  ND2D1BWP30P140LVT U8627 ( .A1(n12302), .A2(i_valid[28]), .ZN(n7767) );
  ND2D1BWP30P140LVT U8628 ( .A1(n12302), .A2(i_valid[27]), .ZN(n7179) );
  ND2D1BWP30P140LVT U8629 ( .A1(n12302), .A2(i_valid[24]), .ZN(n7178) );
  ND2D1BWP30P140LVT U8630 ( .A1(n6228), .A2(i_cmd[226]), .ZN(n7553) );
  ND2D1BWP30P140LVT U8631 ( .A1(n6253), .A2(i_cmd[3]), .ZN(n8541) );
  ND2D1BWP30P140LVT U8632 ( .A1(n6241), .A2(i_cmd[39]), .ZN(n10662) );
  ND2D1BWP30P140LVT U8633 ( .A1(n11040), .A2(i_cmd[36]), .ZN(n11042) );
  ND2D1BWP30P140LVT U8634 ( .A1(n10939), .A2(i_cmd[230]), .ZN(n10941) );
  ND2D1BWP30P140LVT U8635 ( .A1(n10934), .A2(i_cmd[7]), .ZN(n10936) );
  NR2D1BWP30P140LVT U8636 ( .A1(inner_first_stage_valid_reg[44]), .A2(n11057), 
        .ZN(n10902) );
  ND2D1BWP30P140LVT U8637 ( .A1(n12302), .A2(n10889), .ZN(n10892) );
  INVD1BWP30P140LVT U8638 ( .I(inner_first_stage_valid_reg[40]), .ZN(n10907)
         );
  NR2D1BWP30P140LVT U8639 ( .A1(inner_first_stage_valid_reg[23]), .A2(
        inner_first_stage_valid_reg[22]), .ZN(n10889) );
  NR2D1BWP30P140LVT U8640 ( .A1(inner_first_stage_valid_reg[20]), .A2(n11057), 
        .ZN(n10888) );
  NR2D1BWP30P140LVT U8641 ( .A1(i_cmd[228]), .A2(i_cmd[244]), .ZN(n6265) );
  NR2D1BWP30P140LVT U8642 ( .A1(i_cmd[252]), .A2(i_cmd[236]), .ZN(n6266) );
  IND2D1BWP30P140LVT U8643 ( .A1(inner_first_stage_valid_reg[2]), .B1(n8580), 
        .ZN(n8583) );
  INR3D0BWP30P140LVT U8644 ( .A1(n8579), .B1(inner_first_stage_valid_reg[4]), 
        .B2(inner_first_stage_valid_reg[0]), .ZN(n8580) );
  OR2D1BWP30P140LVT U8645 ( .A1(n8583), .A2(inner_first_stage_valid_reg[3]), 
        .Z(n8586) );
  ND2D1BWP30P140LVT U8646 ( .A1(n10856), .A2(n10862), .ZN(n10861) );
  NR2D1BWP30P140LVT U8647 ( .A1(inner_first_stage_valid_reg[12]), .A2(n11181), 
        .ZN(n10856) );
  OR2D1BWP30P140LVT U8648 ( .A1(n10861), .A2(inner_first_stage_valid_reg[8]), 
        .Z(n10857) );
  ND2D1BWP30P140LVT U8649 ( .A1(n10860), .A2(n10859), .ZN(n10864) );
  ND2D1BWP30P140LVT U8650 ( .A1(n10858), .A2(n10859), .ZN(n10865) );
  IND2D1BWP30P140LVT U8651 ( .A1(n10891), .B1(n10888), .ZN(n10883) );
  ND2D1BWP30P140LVT U8652 ( .A1(n7455), .A2(n7454), .ZN(n7456) );
  ND2D1BWP30P140LVT U8653 ( .A1(n7452), .A2(n7454), .ZN(n7453) );
  ND2D1BWP30P140LVT U8654 ( .A1(n7460), .A2(n7459), .ZN(n7461) );
  OR2D1BWP30P140LVT U8655 ( .A1(inner_first_stage_valid_reg[33]), .A2(
        inner_first_stage_valid_reg[37]), .Z(n10878) );
  INVD1BWP30P140LVT U8656 ( .I(inner_first_stage_valid_reg[32]), .ZN(n10877)
         );
  NR2D1BWP30P140LVT U8657 ( .A1(inner_first_stage_valid_reg[42]), .A2(
        inner_first_stage_valid_reg[43]), .ZN(n10904) );
  NR2D1BWP30P140LVT U8658 ( .A1(inner_first_stage_valid_reg[46]), .A2(
        inner_first_stage_valid_reg[47]), .ZN(n10903) );
  ND2D1BWP30P140LVT U8659 ( .A1(n10905), .A2(n10907), .ZN(n10898) );
  ND2D1BWP30P140LVT U8660 ( .A1(n7373), .A2(n7369), .ZN(n7375) );
  NR2D1BWP30P140LVT U8661 ( .A1(inner_first_stage_valid_reg[52]), .A2(n11057), 
        .ZN(n7369) );
  ND2D1BWP30P140LVT U8662 ( .A1(n7378), .A2(n7377), .ZN(n7379) );
  OR2D1BWP30P140LVT U8663 ( .A1(n7375), .A2(inner_first_stage_valid_reg[48]), 
        .Z(n7370) );
  ND2D1BWP30P140LVT U8664 ( .A1(n7371), .A2(n7377), .ZN(n7372) );
  ND2D1BWP30P140LVT U8665 ( .A1(n8828), .A2(n8826), .ZN(n8823) );
  INVD1BWP30P140LVT U8666 ( .I(inner_first_stage_valid_reg[59]), .ZN(n8833) );
  ND2D1BWP30P140LVT U8667 ( .A1(n8834), .A2(n8833), .ZN(n8832) );
  ND2D1BWP30P140LVT U8668 ( .A1(n8825), .A2(n8824), .ZN(n8827) );
  OR2D1BWP30P140LVT U8669 ( .A1(i_cmd[231]), .A2(i_cmd[247]), .Z(n7532) );
  INVD1BWP30P140LVT U8670 ( .I(i_cmd[239]), .ZN(n7530) );
  INVD1BWP30P140LVT U8671 ( .I(i_cmd[255]), .ZN(n7531) );
  OR2D1BWP30P140LVT U8672 ( .A1(i_cmd[199]), .A2(i_cmd[215]), .Z(n6990) );
  OR2D1BWP30P140LVT U8673 ( .A1(i_cmd[183]), .A2(i_cmd[167]), .Z(n6323) );
  OR2D1BWP30P140LVT U8674 ( .A1(i_cmd[151]), .A2(i_cmd[135]), .Z(n10695) );
  INVD1BWP30P140LVT U8675 ( .I(i_cmd[159]), .ZN(n10693) );
  INVD1BWP30P140LVT U8676 ( .I(i_cmd[143]), .ZN(n10697) );
  NR2D1BWP30P140LVT U8677 ( .A1(i_cmd[103]), .A2(i_cmd[119]), .ZN(n6257) );
  OR2D1BWP30P140LVT U8678 ( .A1(i_cmd[71]), .A2(i_cmd[87]), .Z(n8479) );
  OR2D1BWP30P140LVT U8679 ( .A1(i_cmd[39]), .A2(i_cmd[55]), .Z(n10668) );
  OR2D1BWP30P140LVT U8680 ( .A1(i_cmd[23]), .A2(i_cmd[7]), .Z(n10633) );
  INVD1BWP30P140LVT U8681 ( .I(i_cmd[31]), .ZN(n10631) );
  INVD1BWP30P140LVT U8682 ( .I(i_cmd[15]), .ZN(n10635) );
  OR2D1BWP30P140LVT U8683 ( .A1(i_cmd[230]), .A2(i_cmd[246]), .Z(n7560) );
  OR2D1BWP30P140LVT U8684 ( .A1(i_cmd[166]), .A2(i_cmd[182]), .Z(n6370) );
  OR2D1BWP30P140LVT U8685 ( .A1(i_cmd[134]), .A2(i_cmd[150]), .Z(n7867) );
  OR2D1BWP30P140LVT U8686 ( .A1(i_cmd[70]), .A2(i_cmd[86]), .Z(n8472) );
  OR2D1BWP30P140LVT U8687 ( .A1(i_cmd[54]), .A2(i_cmd[38]), .Z(n8320) );
  OR2D1BWP30P140LVT U8688 ( .A1(i_cmd[6]), .A2(i_cmd[22]), .Z(n8487) );
  INVD1BWP30P140LVT U8689 ( .I(i_cmd[14]), .ZN(n8486) );
  INVD1BWP30P140LVT U8690 ( .I(i_cmd[30]), .ZN(n8488) );
  OR2D1BWP30P140LVT U8691 ( .A1(i_cmd[229]), .A2(i_cmd[245]), .Z(n7513) );
  OR2D1BWP30P140LVT U8692 ( .A1(i_cmd[197]), .A2(i_cmd[213]), .Z(n6996) );
  OR2D1BWP30P140LVT U8693 ( .A1(i_cmd[165]), .A2(i_cmd[181]), .Z(n6348) );
  OR2D1BWP30P140LVT U8694 ( .A1(i_cmd[133]), .A2(i_cmd[149]), .Z(n7961) );
  OR2D1BWP30P140LVT U8695 ( .A1(i_cmd[101]), .A2(i_cmd[117]), .Z(n7627) );
  OR2D1BWP30P140LVT U8696 ( .A1(i_cmd[69]), .A2(i_cmd[85]), .Z(n8522) );
  OR2D1BWP30P140LVT U8697 ( .A1(i_cmd[53]), .A2(i_cmd[37]), .Z(n8366) );
  INVD1BWP30P140LVT U8698 ( .I(i_cmd[61]), .ZN(n8365) );
  INVD1BWP30P140LVT U8699 ( .I(i_cmd[45]), .ZN(n8367) );
  OR2D1BWP30P140LVT U8700 ( .A1(i_cmd[5]), .A2(i_cmd[21]), .Z(n8492) );
  INVD1BWP30P140LVT U8701 ( .I(i_cmd[13]), .ZN(n8491) );
  INVD1BWP30P140LVT U8702 ( .I(i_cmd[29]), .ZN(n8493) );
  OR2D1BWP30P140LVT U8703 ( .A1(i_cmd[196]), .A2(i_cmd[212]), .Z(n6341) );
  OR2D1BWP30P140LVT U8704 ( .A1(i_cmd[164]), .A2(i_cmd[180]), .Z(n6285) );
  OR2D1BWP30P140LVT U8705 ( .A1(i_cmd[132]), .A2(i_cmd[148]), .Z(n7914) );
  OR2D1BWP30P140LVT U8706 ( .A1(i_cmd[68]), .A2(i_cmd[84]), .Z(n8692) );
  OR2D1BWP30P140LVT U8707 ( .A1(i_cmd[52]), .A2(i_cmd[36]), .Z(n8243) );
  INVD1BWP30P140LVT U8708 ( .I(i_cmd[60]), .ZN(n8242) );
  INVD1BWP30P140LVT U8709 ( .I(i_cmd[44]), .ZN(n8244) );
  OR2D1BWP30P140LVT U8710 ( .A1(i_cmd[4]), .A2(i_cmd[20]), .Z(n8929) );
  OR2D1BWP30P140LVT U8711 ( .A1(i_cmd[227]), .A2(i_cmd[243]), .Z(n7484) );
  OR2D1BWP30P140LVT U8712 ( .A1(i_cmd[195]), .A2(i_cmd[211]), .Z(n6418) );
  OR2D1BWP30P140LVT U8713 ( .A1(i_cmd[163]), .A2(i_cmd[179]), .Z(n6357) );
  OR2D1BWP30P140LVT U8714 ( .A1(i_cmd[131]), .A2(i_cmd[147]), .Z(n7870) );
  OR2D1BWP30P140LVT U8715 ( .A1(i_cmd[115]), .A2(i_cmd[99]), .Z(n7586) );
  OR2D1BWP30P140LVT U8716 ( .A1(i_cmd[67]), .A2(i_cmd[83]), .Z(n8496) );
  OR2D1BWP30P140LVT U8717 ( .A1(i_cmd[35]), .A2(i_cmd[51]), .Z(n8534) );
  OR2D1BWP30P140LVT U8718 ( .A1(i_cmd[3]), .A2(i_cmd[19]), .Z(n8538) );
  OR2D1BWP30P140LVT U8719 ( .A1(i_cmd[226]), .A2(i_cmd[242]), .Z(n7554) );
  OR2D1BWP30P140LVT U8720 ( .A1(i_cmd[194]), .A2(i_cmd[210]), .Z(n7020) );
  OR2D1BWP30P140LVT U8721 ( .A1(i_cmd[146]), .A2(i_cmd[130]), .Z(n7831) );
  OR2D1BWP30P140LVT U8722 ( .A1(i_cmd[98]), .A2(i_cmd[114]), .Z(n7842) );
  OR2D1BWP30P140LVT U8723 ( .A1(i_cmd[66]), .A2(i_cmd[82]), .Z(n8567) );
  OR2D1BWP30P140LVT U8724 ( .A1(i_cmd[50]), .A2(i_cmd[34]), .Z(n8279) );
  OR2D1BWP30P140LVT U8725 ( .A1(i_cmd[18]), .A2(i_cmd[2]), .Z(n8503) );
  OR2D1BWP30P140LVT U8726 ( .A1(i_cmd[225]), .A2(i_cmd[241]), .Z(n7583) );
  OR2D1BWP30P140LVT U8727 ( .A1(i_cmd[193]), .A2(i_cmd[209]), .Z(n7025) );
  OR2D1BWP30P140LVT U8728 ( .A1(i_cmd[129]), .A2(i_cmd[145]), .Z(n7978) );
  OR2D1BWP30P140LVT U8729 ( .A1(i_cmd[81]), .A2(i_cmd[65]), .Z(n8526) );
  INVD1BWP30P140LVT U8730 ( .I(i_cmd[89]), .ZN(n8525) );
  INVD1BWP30P140LVT U8731 ( .I(i_cmd[73]), .ZN(n8527) );
  OR2D1BWP30P140LVT U8732 ( .A1(i_cmd[33]), .A2(i_cmd[49]), .Z(n8225) );
  OR2D1BWP30P140LVT U8733 ( .A1(i_cmd[1]), .A2(i_cmd[17]), .Z(n8607) );
  ND2OPTIBD1BWP30P140LVT U8734 ( .A1(n10869), .A2(i_valid[29]), .ZN(n7769) );
  NR2D1BWP30P140LVT U8735 ( .A1(i_cmd[232]), .A2(i_cmd[248]), .ZN(n6267) );
  NR2D1BWP30P140LVT U8736 ( .A1(i_cmd[224]), .A2(i_cmd[240]), .ZN(n6268) );
  ND2OPTIBD1BWP30P140LVT U8737 ( .A1(n10869), .A2(i_valid[25]), .ZN(n7183) );
  OR2D1BWP30P140LVT U8738 ( .A1(i_cmd[208]), .A2(i_cmd[192]), .Z(n7182) );
  ND2OPTIBD1BWP30P140LVT U8739 ( .A1(n10869), .A2(i_valid[26]), .ZN(n7181) );
  OR2D1BWP30P140LVT U8740 ( .A1(i_cmd[160]), .A2(i_cmd[176]), .Z(n6692) );
  OR2D1BWP30P140LVT U8741 ( .A1(i_cmd[128]), .A2(i_cmd[144]), .Z(n10398) );
  NR2D1BWP30P140LVT U8742 ( .A1(i_cmd[96]), .A2(i_cmd[112]), .ZN(n6273) );
  OR2D1BWP30P140LVT U8743 ( .A1(i_cmd[64]), .A2(i_cmd[80]), .Z(n10393) );
  OR2D1BWP30P140LVT U8744 ( .A1(i_cmd[32]), .A2(i_cmd[48]), .Z(n10137) );
  OR2D1BWP30P140LVT U8745 ( .A1(i_cmd[0]), .A2(i_cmd[16]), .Z(n10375) );
  ND2D1BWP30P140LVT U8746 ( .A1(n11351), .A2(inner_first_stage_data_reg[162]), 
        .ZN(n11194) );
  ND2D1BWP30P140LVT U8747 ( .A1(n11344), .A2(inner_first_stage_data_reg[36]), 
        .ZN(n11204) );
  ND2D1BWP30P140LVT U8748 ( .A1(n11351), .A2(inner_first_stage_data_reg[175]), 
        .ZN(n11259) );
  ND2D1BWP30P140LVT U8749 ( .A1(n11351), .A2(inner_first_stage_data_reg[176]), 
        .ZN(n11264) );
  ND2D1BWP30P140LVT U8750 ( .A1(n11351), .A2(inner_first_stage_data_reg[184]), 
        .ZN(n11304) );
  ND2D1BWP30P140LVT U8751 ( .A1(n11351), .A2(inner_first_stage_data_reg[190]), 
        .ZN(n11334) );
  AN3D1BWP30P140LVT U8752 ( .A1(inner_first_stage_valid_reg[7]), .A2(n8588), 
        .A3(n8587), .Z(n11343) );
  AN3D1BWP30P140LVT U8753 ( .A1(inner_first_stage_valid_reg[2]), .A2(n8580), 
        .A3(n8584), .Z(n11339) );
  AN3D1BWP30P140LVT U8754 ( .A1(n8579), .A2(inner_first_stage_valid_reg[4]), 
        .A3(n8588), .Z(n11340) );
  AN4D1BWP30P140LVT U8755 ( .A1(n10863), .A2(n12302), .A3(
        inner_first_stage_valid_reg[12]), .A4(n10862), .Z(n11476) );
  AN3D1BWP30P140LVT U8756 ( .A1(n10887), .A2(inner_first_stage_valid_reg[21]), 
        .A3(n10886), .Z(n11615) );
  NR3D0P7BWP30P140LVT U8757 ( .A1(inner_first_stage_valid_reg[38]), .A2(n12303), .A3(n10868), .ZN(n11888) );
  NR3D0P7BWP30P140LVT U8758 ( .A1(inner_first_stage_valid_reg[39]), .A2(n10870), .A3(n10868), .ZN(n11889) );
  AN3D1BWP30P140LVT U8759 ( .A1(inner_first_stage_valid_reg[44]), .A2(n10901), 
        .A3(n10900), .Z(n12021) );
  AN4D1BWP30P140LVT U8760 ( .A1(n7374), .A2(n12302), .A3(
        inner_first_stage_valid_reg[52]), .A4(n7373), .Z(n12156) );
  NR3D0P7BWP30P140LVT U8761 ( .A1(inner_first_stage_valid_reg[62]), .A2(n8826), 
        .A3(n8827), .ZN(n12297) );
  AN3D1BWP30P140LVT U8762 ( .A1(inner_first_stage_valid_reg[60]), .A2(n8830), 
        .A3(n8824), .Z(n12295) );
  NR4D0BWP30P140LVT U8763 ( .A1(i_cmd[255]), .A2(n7532), .A3(n7769), .A4(n7530), .ZN(n8256) );
  NR2D1BWP30P140LVT U8764 ( .A1(n7767), .A2(n10912), .ZN(n8258) );
  ND2D1BWP30P140LVT U8765 ( .A1(n7531), .A2(n7530), .ZN(n10914) );
  ND2D1BWP30P140LVT U8766 ( .A1(i_cmd[231]), .A2(n10910), .ZN(n10912) );
  NR2D1BWP30P140LVT U8767 ( .A1(n7178), .A2(n10921), .ZN(n7335) );
  NR4D0BWP30P140LVT U8768 ( .A1(i_cmd[223]), .A2(n10919), .A3(n7183), .A4(
        n6990), .ZN(n7336) );
  INVD1BWP30P140LVT U8769 ( .I(i_cmd[223]), .ZN(n10918) );
  INVD1BWP30P140LVT U8770 ( .I(i_cmd[207]), .ZN(n10919) );
  ND2D1BWP30P140LVT U8771 ( .A1(i_cmd[199]), .A2(n10915), .ZN(n10921) );
  ND2D1BWP30P140LVT U8772 ( .A1(n10919), .A2(n10918), .ZN(n10916) );
  NR2D1BWP30P140LVT U8773 ( .A1(n6689), .A2(n6320), .ZN(n6878) );
  INVD1BWP30P140LVT U8774 ( .I(i_cmd[191]), .ZN(n6324) );
  INVD1BWP30P140LVT U8775 ( .I(i_cmd[175]), .ZN(n6322) );
  ND2D1BWP30P140LVT U8776 ( .A1(n6322), .A2(n6324), .ZN(n6321) );
  NR2D1BWP30P140LVT U8777 ( .A1(n10691), .A2(n10924), .ZN(n10852) );
  ND2D1BWP30P140LVT U8778 ( .A1(n10697), .A2(n10693), .ZN(n10926) );
  ND2D1BWP30P140LVT U8779 ( .A1(i_cmd[135]), .A2(n10922), .ZN(n10924) );
  NR2D1BWP30P140LVT U8780 ( .A1(n8445), .A2(n8377), .ZN(n10386) );
  NR2D1BWP30P140LVT U8781 ( .A1(n8443), .A2(n8375), .ZN(n10388) );
  NR2D1BWP30P140LVT U8782 ( .A1(n8447), .A2(n8376), .ZN(n10385) );
  NR2D1BWP30P140LVT U8783 ( .A1(n8441), .A2(n8374), .ZN(n10387) );
  INVD1BWP30P140LVT U8784 ( .I(i_cmd[95]), .ZN(n10930) );
  INVD1BWP30P140LVT U8785 ( .I(i_cmd[79]), .ZN(n10931) );
  ND2D1BWP30P140LVT U8786 ( .A1(i_cmd[71]), .A2(n10927), .ZN(n10933) );
  ND2D1BWP30P140LVT U8787 ( .A1(n10931), .A2(n10930), .ZN(n10928) );
  NR2D1BWP30P140LVT U8788 ( .A1(n10663), .A2(n10662), .ZN(n10830) );
  INVD1BWP30P140LVT U8789 ( .I(i_cmd[63]), .ZN(n10669) );
  INVD1BWP30P140LVT U8790 ( .I(i_cmd[47]), .ZN(n10665) );
  ND2D1BWP30P140LVT U8791 ( .A1(n10665), .A2(n10669), .ZN(n10666) );
  NR2D1BWP30P140LVT U8792 ( .A1(n10629), .A2(n10936), .ZN(n10812) );
  ND2D1BWP30P140LVT U8793 ( .A1(n10635), .A2(n10631), .ZN(n10938) );
  NR2D1BWP30P140LVT U8794 ( .A1(n7767), .A2(n10941), .ZN(n8342) );
  NR2D1BWP30P140LVT U8795 ( .A1(n7179), .A2(n7079), .ZN(n7363) );
  NR2D1BWP30P140LVT U8796 ( .A1(n7178), .A2(n7076), .ZN(n7365) );
  NR2D1BWP30P140LVT U8797 ( .A1(n7181), .A2(n7078), .ZN(n7364) );
  NR2D1BWP30P140LVT U8798 ( .A1(n7183), .A2(n7077), .ZN(n7366) );
  NR2D1BWP30P140LVT U8799 ( .A1(n6689), .A2(n10946), .ZN(n6924) );
  ND2D1BWP30P140LVT U8800 ( .A1(i_cmd[166]), .A2(n10944), .ZN(n10946) );
  INVD1BWP30P140LVT U8801 ( .I(i_cmd[158]), .ZN(n10952) );
  INVD1BWP30P140LVT U8802 ( .I(i_cmd[142]), .ZN(n10953) );
  ND2D1BWP30P140LVT U8803 ( .A1(i_cmd[134]), .A2(n10949), .ZN(n10955) );
  ND2D1BWP30P140LVT U8804 ( .A1(n10953), .A2(n10952), .ZN(n10950) );
  NR2D1BWP30P140LVT U8805 ( .A1(n8443), .A2(n8420), .ZN(n10408) );
  NR2D1BWP30P140LVT U8806 ( .A1(n8445), .A2(n8421), .ZN(n10405) );
  NR2D1BWP30P140LVT U8807 ( .A1(n8447), .A2(n8419), .ZN(n10406) );
  NR2D1BWP30P140LVT U8808 ( .A1(n8441), .A2(n8418), .ZN(n10407) );
  INVD1BWP30P140LVT U8809 ( .I(i_cmd[94]), .ZN(n10959) );
  INVD1BWP30P140LVT U8810 ( .I(i_cmd[78]), .ZN(n10960) );
  ND2D1BWP30P140LVT U8811 ( .A1(i_cmd[70]), .A2(n10956), .ZN(n10962) );
  ND2D1BWP30P140LVT U8812 ( .A1(n10960), .A2(n10959), .ZN(n10957) );
  INVD1BWP30P140LVT U8813 ( .I(i_cmd[62]), .ZN(n8319) );
  INVD1BWP30P140LVT U8814 ( .I(i_cmd[46]), .ZN(n8321) );
  ND2D1BWP30P140LVT U8815 ( .A1(n8321), .A2(n8319), .ZN(n8318) );
  ND2D1BWP30P140LVT U8816 ( .A1(n8488), .A2(n8486), .ZN(n10967) );
  ND2D1BWP30P140LVT U8817 ( .A1(i_cmd[6]), .A2(n10963), .ZN(n10965) );
  NR2D1BWP30P140LVT U8818 ( .A1(n7767), .A2(n10970), .ZN(n8233) );
  ND2D1BWP30P140LVT U8819 ( .A1(i_cmd[229]), .A2(n10968), .ZN(n10970) );
  NR4D0BWP30P140LVT U8820 ( .A1(i_cmd[221]), .A2(n7183), .A3(n6995), .A4(n6996), .ZN(n7326) );
  NR2D1BWP30P140LVT U8821 ( .A1(n7178), .A2(n10975), .ZN(n7325) );
  ND2D1BWP30P140LVT U8822 ( .A1(i_cmd[197]), .A2(n10973), .ZN(n10975) );
  ND2D1BWP30P140LVT U8823 ( .A1(n6997), .A2(n6995), .ZN(n10977) );
  NR2D1BWP30P140LVT U8824 ( .A1(n6689), .A2(n10984), .ZN(n6884) );
  INVD1BWP30P140LVT U8825 ( .I(i_cmd[189]), .ZN(n10981) );
  INVD1BWP30P140LVT U8826 ( .I(i_cmd[173]), .ZN(n10982) );
  ND2D1BWP30P140LVT U8827 ( .A1(i_cmd[165]), .A2(n10978), .ZN(n10984) );
  ND2D1BWP30P140LVT U8828 ( .A1(n10982), .A2(n10981), .ZN(n10979) );
  ND2D1BWP30P140LVT U8829 ( .A1(i_cmd[133]), .A2(n10985), .ZN(n10987) );
  INVD1BWP30P140LVT U8830 ( .I(i_cmd[109]), .ZN(n10993) );
  INVD1BWP30P140LVT U8831 ( .I(i_cmd[125]), .ZN(n10994) );
  ND2D1BWP30P140LVT U8832 ( .A1(i_cmd[101]), .A2(n10990), .ZN(n10996) );
  ND2D1BWP30P140LVT U8833 ( .A1(n10994), .A2(n10993), .ZN(n10991) );
  NR2D1BWP30P140LVT U8834 ( .A1(n10394), .A2(n11003), .ZN(n9846) );
  INVD1BWP30P140LVT U8835 ( .I(i_cmd[77]), .ZN(n11000) );
  INVD1BWP30P140LVT U8836 ( .I(i_cmd[93]), .ZN(n11001) );
  ND2D1BWP30P140LVT U8837 ( .A1(i_cmd[69]), .A2(n10997), .ZN(n11003) );
  ND2D1BWP30P140LVT U8838 ( .A1(n11001), .A2(n11000), .ZN(n10998) );
  ND2D1BWP30P140LVT U8839 ( .A1(n8367), .A2(n8365), .ZN(n11008) );
  ND2D1BWP30P140LVT U8840 ( .A1(i_cmd[37]), .A2(n11004), .ZN(n11006) );
  ND2D1BWP30P140LVT U8841 ( .A1(n8493), .A2(n8491), .ZN(n11013) );
  ND2D1BWP30P140LVT U8842 ( .A1(i_cmd[5]), .A2(n11009), .ZN(n11011) );
  NR2D1BWP30P140LVT U8843 ( .A1(n7765), .A2(n7764), .ZN(n9662) );
  NR2D1BWP30P140LVT U8844 ( .A1(n7769), .A2(n7768), .ZN(n9660) );
  NR2D1BWP30P140LVT U8845 ( .A1(n7771), .A2(n7770), .ZN(n9663) );
  NR2D1BWP30P140LVT U8846 ( .A1(n7767), .A2(n7766), .ZN(n9661) );
  NR2D1BWP30P140LVT U8847 ( .A1(n7178), .A2(n11016), .ZN(n6758) );
  NR2D1BWP30P140LVT U8848 ( .A1(n6689), .A2(n11025), .ZN(n6398) );
  INVD1BWP30P140LVT U8849 ( .I(i_cmd[172]), .ZN(n11022) );
  INVD1BWP30P140LVT U8850 ( .I(i_cmd[188]), .ZN(n11023) );
  ND2D1BWP30P140LVT U8851 ( .A1(i_cmd[164]), .A2(n11019), .ZN(n11025) );
  ND2D1BWP30P140LVT U8852 ( .A1(n11023), .A2(n11022), .ZN(n11020) );
  NR2D1BWP30P140LVT U8853 ( .A1(n10691), .A2(n11032), .ZN(n10182) );
  INVD1BWP30P140LVT U8854 ( .I(i_cmd[156]), .ZN(n11029) );
  INVD1BWP30P140LVT U8855 ( .I(i_cmd[140]), .ZN(n11030) );
  ND2D1BWP30P140LVT U8856 ( .A1(i_cmd[132]), .A2(n11026), .ZN(n11032) );
  ND2D1BWP30P140LVT U8857 ( .A1(n11030), .A2(n11029), .ZN(n11027) );
  NR2D1BWP30P140LVT U8858 ( .A1(n8445), .A2(n8444), .ZN(n10427) );
  NR2D1BWP30P140LVT U8859 ( .A1(n8447), .A2(n8446), .ZN(n10428) );
  NR2D1BWP30P140LVT U8860 ( .A1(n8443), .A2(n8442), .ZN(n10430) );
  NR2D1BWP30P140LVT U8861 ( .A1(n8441), .A2(n8440), .ZN(n10429) );
  NR2D1BWP30P140LVT U8862 ( .A1(n10394), .A2(n11039), .ZN(n10052) );
  INVD1BWP30P140LVT U8863 ( .I(i_cmd[76]), .ZN(n11036) );
  INVD1BWP30P140LVT U8864 ( .I(i_cmd[92]), .ZN(n11037) );
  ND2D1BWP30P140LVT U8865 ( .A1(i_cmd[68]), .A2(n11033), .ZN(n11039) );
  ND2D1BWP30P140LVT U8866 ( .A1(n11037), .A2(n11036), .ZN(n11034) );
  NR2D1BWP30P140LVT U8867 ( .A1(n10663), .A2(n11042), .ZN(n10224) );
  ND2D1BWP30P140LVT U8868 ( .A1(n8244), .A2(n8242), .ZN(n11044) );
  NR2D1BWP30P140LVT U8869 ( .A1(n10629), .A2(n11051), .ZN(n10096) );
  INVD1BWP30P140LVT U8870 ( .I(i_cmd[12]), .ZN(n11048) );
  INVD1BWP30P140LVT U8871 ( .I(i_cmd[28]), .ZN(n11049) );
  ND2D1BWP30P140LVT U8872 ( .A1(i_cmd[4]), .A2(n11045), .ZN(n11051) );
  ND2D1BWP30P140LVT U8873 ( .A1(n11049), .A2(n11048), .ZN(n11046) );
  NR4D0BWP30P140LVT U8874 ( .A1(i_cmd[251]), .A2(n11056), .A3(n7769), .A4(
        n7484), .ZN(n8208) );
  NR2D1BWP30P140LVT U8875 ( .A1(n7767), .A2(n11059), .ZN(n8206) );
  INVD1BWP30P140LVT U8876 ( .I(i_cmd[251]), .ZN(n11055) );
  INVD1BWP30P140LVT U8877 ( .I(i_cmd[235]), .ZN(n11056) );
  ND2D1BWP30P140LVT U8878 ( .A1(i_cmd[227]), .A2(n11052), .ZN(n11059) );
  ND2D1BWP30P140LVT U8879 ( .A1(n11056), .A2(n11055), .ZN(n11053) );
  NR4D0BWP30P140LVT U8880 ( .A1(i_cmd[219]), .A2(n7183), .A3(n6419), .A4(n6418), .ZN(n6721) );
  NR2D1BWP30P140LVT U8881 ( .A1(n7178), .A2(n11062), .ZN(n6720) );
  ND2D1BWP30P140LVT U8882 ( .A1(i_cmd[195]), .A2(n11060), .ZN(n11062) );
  ND2D1BWP30P140LVT U8883 ( .A1(n6417), .A2(n6419), .ZN(n11064) );
  NR2D1BWP30P140LVT U8884 ( .A1(n6689), .A2(n11067), .ZN(n6910) );
  ND2D1BWP30P140LVT U8885 ( .A1(i_cmd[163]), .A2(n11065), .ZN(n11067) );
  NR2D1BWP30P140LVT U8886 ( .A1(n10691), .A2(n11072), .ZN(n9934) );
  ND2D1BWP30P140LVT U8887 ( .A1(i_cmd[131]), .A2(n11070), .ZN(n11072) );
  INVD1BWP30P140LVT U8888 ( .I(i_cmd[123]), .ZN(n11078) );
  INVD1BWP30P140LVT U8889 ( .I(i_cmd[107]), .ZN(n11079) );
  ND2D1BWP30P140LVT U8890 ( .A1(i_cmd[99]), .A2(n11075), .ZN(n11081) );
  ND2D1BWP30P140LVT U8891 ( .A1(n11079), .A2(n11078), .ZN(n11076) );
  NR2D1BWP30P140LVT U8892 ( .A1(n10394), .A2(n11088), .ZN(n9756) );
  INVD1BWP30P140LVT U8893 ( .I(i_cmd[75]), .ZN(n11085) );
  INVD1BWP30P140LVT U8894 ( .I(i_cmd[91]), .ZN(n11086) );
  ND2D1BWP30P140LVT U8895 ( .A1(i_cmd[67]), .A2(n11082), .ZN(n11088) );
  ND2D1BWP30P140LVT U8896 ( .A1(n11086), .A2(n11085), .ZN(n11083) );
  NR2D1BWP30P140LVT U8897 ( .A1(n10663), .A2(n11095), .ZN(n9522) );
  INVD1BWP30P140LVT U8898 ( .I(i_cmd[43]), .ZN(n11092) );
  INVD1BWP30P140LVT U8899 ( .I(i_cmd[59]), .ZN(n11093) );
  ND2D1BWP30P140LVT U8900 ( .A1(i_cmd[35]), .A2(n11089), .ZN(n11095) );
  ND2D1BWP30P140LVT U8901 ( .A1(n11093), .A2(n11092), .ZN(n11090) );
  NR2D1BWP30P140LVT U8902 ( .A1(n10629), .A2(n8541), .ZN(n10088) );
  INVD1BWP30P140LVT U8903 ( .I(i_cmd[27]), .ZN(n8539) );
  INVD1BWP30P140LVT U8904 ( .I(i_cmd[11]), .ZN(n8537) );
  ND2D1BWP30P140LVT U8905 ( .A1(n8537), .A2(n8539), .ZN(n8540) );
  NR4D0BWP30P140LVT U8906 ( .A1(i_cmd[250]), .A2(n7555), .A3(n7769), .A4(n7554), .ZN(n8351) );
  NR2D1BWP30P140LVT U8907 ( .A1(n7767), .A2(n7553), .ZN(n8354) );
  INVD1BWP30P140LVT U8908 ( .I(i_cmd[250]), .ZN(n7552) );
  INVD1BWP30P140LVT U8909 ( .I(i_cmd[234]), .ZN(n7555) );
  ND2D1BWP30P140LVT U8910 ( .A1(n7555), .A2(n7552), .ZN(n7551) );
  NR2D1BWP30P140LVT U8911 ( .A1(n7178), .A2(n11098), .ZN(n7303) );
  NR2D1BWP30P140LVT U8912 ( .A1(n6693), .A2(n6411), .ZN(n6620) );
  NR2D1BWP30P140LVT U8913 ( .A1(n6691), .A2(n6409), .ZN(n6619) );
  NR2D1BWP30P140LVT U8914 ( .A1(n6690), .A2(n6410), .ZN(n6618) );
  INVD1BWP30P140LVT U8915 ( .I(i_cmd[154]), .ZN(n7832) );
  INVD1BWP30P140LVT U8916 ( .I(i_cmd[138]), .ZN(n7829) );
  ND2D1BWP30P140LVT U8917 ( .A1(n7829), .A2(n7832), .ZN(n7833) );
  ND2D1BWP30P140LVT U8918 ( .A1(i_cmd[130]), .A2(n6247), .ZN(n7830) );
  ND2D1BWP30P140LVT U8919 ( .A1(i_cmd[98]), .A2(n11101), .ZN(n11103) );
  INVD1BWP30P140LVT U8920 ( .I(i_cmd[90]), .ZN(n8568) );
  INVD1BWP30P140LVT U8921 ( .I(i_cmd[74]), .ZN(n8566) );
  ND2D1BWP30P140LVT U8922 ( .A1(n8566), .A2(n8568), .ZN(n8569) );
  INVD1BWP30P140LVT U8923 ( .I(i_cmd[58]), .ZN(n11109) );
  INVD1BWP30P140LVT U8924 ( .I(i_cmd[42]), .ZN(n11110) );
  ND2D1BWP30P140LVT U8925 ( .A1(i_cmd[34]), .A2(n11106), .ZN(n11112) );
  ND2D1BWP30P140LVT U8926 ( .A1(n11110), .A2(n11109), .ZN(n11107) );
  INVD1BWP30P140LVT U8927 ( .I(i_cmd[26]), .ZN(n8502) );
  INVD1BWP30P140LVT U8928 ( .I(i_cmd[10]), .ZN(n8504) );
  ND2D1BWP30P140LVT U8929 ( .A1(n8504), .A2(n8502), .ZN(n8501) );
  NR4D0BWP30P140LVT U8930 ( .A1(i_cmd[249]), .A2(n11117), .A3(n7769), .A4(
        n7583), .ZN(n8720) );
  NR2D1BWP30P140LVT U8931 ( .A1(n7767), .A2(n11119), .ZN(n8722) );
  INVD1BWP30P140LVT U8932 ( .I(i_cmd[249]), .ZN(n11116) );
  INVD1BWP30P140LVT U8933 ( .I(i_cmd[233]), .ZN(n11117) );
  ND2D1BWP30P140LVT U8934 ( .A1(i_cmd[225]), .A2(n11113), .ZN(n11119) );
  ND2D1BWP30P140LVT U8935 ( .A1(n11117), .A2(n11116), .ZN(n11114) );
  NR2D1BWP30P140LVT U8936 ( .A1(n7178), .A2(n11122), .ZN(n7353) );
  ND2D1BWP30P140LVT U8937 ( .A1(i_cmd[193]), .A2(n11120), .ZN(n11122) );
  NR2D1BWP30P140LVT U8938 ( .A1(n6691), .A2(n6550), .ZN(n6941) );
  NR2D1BWP30P140LVT U8939 ( .A1(n6690), .A2(n6551), .ZN(n6940) );
  NR2D1BWP30P140LVT U8940 ( .A1(n6693), .A2(n6549), .ZN(n6943) );
  NR2D1BWP30P140LVT U8941 ( .A1(n6689), .A2(n6548), .ZN(n6942) );
  INVD1BWP30P140LVT U8942 ( .I(i_cmd[153]), .ZN(n11128) );
  INVD1BWP30P140LVT U8943 ( .I(i_cmd[137]), .ZN(n11129) );
  ND2D1BWP30P140LVT U8944 ( .A1(i_cmd[129]), .A2(n11125), .ZN(n11131) );
  ND2D1BWP30P140LVT U8945 ( .A1(n11129), .A2(n11128), .ZN(n11126) );
  NR2D1BWP30P140LVT U8946 ( .A1(n8443), .A2(n7935), .ZN(n8124) );
  NR2D1BWP30P140LVT U8947 ( .A1(n8445), .A2(n7937), .ZN(n8125) );
  NR2D1BWP30P140LVT U8948 ( .A1(n8447), .A2(n7936), .ZN(n8123) );
  NR2D1BWP30P140LVT U8949 ( .A1(n8441), .A2(n7938), .ZN(n8122) );
  ND2D1BWP30P140LVT U8950 ( .A1(n8527), .A2(n8525), .ZN(n11136) );
  INVD1BWP30P140LVT U8951 ( .I(i_cmd[57]), .ZN(n11140) );
  INVD1BWP30P140LVT U8952 ( .I(i_cmd[41]), .ZN(n11141) );
  ND2D1BWP30P140LVT U8953 ( .A1(i_cmd[33]), .A2(n11137), .ZN(n11143) );
  ND2D1BWP30P140LVT U8954 ( .A1(n11141), .A2(n11140), .ZN(n11138) );
  INVD1BWP30P140LVT U8955 ( .I(i_cmd[9]), .ZN(n11147) );
  INVD1BWP30P140LVT U8956 ( .I(i_cmd[25]), .ZN(n11148) );
  ND2D1BWP30P140LVT U8957 ( .A1(i_cmd[1]), .A2(n11144), .ZN(n11150) );
  ND2D1BWP30P140LVT U8958 ( .A1(n11148), .A2(n11147), .ZN(n11145) );
  NR2D1BWP30P140LVT U8959 ( .A1(n7765), .A2(n7732), .ZN(n9544) );
  NR2D1BWP30P140LVT U8960 ( .A1(n7771), .A2(n7734), .ZN(n9543) );
  NR2D1BWP30P140LVT U8961 ( .A1(n7769), .A2(n7735), .ZN(n9545) );
  NR2D1BWP30P140LVT U8962 ( .A1(n7178), .A2(n11153), .ZN(n7424) );
  NR4D0BWP30P140LVT U8963 ( .A1(i_cmd[216]), .A2(n7184), .A3(n7183), .A4(n7182), .ZN(n7423) );
  ND2D1BWP30P140LVT U8964 ( .A1(i_cmd[192]), .A2(n11151), .ZN(n11153) );
  ND2D1BWP30P140LVT U8965 ( .A1(n7184), .A2(n7180), .ZN(n11155) );
  NR2D1BWP30P140LVT U8966 ( .A1(n6689), .A2(n11158), .ZN(n6986) );
  ND2D1BWP30P140LVT U8967 ( .A1(i_cmd[160]), .A2(n11156), .ZN(n11158) );
  INVD1BWP30P140LVT U8968 ( .I(i_cmd[152]), .ZN(n11164) );
  INVD1BWP30P140LVT U8969 ( .I(i_cmd[136]), .ZN(n11165) );
  ND2D1BWP30P140LVT U8970 ( .A1(i_cmd[128]), .A2(n11161), .ZN(n11167) );
  ND2D1BWP30P140LVT U8971 ( .A1(n11165), .A2(n11164), .ZN(n11162) );
  NR2D1BWP30P140LVT U8972 ( .A1(n8445), .A2(n7428), .ZN(n8041) );
  INVD1BWP30P140LVT U8973 ( .I(i_cmd[88]), .ZN(n11171) );
  INVD1BWP30P140LVT U8974 ( .I(i_cmd[72]), .ZN(n11172) );
  ND2D1BWP30P140LVT U8975 ( .A1(i_cmd[64]), .A2(n11168), .ZN(n11175) );
  ND2D1BWP30P140LVT U8976 ( .A1(n11172), .A2(n11171), .ZN(n11169) );
  INVD1BWP30P140LVT U8977 ( .I(i_cmd[56]), .ZN(n11179) );
  INVD1BWP30P140LVT U8978 ( .I(i_cmd[40]), .ZN(n11180) );
  ND2D1BWP30P140LVT U8979 ( .A1(i_cmd[32]), .A2(n11176), .ZN(n11183) );
  ND2D1BWP30P140LVT U8980 ( .A1(n11180), .A2(n11179), .ZN(n11177) );
  INVD1BWP30P140LVT U8981 ( .I(i_cmd[24]), .ZN(n10373) );
  INVD1BWP30P140LVT U8982 ( .I(i_cmd[8]), .ZN(n10376) );
  ND2D1BWP30P140LVT U8983 ( .A1(n10376), .A2(n10373), .ZN(n10372) );
  ND2D1BWP30P140LVT U8984 ( .A1(i_cmd[0]), .A2(n6250), .ZN(n10374) );
  ND2D1BWP30P140LVT U8985 ( .A1(n11344), .A2(inner_first_stage_data_reg[32]), 
        .ZN(n11184) );
  ND2D1BWP30P140LVT U8986 ( .A1(n11351), .A2(inner_first_stage_data_reg[161]), 
        .ZN(n11189) );
  ND2D1BWP30P140LVT U8987 ( .A1(n11345), .A2(inner_first_stage_data_reg[5]), 
        .ZN(n11209) );
  ND2D1BWP30P140LVT U8988 ( .A1(n11351), .A2(inner_first_stage_data_reg[166]), 
        .ZN(n11214) );
  ND2D1BWP30P140LVT U8989 ( .A1(n11351), .A2(inner_first_stage_data_reg[169]), 
        .ZN(n11229) );
  ND2D1BWP30P140LVT U8990 ( .A1(n11351), .A2(inner_first_stage_data_reg[170]), 
        .ZN(n11234) );
  ND2D1BWP30P140LVT U8991 ( .A1(n11345), .A2(inner_first_stage_data_reg[12]), 
        .ZN(n11244) );
  ND2D1BWP30P140LVT U8992 ( .A1(n11351), .A2(inner_first_stage_data_reg[177]), 
        .ZN(n11269) );
  ND2D1BWP30P140LVT U8993 ( .A1(n11351), .A2(inner_first_stage_data_reg[180]), 
        .ZN(n11284) );
  ND2D1BWP30P140LVT U8994 ( .A1(n11344), .A2(inner_first_stage_data_reg[53]), 
        .ZN(n11289) );
  ND2D1BWP30P140LVT U8995 ( .A1(n11344), .A2(inner_first_stage_data_reg[54]), 
        .ZN(n11294) );
  ND2D1BWP30P140LVT U8996 ( .A1(n11344), .A2(inner_first_stage_data_reg[55]), 
        .ZN(n11299) );
  ND2D1BWP30P140LVT U8997 ( .A1(n11344), .A2(inner_first_stage_data_reg[57]), 
        .ZN(n11309) );
  ND2D1BWP30P140LVT U8998 ( .A1(n11351), .A2(inner_first_stage_data_reg[186]), 
        .ZN(n11314) );
  ND2D1BWP30P140LVT U8999 ( .A1(n11344), .A2(inner_first_stage_data_reg[60]), 
        .ZN(n11324) );
  ND2D1BWP30P140LVT U9000 ( .A1(n11351), .A2(inner_first_stage_data_reg[189]), 
        .ZN(n11329) );
  ND2D1BWP30P140LVT U9001 ( .A1(n11345), .A2(inner_first_stage_data_reg[31]), 
        .ZN(n11346) );
  ND2D1BWP30P140LVT U9002 ( .A1(n8590), .A2(n8589), .ZN(N2228) );
  ND2D1BWP30P140LVT U9003 ( .A1(n10867), .A2(n10866), .ZN(N3078) );
  ND2D1BWP30P140LVT U9004 ( .A1(n10895), .A2(n10894), .ZN(N4952) );
  ND2D1BWP30P140LVT U9005 ( .A1(n7463), .A2(n7462), .ZN(N5802) );
  ND2D1BWP30P140LVT U9006 ( .A1(n10881), .A2(n10880), .ZN(N7676) );
  ND2D1BWP30P140LVT U9007 ( .A1(n10909), .A2(n10908), .ZN(N8526) );
  ND2D1BWP30P140LVT U9008 ( .A1(n7381), .A2(n7380), .ZN(N10400) );
  ND2D1BWP30P140LVT U9009 ( .A1(n8836), .A2(n8835), .ZN(N11250) );
  ND2D1BWP30P140LVT U9010 ( .A1(n10400), .A2(n10399), .ZN(N1423) );
  ND2D1BWP30P140LVT U9011 ( .A1(n10603), .A2(n10602), .ZN(N1424) );
  ND2D1BWP30P140LVT U9012 ( .A1(n10466), .A2(n10465), .ZN(N1425) );
  ND2D1BWP30P140LVT U9013 ( .A1(n10597), .A2(n10596), .ZN(N1426) );
  ND2D1BWP30P140LVT U9014 ( .A1(n10621), .A2(n10620), .ZN(N1427) );
  ND2D1BWP30P140LVT U9015 ( .A1(n10490), .A2(n10489), .ZN(N1428) );
  ND2D1BWP30P140LVT U9016 ( .A1(n10599), .A2(n10598), .ZN(N1429) );
  ND2D1BWP30P140LVT U9017 ( .A1(n10605), .A2(n10604), .ZN(N1430) );
  ND2D1BWP30P140LVT U9018 ( .A1(n10480), .A2(n10479), .ZN(N1431) );
  ND2D1BWP30P140LVT U9019 ( .A1(n10488), .A2(n10487), .ZN(N1432) );
  ND2D1BWP30P140LVT U9020 ( .A1(n10468), .A2(n10467), .ZN(N1433) );
  ND2D1BWP30P140LVT U9021 ( .A1(n10482), .A2(n10481), .ZN(N1434) );
  ND2D1BWP30P140LVT U9022 ( .A1(n10623), .A2(n10622), .ZN(N1435) );
  ND2D1BWP30P140LVT U9023 ( .A1(n10476), .A2(n10475), .ZN(N1436) );
  ND2D1BWP30P140LVT U9024 ( .A1(n10613), .A2(n10612), .ZN(N1437) );
  ND2D1BWP30P140LVT U9025 ( .A1(n10601), .A2(n10600), .ZN(N1438) );
  ND2D1BWP30P140LVT U9026 ( .A1(n10607), .A2(n10606), .ZN(N1439) );
  ND2D1BWP30P140LVT U9027 ( .A1(n10617), .A2(n10616), .ZN(N1440) );
  ND2D1BWP30P140LVT U9028 ( .A1(n10628), .A2(n10627), .ZN(N1441) );
  ND2D1BWP30P140LVT U9029 ( .A1(n10474), .A2(n10473), .ZN(N1442) );
  ND2D1BWP30P140LVT U9030 ( .A1(n10464), .A2(n10463), .ZN(N1443) );
  ND2D1BWP30P140LVT U9031 ( .A1(n10470), .A2(n10469), .ZN(N1444) );
  ND2D1BWP30P140LVT U9032 ( .A1(n10472), .A2(n10471), .ZN(N1445) );
  ND2D1BWP30P140LVT U9033 ( .A1(n10609), .A2(n10608), .ZN(N1446) );
  ND2D1BWP30P140LVT U9034 ( .A1(n10593), .A2(n10592), .ZN(N1447) );
  ND2D1BWP30P140LVT U9035 ( .A1(n10611), .A2(n10610), .ZN(N1448) );
  ND2D1BWP30P140LVT U9036 ( .A1(n10484), .A2(n10483), .ZN(N1449) );
  ND2D1BWP30P140LVT U9037 ( .A1(n10615), .A2(n10614), .ZN(N1450) );
  ND2D1BWP30P140LVT U9038 ( .A1(n10595), .A2(n10594), .ZN(N1451) );
  ND2D1BWP30P140LVT U9039 ( .A1(n10619), .A2(n10618), .ZN(N1452) );
  ND2D1BWP30P140LVT U9040 ( .A1(n10486), .A2(n10485), .ZN(N1453) );
  ND2D1BWP30P140LVT U9041 ( .A1(n10478), .A2(n10477), .ZN(N1454) );
  ND2D1BWP30P140LVT U9042 ( .A1(n10506), .A2(n10505), .ZN(N983) );
  ND2D1BWP30P140LVT U9043 ( .A1(n10492), .A2(n10491), .ZN(N984) );
  ND2D1BWP30P140LVT U9044 ( .A1(n10498), .A2(n10497), .ZN(N985) );
  ND2D1BWP30P140LVT U9045 ( .A1(n10548), .A2(n10547), .ZN(N986) );
  ND2D1BWP30P140LVT U9046 ( .A1(n10508), .A2(n10507), .ZN(N987) );
  ND2D1BWP30P140LVT U9047 ( .A1(n10542), .A2(n10541), .ZN(N988) );
  ND2D1BWP30P140LVT U9048 ( .A1(n10544), .A2(n10543), .ZN(N989) );
  ND2D1BWP30P140LVT U9049 ( .A1(n10518), .A2(n10517), .ZN(N990) );
  ND2D1BWP30P140LVT U9050 ( .A1(n10538), .A2(n10537), .ZN(N991) );
  ND2D1BWP30P140LVT U9051 ( .A1(n10546), .A2(n10545), .ZN(N992) );
  ND2D1BWP30P140LVT U9052 ( .A1(n10504), .A2(n10503), .ZN(N993) );
  ND2D1BWP30P140LVT U9053 ( .A1(n10534), .A2(n10533), .ZN(N994) );
  ND2D1BWP30P140LVT U9054 ( .A1(n10524), .A2(n10523), .ZN(N995) );
  ND2D1BWP30P140LVT U9055 ( .A1(n10536), .A2(n10535), .ZN(N996) );
  ND2D1BWP30P140LVT U9056 ( .A1(n10516), .A2(n10515), .ZN(N997) );
  ND2D1BWP30P140LVT U9057 ( .A1(n10496), .A2(n10495), .ZN(N998) );
  ND2D1BWP30P140LVT U9058 ( .A1(n10520), .A2(n10519), .ZN(N999) );
  ND2D1BWP30P140LVT U9059 ( .A1(n10550), .A2(n10549), .ZN(N1000) );
  ND2D1BWP30P140LVT U9060 ( .A1(n10522), .A2(n10521), .ZN(N1001) );
  ND2D1BWP30P140LVT U9061 ( .A1(n10540), .A2(n10539), .ZN(N1002) );
  ND2D1BWP30P140LVT U9062 ( .A1(n10526), .A2(n10525), .ZN(N1003) );
  ND2D1BWP30P140LVT U9063 ( .A1(n10556), .A2(n10555), .ZN(N1004) );
  ND2D1BWP30P140LVT U9064 ( .A1(n10514), .A2(n10513), .ZN(N1005) );
  ND2D1BWP30P140LVT U9065 ( .A1(n10512), .A2(n10511), .ZN(N1006) );
  ND2D1BWP30P140LVT U9066 ( .A1(n10530), .A2(n10529), .ZN(N1007) );
  ND2D1BWP30P140LVT U9067 ( .A1(n10528), .A2(n10527), .ZN(N1008) );
  ND2D1BWP30P140LVT U9068 ( .A1(n10532), .A2(n10531), .ZN(N1009) );
  ND2D1BWP30P140LVT U9069 ( .A1(n10510), .A2(n10509), .ZN(N1010) );
  ND2D1BWP30P140LVT U9070 ( .A1(n10494), .A2(n10493), .ZN(N1011) );
  ND2D1BWP30P140LVT U9071 ( .A1(n10502), .A2(n10501), .ZN(N1012) );
  ND2D1BWP30P140LVT U9072 ( .A1(n10397), .A2(n10396), .ZN(N1013) );
  ND2D1BWP30P140LVT U9073 ( .A1(n10500), .A2(n10499), .ZN(N1014) );
  ND2D1BWP30P140LVT U9074 ( .A1(n10359), .A2(n10358), .ZN(N763) );
  ND2D1BWP30P140LVT U9075 ( .A1(n10362), .A2(n10361), .ZN(N764) );
  ND2D1BWP30P140LVT U9076 ( .A1(n10371), .A2(n10370), .ZN(N769) );
  ND2D1BWP30P140LVT U9077 ( .A1(n10307), .A2(n10306), .ZN(N777) );
  ND2D1BWP30P140LVT U9078 ( .A1(n10309), .A2(n10308), .ZN(N781) );
  ND2D1BWP30P140LVT U9079 ( .A1(n10364), .A2(n10363), .ZN(N782) );
  ND2D1BWP30P140LVT U9080 ( .A1(n10311), .A2(n10310), .ZN(N786) );
  ND2D1BWP30P140LVT U9081 ( .A1(n10305), .A2(n10304), .ZN(N787) );
  ND2D1BWP30P140LVT U9082 ( .A1(n10313), .A2(n10312), .ZN(N789) );
  ND2D1BWP30P140LVT U9083 ( .A1(n10366), .A2(n10365), .ZN(N791) );
  ND2D1BWP30P140LVT U9084 ( .A1(n10378), .A2(n10377), .ZN(N543) );
  ND2D1BWP30P140LVT U9085 ( .A1(n10570), .A2(n10569), .ZN(N544) );
  ND2D1BWP30P140LVT U9086 ( .A1(n10574), .A2(n10573), .ZN(N545) );
  ND2D1BWP30P140LVT U9087 ( .A1(n10560), .A2(n10559), .ZN(N546) );
  ND2D1BWP30P140LVT U9088 ( .A1(n10566), .A2(n10565), .ZN(N547) );
  ND2D1BWP30P140LVT U9089 ( .A1(n10562), .A2(n10561), .ZN(N548) );
  ND2D1BWP30P140LVT U9090 ( .A1(n10558), .A2(n10557), .ZN(N549) );
  ND2D1BWP30P140LVT U9091 ( .A1(n10448), .A2(n10447), .ZN(N550) );
  ND2D1BWP30P140LVT U9092 ( .A1(n10582), .A2(n10581), .ZN(N551) );
  ND2D1BWP30P140LVT U9093 ( .A1(n10450), .A2(n10449), .ZN(N552) );
  ND2D1BWP30P140LVT U9094 ( .A1(n10578), .A2(n10577), .ZN(N553) );
  ND2D1BWP30P140LVT U9095 ( .A1(n10434), .A2(n10433), .ZN(N554) );
  ND2D1BWP30P140LVT U9096 ( .A1(n10580), .A2(n10579), .ZN(N555) );
  ND2D1BWP30P140LVT U9097 ( .A1(n10438), .A2(n10437), .ZN(N556) );
  ND2D1BWP30P140LVT U9098 ( .A1(n10442), .A2(n10441), .ZN(N557) );
  ND2D1BWP30P140LVT U9099 ( .A1(n10568), .A2(n10567), .ZN(N558) );
  ND2D1BWP30P140LVT U9100 ( .A1(n10436), .A2(n10435), .ZN(N559) );
  ND2D1BWP30P140LVT U9101 ( .A1(n10444), .A2(n10443), .ZN(N560) );
  ND2D1BWP30P140LVT U9102 ( .A1(n10456), .A2(n10455), .ZN(N561) );
  ND2D1BWP30P140LVT U9103 ( .A1(n10458), .A2(n10457), .ZN(N562) );
  ND2D1BWP30P140LVT U9104 ( .A1(n10462), .A2(n10461), .ZN(N563) );
  ND2D1BWP30P140LVT U9105 ( .A1(n10584), .A2(n10583), .ZN(N564) );
  ND2D1BWP30P140LVT U9106 ( .A1(n10564), .A2(n10563), .ZN(N565) );
  ND2D1BWP30P140LVT U9107 ( .A1(n10452), .A2(n10451), .ZN(N566) );
  ND2D1BWP30P140LVT U9108 ( .A1(n10454), .A2(n10453), .ZN(N567) );
  ND2D1BWP30P140LVT U9109 ( .A1(n10572), .A2(n10571), .ZN(N568) );
  ND2D1BWP30P140LVT U9110 ( .A1(n10576), .A2(n10575), .ZN(N569) );
  ND2D1BWP30P140LVT U9111 ( .A1(n10586), .A2(n10585), .ZN(N570) );
  ND2D1BWP30P140LVT U9112 ( .A1(n10446), .A2(n10445), .ZN(N571) );
  ND2D1BWP30P140LVT U9113 ( .A1(n10460), .A2(n10459), .ZN(N572) );
  ND2D1BWP30P140LVT U9114 ( .A1(n10440), .A2(n10439), .ZN(N573) );
  ND2D1BWP30P140LVT U9115 ( .A1(n10591), .A2(n10590), .ZN(N574) );
  NR2D1BWP30P140LVT U9116 ( .A1(n8443), .A2(n7431), .ZN(n7434) );
  NR2D1BWP30P140LVT U9117 ( .A1(n8441), .A2(n7429), .ZN(n6212) );
  NR2D1BWP30P140LVT U9118 ( .A1(n10663), .A2(n11143), .ZN(n6213) );
  NR2D1BWP30P140LVT U9119 ( .A1(n8441), .A2(n10996), .ZN(n6214) );
  NR2D1BWP30P140LVT U9120 ( .A1(n8441), .A2(n11081), .ZN(n6215) );
  NR2D1BWP30P140LVT U9121 ( .A1(n10394), .A2(n11134), .ZN(n6216) );
  NR2D1BWP30P140LVT U9122 ( .A1(n10394), .A2(n10933), .ZN(n6217) );
  NR2D1BWP30P140LVT U9123 ( .A1(n10629), .A2(n8505), .ZN(n6218) );
  NR2D1BWP30P140LVT U9124 ( .A1(n10394), .A2(n8570), .ZN(n6219) );
  NR2D1BWP30P140LVT U9125 ( .A1(n10691), .A2(n11167), .ZN(n6220) );
  NR2D1BWP30P140LVT U9126 ( .A1(n10629), .A2(n10374), .ZN(n6221) );
  NR2D1BWP30P140LVT U9127 ( .A1(n10691), .A2(n7830), .ZN(n6222) );
  NR2D1BWP30P140LVT U9128 ( .A1(n10629), .A2(n10965), .ZN(n6223) );
  NR2D1BWP30P140LVT U9129 ( .A1(n8441), .A2(n11103), .ZN(n6224) );
  NR2D1BWP30P140LVT U9130 ( .A1(n6689), .A2(n6412), .ZN(n6225) );
  NR2D1BWP30P140LVT U9131 ( .A1(n7767), .A2(n7733), .ZN(n6226) );
  NR2D1BWP30P140LVT U9132 ( .A1(n10394), .A2(n10962), .ZN(n6227) );
  NR2D1BWP30P140LVT U9133 ( .A1(n10663), .A2(n11183), .ZN(n10360) );
  NR2D1BWP30P140LVT U9134 ( .A1(n10691), .A2(n11131), .ZN(n10006) );
  NR2D1BWP30P140LVT U9135 ( .A1(n10663), .A2(n11112), .ZN(n10026) );
  NR2D1BWP30P140LVT U9136 ( .A1(n10629), .A2(n11150), .ZN(n9969) );
  NR2D1BWP30P140LVT U9137 ( .A1(n10629), .A2(n11011), .ZN(n10116) );
  INR4D1BWP30P140LVT U9138 ( .A1(inner_first_stage_valid_reg[48]), .B1(
        inner_first_stage_valid_reg[55]), .B2(inner_first_stage_valid_reg[54]), 
        .B3(n7375), .ZN(n7376) );
  NR2D1BWP30P140LVT U9139 ( .A1(n8447), .A2(n7430), .ZN(n7443) );
  INVD2BWP30P140LVT U9140 ( .I(n6239), .ZN(n12302) );
  NR2D1BWP30P140LVT U9141 ( .A1(n10394), .A2(n11175), .ZN(n10552) );
  NR2D1BWP30P140LVT U9142 ( .A1(n10663), .A2(n8322), .ZN(n9318) );
  NR2D1BWP30P140LVT U9143 ( .A1(n10663), .A2(n11006), .ZN(n10134) );
  NR2D1BWP30P140LVT U9144 ( .A1(n10691), .A2(n10955), .ZN(n10245) );
  NR2D1BWP30P140LVT U9145 ( .A1(n10691), .A2(n10987), .ZN(n10272) );
  IND2D4BWP30P140LVT U9146 ( .A1(rst), .B1(i_en), .ZN(n6239) );
  NR3D0P7BWP30P140LVT U9147 ( .A1(i_cmd[242]), .A2(i_cmd[234]), .A3(i_cmd[250]), .ZN(n6228) );
  AOI211D1BWP30P140LVT U9148 ( .A1(i_cmd[242]), .A2(n7551), .B(n6228), .C(
        i_cmd[226]), .ZN(n6229) );
  OAI21D1BWP30P140LVT U9149 ( .A1(n7555), .A2(n7552), .B(n6229), .ZN(n6230) );
  INVD2BWP30P140LVT U9150 ( .I(n12302), .ZN(n11181) );
  AOI21D1BWP30P140LVT U9151 ( .A1(n7553), .A2(n6230), .B(n11181), .ZN(N4806)
         );
  NR3D0P7BWP30P140LVT U9152 ( .A1(i_cmd[82]), .A2(i_cmd[74]), .A3(i_cmd[90]), 
        .ZN(n6231) );
  ND2D1BWP30P140LVT U9153 ( .A1(n6231), .A2(i_cmd[66]), .ZN(n8570) );
  AOI211D1BWP30P140LVT U9154 ( .A1(i_cmd[82]), .A2(n8569), .B(n6231), .C(
        i_cmd[66]), .ZN(n6232) );
  OAI21D1BWP30P140LVT U9155 ( .A1(n8566), .A2(n8568), .B(n6232), .ZN(n6233) );
  AOI21D1BWP30P140LVT U9156 ( .A1(n8570), .A2(n6233), .B(n11181), .ZN(N3726)
         );
  NR3D0P7BWP30P140LVT U9157 ( .A1(i_cmd[18]), .A2(i_cmd[10]), .A3(i_cmd[26]), 
        .ZN(n6234) );
  ND2D1BWP30P140LVT U9158 ( .A1(n6234), .A2(i_cmd[2]), .ZN(n8505) );
  AOI211D1BWP30P140LVT U9159 ( .A1(i_cmd[18]), .A2(n8501), .B(n6234), .C(
        i_cmd[2]), .ZN(n6235) );
  OAI21D1BWP30P140LVT U9160 ( .A1(n8504), .A2(n8502), .B(n6235), .ZN(n6236) );
  AOI21D1BWP30P140LVT U9161 ( .A1(n8505), .A2(n6236), .B(n11181), .ZN(N3294)
         );
  NR3D0P7BWP30P140LVT U9162 ( .A1(i_cmd[183]), .A2(i_cmd[175]), .A3(i_cmd[191]), .ZN(n6237) );
  ND2D1BWP30P140LVT U9163 ( .A1(n6237), .A2(i_cmd[167]), .ZN(n6320) );
  AOI211D1BWP30P140LVT U9164 ( .A1(i_cmd[183]), .A2(n6321), .B(n6237), .C(
        i_cmd[167]), .ZN(n6238) );
  OAI21D1BWP30P140LVT U9165 ( .A1(n6322), .A2(n6324), .B(n6238), .ZN(n6240) );
  AOI21D1BWP30P140LVT U9166 ( .A1(n6320), .A2(n6240), .B(n11173), .ZN(N10928)
         );
  NR3D0P7BWP30P140LVT U9167 ( .A1(i_cmd[55]), .A2(i_cmd[47]), .A3(i_cmd[63]), 
        .ZN(n6241) );
  AOI211D1BWP30P140LVT U9168 ( .A1(i_cmd[55]), .A2(n10666), .B(n6241), .C(
        i_cmd[39]), .ZN(n6242) );
  OAI21D1BWP30P140LVT U9169 ( .A1(n10665), .A2(n10669), .B(n6242), .ZN(n6243)
         );
  AOI21D1BWP30P140LVT U9170 ( .A1(n10662), .A2(n6243), .B(n11173), .ZN(N10576)
         );
  NR3D0P7BWP30P140LVT U9171 ( .A1(i_cmd[54]), .A2(i_cmd[46]), .A3(i_cmd[62]), 
        .ZN(n6244) );
  ND2D1BWP30P140LVT U9172 ( .A1(n6244), .A2(i_cmd[38]), .ZN(n8322) );
  OAI21D1BWP30P140LVT U9173 ( .A1(n6244), .A2(i_cmd[38]), .B(n8322), .ZN(n6245) );
  OAI211D1BWP30P140LVT U9174 ( .A1(n8321), .A2(n8319), .B(n10869), .C(n6245), 
        .ZN(n6246) );
  AOI21D1BWP30P140LVT U9175 ( .A1(i_cmd[54]), .A2(n8318), .B(n6246), .ZN(N8958) );
  NR3D0P7BWP30P140LVT U9176 ( .A1(i_cmd[146]), .A2(i_cmd[138]), .A3(i_cmd[154]), .ZN(n6247) );
  OAI21D1BWP30P140LVT U9177 ( .A1(i_cmd[130]), .A2(n6247), .B(n7830), .ZN(
        n6248) );
  OAI211D1BWP30P140LVT U9178 ( .A1(n7829), .A2(n7832), .B(n10869), .C(n6248), 
        .ZN(n6249) );
  AOI21D1BWP30P140LVT U9179 ( .A1(i_cmd[146]), .A2(n7833), .B(n6249), .ZN(
        N4158) );
  NR3D0P7BWP30P140LVT U9180 ( .A1(i_cmd[8]), .A2(i_cmd[24]), .A3(i_cmd[16]), 
        .ZN(n6250) );
  OAI21D1BWP30P140LVT U9181 ( .A1(i_cmd[0]), .A2(n6250), .B(n10374), .ZN(n6251) );
  OAI211D1BWP30P140LVT U9182 ( .A1(n10376), .A2(n10373), .B(n10869), .C(n6251), 
        .ZN(n6252) );
  AOI21D1BWP30P140LVT U9183 ( .A1(i_cmd[16]), .A2(n10372), .B(n6252), .ZN(N542) );
  NR3D0P7BWP30P140LVT U9184 ( .A1(i_cmd[19]), .A2(i_cmd[11]), .A3(i_cmd[27]), 
        .ZN(n6253) );
  OAI21D1BWP30P140LVT U9185 ( .A1(n6253), .A2(i_cmd[3]), .B(n8541), .ZN(n6254)
         );
  OAI211D1BWP30P140LVT U9186 ( .A1(n8537), .A2(n8539), .B(n10869), .C(n6254), 
        .ZN(n6255) );
  AOI21D1BWP30P140LVT U9187 ( .A1(i_cmd[19]), .A2(n8540), .B(n6255), .ZN(N5040) );
  NR2D1BWP30P140LVT U9188 ( .A1(i_cmd[127]), .A2(i_cmd[111]), .ZN(n6256) );
  IND3D1BWP30P140LVT U9189 ( .A1(i_cmd[119]), .B1(i_cmd[103]), .B2(n6256), 
        .ZN(n8374) );
  IND3D1BWP30P140LVT U9190 ( .A1(i_cmd[103]), .B1(i_cmd[119]), .B2(n6256), 
        .ZN(n8375) );
  IND3D1BWP30P140LVT U9191 ( .A1(i_cmd[111]), .B1(i_cmd[127]), .B2(n6257), 
        .ZN(n8376) );
  IND3D1BWP30P140LVT U9192 ( .A1(i_cmd[127]), .B1(i_cmd[111]), .B2(n6257), 
        .ZN(n8377) );
  AN4D0BWP30P140LVT U9193 ( .A1(n8374), .A2(n8375), .A3(n8376), .A4(n8377), 
        .Z(n6258) );
  NR2D1BWP30P140LVT U9194 ( .A1(n6258), .A2(n11057), .ZN(N10752) );
  NR2D1BWP30P140LVT U9195 ( .A1(i_cmd[206]), .A2(i_cmd[222]), .ZN(n6259) );
  IND3D1BWP30P140LVT U9196 ( .A1(i_cmd[198]), .B1(i_cmd[214]), .B2(n6259), 
        .ZN(n7078) );
  NR2D1BWP30P140LVT U9197 ( .A1(i_cmd[198]), .A2(i_cmd[214]), .ZN(n6260) );
  IND3D1BWP30P140LVT U9198 ( .A1(i_cmd[206]), .B1(i_cmd[222]), .B2(n6260), 
        .ZN(n7079) );
  IND3D1BWP30P140LVT U9199 ( .A1(i_cmd[214]), .B1(i_cmd[198]), .B2(n6259), 
        .ZN(n7076) );
  IND3D1BWP30P140LVT U9200 ( .A1(i_cmd[222]), .B1(i_cmd[206]), .B2(n6260), 
        .ZN(n7077) );
  AN4D0BWP30P140LVT U9201 ( .A1(n7078), .A2(n7079), .A3(n7076), .A4(n7077), 
        .Z(n6261) );
  NR2D1BWP30P140LVT U9202 ( .A1(n6261), .A2(n11057), .ZN(N10038) );
  NR2D1BWP30P140LVT U9203 ( .A1(i_cmd[126]), .A2(i_cmd[110]), .ZN(n6263) );
  IND3D1BWP30P140LVT U9204 ( .A1(i_cmd[102]), .B1(i_cmd[118]), .B2(n6263), 
        .ZN(n8420) );
  NR2D1BWP30P140LVT U9205 ( .A1(i_cmd[102]), .A2(i_cmd[118]), .ZN(n6262) );
  IND3D1BWP30P140LVT U9206 ( .A1(i_cmd[126]), .B1(i_cmd[110]), .B2(n6262), 
        .ZN(n8421) );
  IND3D1BWP30P140LVT U9207 ( .A1(i_cmd[110]), .B1(i_cmd[126]), .B2(n6262), 
        .ZN(n8419) );
  IND3D1BWP30P140LVT U9208 ( .A1(i_cmd[118]), .B1(i_cmd[102]), .B2(n6263), 
        .ZN(n8418) );
  AN4D0BWP30P140LVT U9209 ( .A1(n8420), .A2(n8421), .A3(n8419), .A4(n8418), 
        .Z(n6264) );
  NR2D1BWP30P140LVT U9210 ( .A1(n6264), .A2(n11057), .ZN(N9390) );
  IND3D1BWP30P140LVT U9211 ( .A1(i_cmd[236]), .B1(i_cmd[252]), .B2(n6265), 
        .ZN(n7770) );
  IND3D1BWP30P140LVT U9212 ( .A1(i_cmd[252]), .B1(n6265), .B2(i_cmd[236]), 
        .ZN(n7768) );
  IND3D1BWP30P140LVT U9213 ( .A1(i_cmd[244]), .B1(i_cmd[228]), .B2(n6266), 
        .ZN(n7766) );
  IND3D1BWP30P140LVT U9214 ( .A1(i_cmd[228]), .B1(i_cmd[244]), .B2(n6266), 
        .ZN(n7764) );
  AN4D0BWP30P140LVT U9215 ( .A1(n7770), .A2(n7768), .A3(n7766), .A4(n7764), 
        .Z(n12304) );
  IND3D1BWP30P140LVT U9216 ( .A1(i_cmd[248]), .B1(i_cmd[232]), .B2(n6268), 
        .ZN(n7735) );
  IND3D1BWP30P140LVT U9217 ( .A1(i_cmd[224]), .B1(i_cmd[240]), .B2(n6267), 
        .ZN(n7732) );
  IND3D1BWP30P140LVT U9218 ( .A1(i_cmd[240]), .B1(i_cmd[224]), .B2(n6267), 
        .ZN(n7733) );
  IND3D1BWP30P140LVT U9219 ( .A1(i_cmd[232]), .B1(i_cmd[248]), .B2(n6268), 
        .ZN(n7734) );
  AN4D0BWP30P140LVT U9220 ( .A1(n7735), .A2(n7732), .A3(n7733), .A4(n7734), 
        .Z(n6269) );
  NR2D1BWP30P140LVT U9221 ( .A1(n6269), .A2(n11057), .ZN(N2082) );
  NR2D1BWP30P140LVT U9222 ( .A1(i_cmd[108]), .A2(i_cmd[124]), .ZN(n6271) );
  IND3D1BWP30P140LVT U9223 ( .A1(i_cmd[100]), .B1(i_cmd[116]), .B2(n6271), 
        .ZN(n8442) );
  NR2D1BWP30P140LVT U9224 ( .A1(i_cmd[116]), .A2(i_cmd[100]), .ZN(n6270) );
  IND3D1BWP30P140LVT U9225 ( .A1(i_cmd[108]), .B1(i_cmd[124]), .B2(n6270), 
        .ZN(n8446) );
  IND3D1BWP30P140LVT U9226 ( .A1(i_cmd[124]), .B1(i_cmd[108]), .B2(n6270), 
        .ZN(n8444) );
  IND3D1BWP30P140LVT U9227 ( .A1(i_cmd[116]), .B1(n6271), .B2(i_cmd[100]), 
        .ZN(n8440) );
  AN4D0BWP30P140LVT U9228 ( .A1(n8442), .A2(n8446), .A3(n8444), .A4(n8440), 
        .Z(n6272) );
  NR2D1BWP30P140LVT U9229 ( .A1(n6272), .A2(n11057), .ZN(N6666) );
  IND3D1BWP30P140LVT U9230 ( .A1(i_cmd[120]), .B1(i_cmd[104]), .B2(n6273), 
        .ZN(n7428) );
  NR2D1BWP30P140LVT U9231 ( .A1(i_cmd[104]), .A2(i_cmd[120]), .ZN(n6274) );
  IND3D1BWP30P140LVT U9232 ( .A1(i_cmd[96]), .B1(i_cmd[112]), .B2(n6274), .ZN(
        n7431) );
  IND3D1BWP30P140LVT U9233 ( .A1(i_cmd[104]), .B1(n6273), .B2(i_cmd[120]), 
        .ZN(n7430) );
  IND3D1BWP30P140LVT U9234 ( .A1(i_cmd[112]), .B1(i_cmd[96]), .B2(n6274), .ZN(
        n7429) );
  AN4D0BWP30P140LVT U9235 ( .A1(n7428), .A2(n7431), .A3(n7430), .A4(n7429), 
        .Z(n6275) );
  NR2D1BWP30P140LVT U9236 ( .A1(n6275), .A2(n11057), .ZN(N1202) );
  NR2D1BWP30P140LVT U9237 ( .A1(i_cmd[162]), .A2(i_cmd[178]), .ZN(n6277) );
  IND3D1BWP30P140LVT U9238 ( .A1(i_cmd[186]), .B1(i_cmd[170]), .B2(n6277), 
        .ZN(n6411) );
  NR2D1BWP30P140LVT U9239 ( .A1(i_cmd[170]), .A2(i_cmd[186]), .ZN(n6276) );
  IND3D1BWP30P140LVT U9240 ( .A1(i_cmd[162]), .B1(i_cmd[178]), .B2(n6276), 
        .ZN(n6409) );
  IND3D1BWP30P140LVT U9241 ( .A1(i_cmd[178]), .B1(i_cmd[162]), .B2(n6276), 
        .ZN(n6412) );
  IND3D1BWP30P140LVT U9242 ( .A1(i_cmd[170]), .B1(i_cmd[186]), .B2(n6277), 
        .ZN(n6410) );
  AN4D0BWP30P140LVT U9243 ( .A1(n6411), .A2(n6409), .A3(n6412), .A4(n6410), 
        .Z(n6278) );
  NR2D1BWP30P140LVT U9244 ( .A1(n6278), .A2(n11181), .ZN(N4374) );
  NR2D1BWP30P140LVT U9245 ( .A1(i_cmd[97]), .A2(i_cmd[113]), .ZN(n6279) );
  IND3D1BWP30P140LVT U9246 ( .A1(i_cmd[105]), .B1(i_cmd[121]), .B2(n6279), 
        .ZN(n7936) );
  NR2D1BWP30P140LVT U9247 ( .A1(i_cmd[121]), .A2(i_cmd[105]), .ZN(n6280) );
  IND3D1BWP30P140LVT U9248 ( .A1(i_cmd[97]), .B1(i_cmd[113]), .B2(n6280), .ZN(
        n7935) );
  IND3D1BWP30P140LVT U9249 ( .A1(i_cmd[121]), .B1(n6279), .B2(i_cmd[105]), 
        .ZN(n7937) );
  IND3D1BWP30P140LVT U9250 ( .A1(i_cmd[113]), .B1(i_cmd[97]), .B2(n6280), .ZN(
        n7938) );
  AN4D0BWP30P140LVT U9251 ( .A1(n7936), .A2(n7935), .A3(n7937), .A4(n7938), 
        .Z(n6281) );
  NR2D1BWP30P140LVT U9252 ( .A1(n6281), .A2(n11181), .ZN(N2580) );
  NR2D1BWP30P140LVT U9253 ( .A1(i_cmd[177]), .A2(i_cmd[161]), .ZN(n6283) );
  IND3D1BWP30P140LVT U9254 ( .A1(i_cmd[185]), .B1(i_cmd[169]), .B2(n6283), 
        .ZN(n6549) );
  NR2D1BWP30P140LVT U9255 ( .A1(i_cmd[169]), .A2(i_cmd[185]), .ZN(n6282) );
  IND3D1BWP30P140LVT U9256 ( .A1(i_cmd[177]), .B1(i_cmd[161]), .B2(n6282), 
        .ZN(n6548) );
  IND3D1BWP30P140LVT U9257 ( .A1(i_cmd[161]), .B1(i_cmd[177]), .B2(n6282), 
        .ZN(n6550) );
  IND3D1BWP30P140LVT U9258 ( .A1(i_cmd[169]), .B1(i_cmd[185]), .B2(n6283), 
        .ZN(n6551) );
  AN4D0BWP30P140LVT U9259 ( .A1(n6549), .A2(n6548), .A3(n6550), .A4(n6551), 
        .Z(n6284) );
  NR2D1BWP30P140LVT U9260 ( .A1(n6284), .A2(n11181), .ZN(N2756) );
  NR4D1BWP30P140LVT U9261 ( .A1(i_cmd[172]), .A2(n11023), .A3(n6690), .A4(
        n6285), .ZN(n6397) );
  NR4D1BWP30P140LVT U9262 ( .A1(i_cmd[188]), .A2(n6693), .A3(n11022), .A4(
        n6285), .ZN(n6395) );
  AOI22D1BWP30P140LVT U9263 ( .A1(i_data_bus[765]), .A2(n6397), .B1(
        i_data_bus[701]), .B2(n6395), .ZN(n6287) );
  INR4D1BWP30P140LVT U9264 ( .A1(i_cmd[180]), .B1(i_cmd[164]), .B2(n6691), 
        .B3(n11020), .ZN(n6396) );
  NR3D0P7BWP30P140LVT U9265 ( .A1(i_cmd[180]), .A2(i_cmd[188]), .A3(i_cmd[172]), .ZN(n11019) );
  AOI22D1BWP30P140LVT U9266 ( .A1(i_data_bus[733]), .A2(n6396), .B1(
        i_data_bus[669]), .B2(n6398), .ZN(n6286) );
  ND2D1BWP30P140LVT U9267 ( .A1(n6287), .A2(n6286), .ZN(N7128) );
  AOI22D1BWP30P140LVT U9268 ( .A1(i_data_bus[762]), .A2(n6397), .B1(
        i_data_bus[698]), .B2(n6395), .ZN(n6289) );
  AOI22D1BWP30P140LVT U9269 ( .A1(i_data_bus[730]), .A2(n6396), .B1(
        i_data_bus[666]), .B2(n6398), .ZN(n6288) );
  ND2D1BWP30P140LVT U9270 ( .A1(n6289), .A2(n6288), .ZN(N7125) );
  AOI22D1BWP30P140LVT U9271 ( .A1(i_data_bus[673]), .A2(n6395), .B1(
        i_data_bus[705]), .B2(n6396), .ZN(n6291) );
  AOI22D1BWP30P140LVT U9272 ( .A1(i_data_bus[737]), .A2(n6397), .B1(
        i_data_bus[641]), .B2(n6398), .ZN(n6290) );
  ND2D1BWP30P140LVT U9273 ( .A1(n6291), .A2(n6290), .ZN(N7100) );
  AOI22D1BWP30P140LVT U9274 ( .A1(i_data_bus[753]), .A2(n6397), .B1(
        i_data_bus[721]), .B2(n6396), .ZN(n6293) );
  AOI22D1BWP30P140LVT U9275 ( .A1(i_data_bus[689]), .A2(n6395), .B1(
        i_data_bus[657]), .B2(n6398), .ZN(n6292) );
  ND2D1BWP30P140LVT U9276 ( .A1(n6293), .A2(n6292), .ZN(N7116) );
  AOI22D1BWP30P140LVT U9277 ( .A1(i_data_bus[744]), .A2(n6397), .B1(
        i_data_bus[712]), .B2(n6396), .ZN(n6295) );
  AOI22D1BWP30P140LVT U9278 ( .A1(i_data_bus[680]), .A2(n6395), .B1(
        i_data_bus[648]), .B2(n6398), .ZN(n6294) );
  ND2D1BWP30P140LVT U9279 ( .A1(n6295), .A2(n6294), .ZN(N7107) );
  AOI22D1BWP30P140LVT U9280 ( .A1(i_data_bus[738]), .A2(n6397), .B1(
        i_data_bus[706]), .B2(n6396), .ZN(n6297) );
  AOI22D1BWP30P140LVT U9281 ( .A1(i_data_bus[674]), .A2(n6395), .B1(
        i_data_bus[642]), .B2(n6398), .ZN(n6296) );
  ND2D1BWP30P140LVT U9282 ( .A1(n6297), .A2(n6296), .ZN(N7101) );
  AOI22D1BWP30P140LVT U9283 ( .A1(i_data_bus[720]), .A2(n6396), .B1(
        i_data_bus[752]), .B2(n6397), .ZN(n6299) );
  AOI22D1BWP30P140LVT U9284 ( .A1(i_data_bus[688]), .A2(n6395), .B1(
        i_data_bus[656]), .B2(n6398), .ZN(n6298) );
  ND2D1BWP30P140LVT U9285 ( .A1(n6299), .A2(n6298), .ZN(N7115) );
  AOI22D1BWP30P140LVT U9286 ( .A1(i_data_bus[710]), .A2(n6396), .B1(
        i_data_bus[742]), .B2(n6397), .ZN(n6301) );
  AOI22D1BWP30P140LVT U9287 ( .A1(i_data_bus[678]), .A2(n6395), .B1(
        i_data_bus[646]), .B2(n6398), .ZN(n6300) );
  ND2D1BWP30P140LVT U9288 ( .A1(n6301), .A2(n6300), .ZN(N7105) );
  AOI22D1BWP30P140LVT U9289 ( .A1(i_data_bus[734]), .A2(n6396), .B1(
        i_data_bus[670]), .B2(n6398), .ZN(n6303) );
  AOI22D1BWP30P140LVT U9290 ( .A1(i_data_bus[766]), .A2(n6397), .B1(
        i_data_bus[702]), .B2(n6395), .ZN(n6302) );
  ND2D1BWP30P140LVT U9291 ( .A1(n6303), .A2(n6302), .ZN(N7129) );
  AOI22D1BWP30P140LVT U9292 ( .A1(i_data_bus[728]), .A2(n6396), .B1(
        i_data_bus[760]), .B2(n6397), .ZN(n6305) );
  AOI22D1BWP30P140LVT U9293 ( .A1(i_data_bus[664]), .A2(n6398), .B1(
        i_data_bus[696]), .B2(n6395), .ZN(n6304) );
  ND2D1BWP30P140LVT U9294 ( .A1(n6305), .A2(n6304), .ZN(N7123) );
  AOI22D1BWP30P140LVT U9295 ( .A1(i_data_bus[754]), .A2(n6397), .B1(
        i_data_bus[658]), .B2(n6398), .ZN(n6307) );
  AOI22D1BWP30P140LVT U9296 ( .A1(i_data_bus[722]), .A2(n6396), .B1(
        i_data_bus[690]), .B2(n6395), .ZN(n6306) );
  ND2D1BWP30P140LVT U9297 ( .A1(n6307), .A2(n6306), .ZN(N7117) );
  AOI22D1BWP30P140LVT U9298 ( .A1(i_data_bus[652]), .A2(n6398), .B1(
        i_data_bus[748]), .B2(n6397), .ZN(n6309) );
  AOI22D1BWP30P140LVT U9299 ( .A1(i_data_bus[716]), .A2(n6396), .B1(
        i_data_bus[684]), .B2(n6395), .ZN(n6308) );
  ND2D1BWP30P140LVT U9300 ( .A1(n6309), .A2(n6308), .ZN(N7111) );
  AOI22D1BWP30P140LVT U9301 ( .A1(i_data_bus[715]), .A2(n6396), .B1(
        i_data_bus[747]), .B2(n6397), .ZN(n6311) );
  AOI22D1BWP30P140LVT U9302 ( .A1(i_data_bus[651]), .A2(n6398), .B1(
        i_data_bus[683]), .B2(n6395), .ZN(n6310) );
  ND2D1BWP30P140LVT U9303 ( .A1(n6311), .A2(n6310), .ZN(N7110) );
  AOI22D1BWP30P140LVT U9304 ( .A1(i_data_bus[743]), .A2(n6397), .B1(
        i_data_bus[647]), .B2(n6398), .ZN(n6313) );
  AOI22D1BWP30P140LVT U9305 ( .A1(i_data_bus[711]), .A2(n6396), .B1(
        i_data_bus[679]), .B2(n6395), .ZN(n6312) );
  ND2D1BWP30P140LVT U9306 ( .A1(n6313), .A2(n6312), .ZN(N7106) );
  AOI22D1BWP30P140LVT U9307 ( .A1(i_data_bus[741]), .A2(n6397), .B1(
        i_data_bus[645]), .B2(n6398), .ZN(n6315) );
  AOI22D1BWP30P140LVT U9308 ( .A1(i_data_bus[709]), .A2(n6396), .B1(
        i_data_bus[677]), .B2(n6395), .ZN(n6314) );
  ND2D1BWP30P140LVT U9309 ( .A1(n6315), .A2(n6314), .ZN(N7104) );
  AOI22D1BWP30P140LVT U9310 ( .A1(i_data_bus[708]), .A2(n6396), .B1(
        i_data_bus[740]), .B2(n6397), .ZN(n6317) );
  AOI22D1BWP30P140LVT U9311 ( .A1(i_data_bus[644]), .A2(n6398), .B1(
        i_data_bus[676]), .B2(n6395), .ZN(n6316) );
  ND2D1BWP30P140LVT U9312 ( .A1(n6317), .A2(n6316), .ZN(N7103) );
  AOI22D1BWP30P140LVT U9313 ( .A1(i_data_bus[739]), .A2(n6397), .B1(
        i_data_bus[707]), .B2(n6396), .ZN(n6319) );
  AOI22D1BWP30P140LVT U9314 ( .A1(i_data_bus[643]), .A2(n6398), .B1(
        i_data_bus[675]), .B2(n6395), .ZN(n6318) );
  ND2D1BWP30P140LVT U9315 ( .A1(n6319), .A2(n6318), .ZN(N7102) );
  INR4D1BWP30P140LVT U9316 ( .A1(i_cmd[183]), .B1(i_cmd[167]), .B2(n6691), 
        .B3(n6321), .ZN(n6876) );
  AOI22D1BWP30P140LVT U9317 ( .A1(i_data_bus[655]), .A2(n6878), .B1(
        i_data_bus[719]), .B2(n6876), .ZN(n6326) );
  NR4D1BWP30P140LVT U9318 ( .A1(i_cmd[191]), .A2(n6322), .A3(n6693), .A4(n6323), .ZN(n6877) );
  NR4D1BWP30P140LVT U9319 ( .A1(i_cmd[175]), .A2(n6690), .A3(n6324), .A4(n6323), .ZN(n6879) );
  AOI22D1BWP30P140LVT U9320 ( .A1(i_data_bus[687]), .A2(n6877), .B1(
        i_data_bus[751]), .B2(n6879), .ZN(n6325) );
  ND2D1BWP30P140LVT U9321 ( .A1(n6326), .A2(n6325), .ZN(N10944) );
  AOI22D1BWP30P140LVT U9322 ( .A1(i_data_bus[668]), .A2(n6398), .B1(
        i_data_bus[700]), .B2(n6395), .ZN(n6328) );
  AOI22D1BWP30P140LVT U9323 ( .A1(i_data_bus[764]), .A2(n6397), .B1(
        i_data_bus[732]), .B2(n6396), .ZN(n6327) );
  ND2D1BWP30P140LVT U9324 ( .A1(n6328), .A2(n6327), .ZN(N7127) );
  AOI22D1BWP30P140LVT U9325 ( .A1(i_data_bus[761]), .A2(n6397), .B1(
        i_data_bus[665]), .B2(n6398), .ZN(n6330) );
  AOI22D1BWP30P140LVT U9326 ( .A1(i_data_bus[697]), .A2(n6395), .B1(
        i_data_bus[729]), .B2(n6396), .ZN(n6329) );
  ND2D1BWP30P140LVT U9327 ( .A1(n6330), .A2(n6329), .ZN(N7124) );
  AOI22D1BWP30P140LVT U9328 ( .A1(i_data_bus[663]), .A2(n6398), .B1(
        i_data_bus[695]), .B2(n6395), .ZN(n6332) );
  AOI22D1BWP30P140LVT U9329 ( .A1(i_data_bus[759]), .A2(n6397), .B1(
        i_data_bus[727]), .B2(n6396), .ZN(n6331) );
  ND2D1BWP30P140LVT U9330 ( .A1(n6332), .A2(n6331), .ZN(N7122) );
  AOI22D1BWP30P140LVT U9331 ( .A1(i_data_bus[659]), .A2(n6398), .B1(
        i_data_bus[691]), .B2(n6395), .ZN(n6334) );
  AOI22D1BWP30P140LVT U9332 ( .A1(i_data_bus[755]), .A2(n6397), .B1(
        i_data_bus[723]), .B2(n6396), .ZN(n6333) );
  ND2D1BWP30P140LVT U9333 ( .A1(n6334), .A2(n6333), .ZN(N7118) );
  AOI22D1BWP30P140LVT U9334 ( .A1(i_data_bus[653]), .A2(n6398), .B1(
        i_data_bus[749]), .B2(n6397), .ZN(n6336) );
  AOI22D1BWP30P140LVT U9335 ( .A1(i_data_bus[685]), .A2(n6395), .B1(
        i_data_bus[717]), .B2(n6396), .ZN(n6335) );
  ND2D1BWP30P140LVT U9336 ( .A1(n6336), .A2(n6335), .ZN(N7112) );
  AOI22D1BWP30P140LVT U9337 ( .A1(i_data_bus[746]), .A2(n6397), .B1(
        i_data_bus[682]), .B2(n6395), .ZN(n6338) );
  AOI22D1BWP30P140LVT U9338 ( .A1(i_data_bus[650]), .A2(n6398), .B1(
        i_data_bus[714]), .B2(n6396), .ZN(n6337) );
  ND2D1BWP30P140LVT U9339 ( .A1(n6338), .A2(n6337), .ZN(N7109) );
  AOI22D1BWP30P140LVT U9340 ( .A1(i_data_bus[681]), .A2(n6395), .B1(
        i_data_bus[745]), .B2(n6397), .ZN(n6340) );
  AOI22D1BWP30P140LVT U9341 ( .A1(i_data_bus[649]), .A2(n6398), .B1(
        i_data_bus[713]), .B2(n6396), .ZN(n6339) );
  ND2D1BWP30P140LVT U9342 ( .A1(n6340), .A2(n6339), .ZN(N7108) );
  OR2D1BWP30P140LVT U9343 ( .A1(i_cmd[204]), .A2(i_cmd[220]), .Z(n11018) );
  INR4D1BWP30P140LVT U9344 ( .A1(i_cmd[212]), .B1(i_cmd[196]), .B2(n7181), 
        .B3(n11018), .ZN(n6760) );
  INR4D1BWP30P140LVT U9345 ( .A1(i_cmd[220]), .B1(i_cmd[204]), .B2(n7179), 
        .B3(n6341), .ZN(n6761) );
  AOI22D1BWP30P140LVT U9346 ( .A1(i_data_bus[852]), .A2(n6760), .B1(
        i_data_bus[884]), .B2(n6761), .ZN(n6343) );
  INR4D1BWP30P140LVT U9347 ( .A1(i_cmd[204]), .B1(i_cmd[220]), .B2(n7183), 
        .B3(n6341), .ZN(n6759) );
  NR3D0P7BWP30P140LVT U9348 ( .A1(i_cmd[212]), .A2(i_cmd[204]), .A3(i_cmd[220]), .ZN(n11014) );
  ND2D1BWP30P140LVT U9349 ( .A1(n11014), .A2(i_cmd[196]), .ZN(n11016) );
  AOI22D1BWP30P140LVT U9350 ( .A1(i_data_bus[820]), .A2(n6759), .B1(
        i_data_bus[788]), .B2(n6758), .ZN(n6342) );
  ND2D1BWP30P140LVT U9351 ( .A1(n6343), .A2(n6342), .ZN(N7335) );
  AOI22D1BWP30P140LVT U9352 ( .A1(i_data_bus[813]), .A2(n6759), .B1(
        i_data_bus[877]), .B2(n6761), .ZN(n6345) );
  AOI22D1BWP30P140LVT U9353 ( .A1(i_data_bus[845]), .A2(n6760), .B1(
        i_data_bus[781]), .B2(n6758), .ZN(n6344) );
  ND2D1BWP30P140LVT U9354 ( .A1(n6345), .A2(n6344), .ZN(N7328) );
  AOI22D1BWP30P140LVT U9355 ( .A1(i_data_bus[812]), .A2(n6759), .B1(
        i_data_bus[876]), .B2(n6761), .ZN(n6347) );
  AOI22D1BWP30P140LVT U9356 ( .A1(i_data_bus[844]), .A2(n6760), .B1(
        i_data_bus[780]), .B2(n6758), .ZN(n6346) );
  ND2D1BWP30P140LVT U9357 ( .A1(n6347), .A2(n6346), .ZN(N7327) );
  NR3D0P7BWP30P140LVT U9358 ( .A1(i_cmd[173]), .A2(i_cmd[189]), .A3(i_cmd[181]), .ZN(n10978) );
  INR4D1BWP30P140LVT U9359 ( .A1(i_cmd[181]), .B1(i_cmd[165]), .B2(n6691), 
        .B3(n10979), .ZN(n6883) );
  AOI22D1BWP30P140LVT U9360 ( .A1(i_data_bus[667]), .A2(n6884), .B1(
        i_data_bus[731]), .B2(n6883), .ZN(n6350) );
  NR4D1BWP30P140LVT U9361 ( .A1(i_cmd[189]), .A2(n10982), .A3(n6693), .A4(
        n6348), .ZN(n6882) );
  NR4D1BWP30P140LVT U9362 ( .A1(i_cmd[173]), .A2(n6690), .A3(n10981), .A4(
        n6348), .ZN(n6885) );
  AOI22D1BWP30P140LVT U9363 ( .A1(i_data_bus[699]), .A2(n6882), .B1(
        i_data_bus[763]), .B2(n6885), .ZN(n6349) );
  ND2D1BWP30P140LVT U9364 ( .A1(n6350), .A2(n6349), .ZN(N8232) );
  AOI22D1BWP30P140LVT U9365 ( .A1(i_data_bus[664]), .A2(n6884), .B1(
        i_data_bus[696]), .B2(n6882), .ZN(n6352) );
  AOI22D1BWP30P140LVT U9366 ( .A1(i_data_bus[728]), .A2(n6883), .B1(
        i_data_bus[760]), .B2(n6885), .ZN(n6351) );
  ND2D1BWP30P140LVT U9367 ( .A1(n6352), .A2(n6351), .ZN(N8229) );
  AOI22D1BWP30P140LVT U9368 ( .A1(i_data_bus[655]), .A2(n6884), .B1(
        i_data_bus[687]), .B2(n6882), .ZN(n6354) );
  AOI22D1BWP30P140LVT U9369 ( .A1(i_data_bus[719]), .A2(n6883), .B1(
        i_data_bus[751]), .B2(n6885), .ZN(n6353) );
  ND2D1BWP30P140LVT U9370 ( .A1(n6354), .A2(n6353), .ZN(N8220) );
  AOI22D1BWP30P140LVT U9371 ( .A1(i_data_bus[654]), .A2(n6884), .B1(
        i_data_bus[718]), .B2(n6883), .ZN(n6356) );
  AOI22D1BWP30P140LVT U9372 ( .A1(i_data_bus[686]), .A2(n6882), .B1(
        i_data_bus[750]), .B2(n6885), .ZN(n6355) );
  ND2D1BWP30P140LVT U9373 ( .A1(n6356), .A2(n6355), .ZN(N8219) );
  NR3D0P7BWP30P140LVT U9374 ( .A1(i_cmd[171]), .A2(i_cmd[187]), .A3(i_cmd[179]), .ZN(n11065) );
  OR2D1BWP30P140LVT U9375 ( .A1(i_cmd[171]), .A2(i_cmd[187]), .Z(n11069) );
  INR4D1BWP30P140LVT U9376 ( .A1(i_cmd[179]), .B1(i_cmd[163]), .B2(n6691), 
        .B3(n11069), .ZN(n6911) );
  AOI22D1BWP30P140LVT U9377 ( .A1(i_data_bus[653]), .A2(n6910), .B1(
        i_data_bus[717]), .B2(n6911), .ZN(n6359) );
  INR4D1BWP30P140LVT U9378 ( .A1(i_cmd[171]), .B1(i_cmd[187]), .B2(n6693), 
        .B3(n6357), .ZN(n6909) );
  INR4D1BWP30P140LVT U9379 ( .A1(i_cmd[187]), .B1(i_cmd[171]), .B2(n6690), 
        .B3(n6357), .ZN(n6908) );
  AOI22D1BWP30P140LVT U9380 ( .A1(i_data_bus[685]), .A2(n6909), .B1(
        i_data_bus[749]), .B2(n6908), .ZN(n6358) );
  ND2D1BWP30P140LVT U9381 ( .A1(n6359), .A2(n6358), .ZN(N5494) );
  AOI22D1BWP30P140LVT U9382 ( .A1(i_data_bus[651]), .A2(n6910), .B1(
        i_data_bus[683]), .B2(n6909), .ZN(n6361) );
  AOI22D1BWP30P140LVT U9383 ( .A1(i_data_bus[715]), .A2(n6911), .B1(
        i_data_bus[747]), .B2(n6908), .ZN(n6360) );
  ND2D1BWP30P140LVT U9384 ( .A1(n6361), .A2(n6360), .ZN(N5492) );
  AOI22D1BWP30P140LVT U9385 ( .A1(i_data_bus[650]), .A2(n6910), .B1(
        i_data_bus[682]), .B2(n6909), .ZN(n6363) );
  AOI22D1BWP30P140LVT U9386 ( .A1(i_data_bus[746]), .A2(n6908), .B1(
        i_data_bus[714]), .B2(n6911), .ZN(n6362) );
  ND2D1BWP30P140LVT U9387 ( .A1(n6363), .A2(n6362), .ZN(N5491) );
  AOI22D1BWP30P140LVT U9388 ( .A1(i_data_bus[670]), .A2(n6878), .B1(
        i_data_bus[702]), .B2(n6877), .ZN(n6365) );
  AOI22D1BWP30P140LVT U9389 ( .A1(i_data_bus[766]), .A2(n6879), .B1(
        i_data_bus[734]), .B2(n6876), .ZN(n6364) );
  ND2D1BWP30P140LVT U9390 ( .A1(n6365), .A2(n6364), .ZN(N10959) );
  AOI22D1BWP30P140LVT U9391 ( .A1(i_data_bus[654]), .A2(n6878), .B1(
        i_data_bus[686]), .B2(n6877), .ZN(n6367) );
  AOI22D1BWP30P140LVT U9392 ( .A1(i_data_bus[750]), .A2(n6879), .B1(
        i_data_bus[718]), .B2(n6876), .ZN(n6366) );
  ND2D1BWP30P140LVT U9393 ( .A1(n6367), .A2(n6366), .ZN(N10943) );
  AOI22D1BWP30P140LVT U9394 ( .A1(i_data_bus[650]), .A2(n6878), .B1(
        i_data_bus[746]), .B2(n6879), .ZN(n6369) );
  AOI22D1BWP30P140LVT U9395 ( .A1(i_data_bus[682]), .A2(n6877), .B1(
        i_data_bus[714]), .B2(n6876), .ZN(n6368) );
  ND2D1BWP30P140LVT U9396 ( .A1(n6369), .A2(n6368), .ZN(N10939) );
  NR3D0P7BWP30P140LVT U9397 ( .A1(i_cmd[174]), .A2(i_cmd[190]), .A3(i_cmd[182]), .ZN(n10944) );
  INR4D1BWP30P140LVT U9398 ( .A1(i_cmd[174]), .B1(i_cmd[190]), .B2(n6693), 
        .B3(n6370), .ZN(n6923) );
  AOI22D1BWP30P140LVT U9399 ( .A1(i_data_bus[670]), .A2(n6924), .B1(
        i_data_bus[702]), .B2(n6923), .ZN(n6372) );
  INR4D1BWP30P140LVT U9400 ( .A1(i_cmd[190]), .B1(i_cmd[174]), .B2(n6690), 
        .B3(n6370), .ZN(n6925) );
  OR2D1BWP30P140LVT U9401 ( .A1(i_cmd[174]), .A2(i_cmd[190]), .Z(n10948) );
  INR4D1BWP30P140LVT U9402 ( .A1(i_cmd[182]), .B1(i_cmd[166]), .B2(n6691), 
        .B3(n10948), .ZN(n6922) );
  AOI22D1BWP30P140LVT U9403 ( .A1(i_data_bus[766]), .A2(n6925), .B1(
        i_data_bus[734]), .B2(n6922), .ZN(n6371) );
  ND2D1BWP30P140LVT U9404 ( .A1(n6372), .A2(n6371), .ZN(N9853) );
  AOI22D1BWP30P140LVT U9405 ( .A1(i_data_bus[668]), .A2(n6924), .B1(
        i_data_bus[700]), .B2(n6923), .ZN(n6374) );
  AOI22D1BWP30P140LVT U9406 ( .A1(i_data_bus[764]), .A2(n6925), .B1(
        i_data_bus[732]), .B2(n6922), .ZN(n6373) );
  ND2D1BWP30P140LVT U9407 ( .A1(n6374), .A2(n6373), .ZN(N9851) );
  AOI22D1BWP30P140LVT U9408 ( .A1(i_data_bus[663]), .A2(n6924), .B1(
        i_data_bus[695]), .B2(n6923), .ZN(n6376) );
  AOI22D1BWP30P140LVT U9409 ( .A1(i_data_bus[759]), .A2(n6925), .B1(
        i_data_bus[727]), .B2(n6922), .ZN(n6375) );
  ND2D1BWP30P140LVT U9410 ( .A1(n6376), .A2(n6375), .ZN(N9846) );
  AOI22D1BWP30P140LVT U9411 ( .A1(i_data_bus[653]), .A2(n6924), .B1(
        i_data_bus[717]), .B2(n6922), .ZN(n6378) );
  AOI22D1BWP30P140LVT U9412 ( .A1(i_data_bus[685]), .A2(n6923), .B1(
        i_data_bus[749]), .B2(n6925), .ZN(n6377) );
  ND2D1BWP30P140LVT U9413 ( .A1(n6378), .A2(n6377), .ZN(N9836) );
  AOI22D1BWP30P140LVT U9414 ( .A1(i_data_bus[652]), .A2(n6924), .B1(
        i_data_bus[684]), .B2(n6923), .ZN(n6380) );
  AOI22D1BWP30P140LVT U9415 ( .A1(i_data_bus[716]), .A2(n6922), .B1(
        i_data_bus[748]), .B2(n6925), .ZN(n6379) );
  ND2D1BWP30P140LVT U9416 ( .A1(n6380), .A2(n6379), .ZN(N9835) );
  AOI22D1BWP30P140LVT U9417 ( .A1(i_data_bus[735]), .A2(n6396), .B1(
        i_data_bus[671]), .B2(n6398), .ZN(n6382) );
  AOI22D1BWP30P140LVT U9418 ( .A1(i_data_bus[703]), .A2(n6395), .B1(
        i_data_bus[767]), .B2(n6397), .ZN(n6381) );
  ND2D1BWP30P140LVT U9419 ( .A1(n6382), .A2(n6381), .ZN(N7130) );
  AOI22D1BWP30P140LVT U9420 ( .A1(i_data_bus[667]), .A2(n6398), .B1(
        i_data_bus[699]), .B2(n6395), .ZN(n6384) );
  AOI22D1BWP30P140LVT U9421 ( .A1(i_data_bus[731]), .A2(n6396), .B1(
        i_data_bus[763]), .B2(n6397), .ZN(n6383) );
  ND2D1BWP30P140LVT U9422 ( .A1(n6384), .A2(n6383), .ZN(N7126) );
  AOI22D1BWP30P140LVT U9423 ( .A1(i_data_bus[694]), .A2(n6395), .B1(
        i_data_bus[726]), .B2(n6396), .ZN(n6386) );
  AOI22D1BWP30P140LVT U9424 ( .A1(i_data_bus[662]), .A2(n6398), .B1(
        i_data_bus[758]), .B2(n6397), .ZN(n6385) );
  ND2D1BWP30P140LVT U9425 ( .A1(n6386), .A2(n6385), .ZN(N7121) );
  AOI22D1BWP30P140LVT U9426 ( .A1(i_data_bus[725]), .A2(n6396), .B1(
        i_data_bus[661]), .B2(n6398), .ZN(n6388) );
  AOI22D1BWP30P140LVT U9427 ( .A1(i_data_bus[693]), .A2(n6395), .B1(
        i_data_bus[757]), .B2(n6397), .ZN(n6387) );
  ND2D1BWP30P140LVT U9428 ( .A1(n6388), .A2(n6387), .ZN(N7120) );
  AOI22D1BWP30P140LVT U9429 ( .A1(i_data_bus[724]), .A2(n6396), .B1(
        i_data_bus[660]), .B2(n6398), .ZN(n6390) );
  AOI22D1BWP30P140LVT U9430 ( .A1(i_data_bus[692]), .A2(n6395), .B1(
        i_data_bus[756]), .B2(n6397), .ZN(n6389) );
  ND2D1BWP30P140LVT U9431 ( .A1(n6390), .A2(n6389), .ZN(N7119) );
  AOI22D1BWP30P140LVT U9432 ( .A1(i_data_bus[687]), .A2(n6395), .B1(
        i_data_bus[719]), .B2(n6396), .ZN(n6392) );
  AOI22D1BWP30P140LVT U9433 ( .A1(i_data_bus[655]), .A2(n6398), .B1(
        i_data_bus[751]), .B2(n6397), .ZN(n6391) );
  ND2D1BWP30P140LVT U9434 ( .A1(n6392), .A2(n6391), .ZN(N7114) );
  AOI22D1BWP30P140LVT U9435 ( .A1(i_data_bus[654]), .A2(n6398), .B1(
        i_data_bus[718]), .B2(n6396), .ZN(n6394) );
  AOI22D1BWP30P140LVT U9436 ( .A1(i_data_bus[686]), .A2(n6395), .B1(
        i_data_bus[750]), .B2(n6397), .ZN(n6393) );
  ND2D1BWP30P140LVT U9437 ( .A1(n6394), .A2(n6393), .ZN(N7113) );
  AOI22D1BWP30P140LVT U9438 ( .A1(i_data_bus[704]), .A2(n6396), .B1(
        i_data_bus[672]), .B2(n6395), .ZN(n6400) );
  AOI22D1BWP30P140LVT U9439 ( .A1(i_data_bus[640]), .A2(n6398), .B1(
        i_data_bus[736]), .B2(n6397), .ZN(n6399) );
  ND2D1BWP30P140LVT U9440 ( .A1(n6400), .A2(n6399), .ZN(N7099) );
  AOI22D1BWP30P140LVT U9441 ( .A1(i_data_bus[664]), .A2(n6910), .B1(
        i_data_bus[728]), .B2(n6911), .ZN(n6402) );
  AOI22D1BWP30P140LVT U9442 ( .A1(i_data_bus[760]), .A2(n6908), .B1(
        i_data_bus[696]), .B2(n6909), .ZN(n6401) );
  ND2D1BWP30P140LVT U9443 ( .A1(n6402), .A2(n6401), .ZN(N5505) );
  AOI22D1BWP30P140LVT U9444 ( .A1(i_data_bus[663]), .A2(n6910), .B1(
        i_data_bus[727]), .B2(n6911), .ZN(n6404) );
  AOI22D1BWP30P140LVT U9445 ( .A1(i_data_bus[759]), .A2(n6908), .B1(
        i_data_bus[695]), .B2(n6909), .ZN(n6403) );
  ND2D1BWP30P140LVT U9446 ( .A1(n6404), .A2(n6403), .ZN(N5504) );
  AOI22D1BWP30P140LVT U9447 ( .A1(i_data_bus[659]), .A2(n6910), .B1(
        i_data_bus[723]), .B2(n6911), .ZN(n6406) );
  AOI22D1BWP30P140LVT U9448 ( .A1(i_data_bus[755]), .A2(n6908), .B1(
        i_data_bus[691]), .B2(n6909), .ZN(n6405) );
  ND2D1BWP30P140LVT U9449 ( .A1(n6406), .A2(n6405), .ZN(N5500) );
  AOI22D1BWP30P140LVT U9450 ( .A1(i_data_bus[652]), .A2(n6910), .B1(
        i_data_bus[748]), .B2(n6908), .ZN(n6408) );
  AOI22D1BWP30P140LVT U9451 ( .A1(i_data_bus[716]), .A2(n6911), .B1(
        i_data_bus[684]), .B2(n6909), .ZN(n6407) );
  ND2D1BWP30P140LVT U9452 ( .A1(n6408), .A2(n6407), .ZN(N5493) );
  AOI22D1BWP30P140LVT U9453 ( .A1(i_data_bus[709]), .A2(n6619), .B1(
        i_data_bus[741]), .B2(n6618), .ZN(n6414) );
  AOI22D1BWP30P140LVT U9454 ( .A1(i_data_bus[677]), .A2(n6620), .B1(
        i_data_bus[645]), .B2(n6225), .ZN(n6413) );
  ND2D1BWP30P140LVT U9455 ( .A1(n6414), .A2(n6413), .ZN(N4380) );
  AOI22D1BWP30P140LVT U9456 ( .A1(i_data_bus[693]), .A2(n6620), .B1(
        i_data_bus[757]), .B2(n6618), .ZN(n6416) );
  AOI22D1BWP30P140LVT U9457 ( .A1(i_data_bus[725]), .A2(n6619), .B1(
        i_data_bus[661]), .B2(n6225), .ZN(n6415) );
  ND2D1BWP30P140LVT U9458 ( .A1(n6416), .A2(n6415), .ZN(N4396) );
  INVD1BWP30P140LVT U9459 ( .I(i_cmd[219]), .ZN(n6417) );
  INVD1BWP30P140LVT U9460 ( .I(i_cmd[203]), .ZN(n6419) );
  INR4D1BWP30P140LVT U9461 ( .A1(i_cmd[211]), .B1(i_cmd[195]), .B2(n7181), 
        .B3(n11064), .ZN(n6722) );
  NR4D1BWP30P140LVT U9462 ( .A1(i_cmd[203]), .A2(n6417), .A3(n7179), .A4(n6418), .ZN(n6723) );
  AOI22D1BWP30P140LVT U9463 ( .A1(i_data_bus[852]), .A2(n6722), .B1(
        i_data_bus[884]), .B2(n6723), .ZN(n6421) );
  NR3D0P7BWP30P140LVT U9464 ( .A1(i_cmd[211]), .A2(i_cmd[219]), .A3(i_cmd[203]), .ZN(n11060) );
  AOI22D1BWP30P140LVT U9465 ( .A1(i_data_bus[820]), .A2(n6721), .B1(
        i_data_bus[788]), .B2(n6720), .ZN(n6420) );
  ND2D1BWP30P140LVT U9466 ( .A1(n6421), .A2(n6420), .ZN(N5589) );
  AOI22D1BWP30P140LVT U9467 ( .A1(i_data_bus[812]), .A2(n6721), .B1(
        i_data_bus[876]), .B2(n6723), .ZN(n6423) );
  AOI22D1BWP30P140LVT U9468 ( .A1(i_data_bus[844]), .A2(n6722), .B1(
        i_data_bus[780]), .B2(n6720), .ZN(n6422) );
  ND2D1BWP30P140LVT U9469 ( .A1(n6423), .A2(n6422), .ZN(N5581) );
  AOI22D1BWP30P140LVT U9470 ( .A1(i_data_bus[659]), .A2(n6924), .B1(
        i_data_bus[755]), .B2(n6925), .ZN(n6425) );
  AOI22D1BWP30P140LVT U9471 ( .A1(i_data_bus[723]), .A2(n6922), .B1(
        i_data_bus[691]), .B2(n6923), .ZN(n6424) );
  ND2D1BWP30P140LVT U9472 ( .A1(n6425), .A2(n6424), .ZN(N9842) );
  AOI22D1BWP30P140LVT U9473 ( .A1(i_data_bus[650]), .A2(n6924), .B1(
        i_data_bus[714]), .B2(n6922), .ZN(n6427) );
  AOI22D1BWP30P140LVT U9474 ( .A1(i_data_bus[746]), .A2(n6925), .B1(
        i_data_bus[682]), .B2(n6923), .ZN(n6426) );
  ND2D1BWP30P140LVT U9475 ( .A1(n6427), .A2(n6426), .ZN(N9833) );
  AOI22D1BWP30P140LVT U9476 ( .A1(i_data_bus[668]), .A2(n6884), .B1(
        i_data_bus[764]), .B2(n6885), .ZN(n6429) );
  AOI22D1BWP30P140LVT U9477 ( .A1(i_data_bus[732]), .A2(n6883), .B1(
        i_data_bus[700]), .B2(n6882), .ZN(n6428) );
  ND2D1BWP30P140LVT U9478 ( .A1(n6429), .A2(n6428), .ZN(N8233) );
  AOI22D1BWP30P140LVT U9479 ( .A1(i_data_bus[663]), .A2(n6884), .B1(
        i_data_bus[759]), .B2(n6885), .ZN(n6431) );
  AOI22D1BWP30P140LVT U9480 ( .A1(i_data_bus[727]), .A2(n6883), .B1(
        i_data_bus[695]), .B2(n6882), .ZN(n6430) );
  ND2D1BWP30P140LVT U9481 ( .A1(n6431), .A2(n6430), .ZN(N8228) );
  AOI22D1BWP30P140LVT U9482 ( .A1(i_data_bus[659]), .A2(n6884), .B1(
        i_data_bus[723]), .B2(n6883), .ZN(n6433) );
  AOI22D1BWP30P140LVT U9483 ( .A1(i_data_bus[755]), .A2(n6885), .B1(
        i_data_bus[691]), .B2(n6882), .ZN(n6432) );
  ND2D1BWP30P140LVT U9484 ( .A1(n6433), .A2(n6432), .ZN(N8224) );
  AOI22D1BWP30P140LVT U9485 ( .A1(i_data_bus[668]), .A2(n6878), .B1(
        i_data_bus[732]), .B2(n6876), .ZN(n6435) );
  AOI22D1BWP30P140LVT U9486 ( .A1(i_data_bus[764]), .A2(n6879), .B1(
        i_data_bus[700]), .B2(n6877), .ZN(n6434) );
  ND2D1BWP30P140LVT U9487 ( .A1(n6435), .A2(n6434), .ZN(N10957) );
  AOI22D1BWP30P140LVT U9488 ( .A1(i_data_bus[663]), .A2(n6878), .B1(
        i_data_bus[727]), .B2(n6876), .ZN(n6437) );
  AOI22D1BWP30P140LVT U9489 ( .A1(i_data_bus[759]), .A2(n6879), .B1(
        i_data_bus[695]), .B2(n6877), .ZN(n6436) );
  ND2D1BWP30P140LVT U9490 ( .A1(n6437), .A2(n6436), .ZN(N10952) );
  AOI22D1BWP30P140LVT U9491 ( .A1(i_data_bus[661]), .A2(n6878), .B1(
        i_data_bus[757]), .B2(n6879), .ZN(n6439) );
  AOI22D1BWP30P140LVT U9492 ( .A1(i_data_bus[725]), .A2(n6876), .B1(
        i_data_bus[693]), .B2(n6877), .ZN(n6438) );
  ND2D1BWP30P140LVT U9493 ( .A1(n6439), .A2(n6438), .ZN(N10950) );
  AOI22D1BWP30P140LVT U9494 ( .A1(i_data_bus[641]), .A2(n6878), .B1(
        i_data_bus[705]), .B2(n6876), .ZN(n6441) );
  AOI22D1BWP30P140LVT U9495 ( .A1(i_data_bus[737]), .A2(n6879), .B1(
        i_data_bus[673]), .B2(n6877), .ZN(n6440) );
  ND2D1BWP30P140LVT U9496 ( .A1(n6441), .A2(n6440), .ZN(N10930) );
  AOI22D1BWP30P140LVT U9497 ( .A1(i_data_bus[766]), .A2(n6618), .B1(
        i_data_bus[702]), .B2(n6620), .ZN(n6443) );
  AOI22D1BWP30P140LVT U9498 ( .A1(i_data_bus[734]), .A2(n6619), .B1(
        i_data_bus[670]), .B2(n6225), .ZN(n6442) );
  ND2D1BWP30P140LVT U9499 ( .A1(n6443), .A2(n6442), .ZN(N4405) );
  AOI22D1BWP30P140LVT U9500 ( .A1(i_data_bus[765]), .A2(n6618), .B1(
        i_data_bus[701]), .B2(n6620), .ZN(n6445) );
  AOI22D1BWP30P140LVT U9501 ( .A1(i_data_bus[733]), .A2(n6619), .B1(
        i_data_bus[669]), .B2(n6225), .ZN(n6444) );
  ND2D1BWP30P140LVT U9502 ( .A1(n6445), .A2(n6444), .ZN(N4404) );
  AOI22D1BWP30P140LVT U9503 ( .A1(i_data_bus[740]), .A2(n6618), .B1(
        i_data_bus[676]), .B2(n6620), .ZN(n6447) );
  AOI22D1BWP30P140LVT U9504 ( .A1(i_data_bus[708]), .A2(n6619), .B1(
        i_data_bus[644]), .B2(n6225), .ZN(n6446) );
  ND2D1BWP30P140LVT U9505 ( .A1(n6447), .A2(n6446), .ZN(N4379) );
  AOI22D1BWP30P140LVT U9506 ( .A1(i_data_bus[761]), .A2(n6618), .B1(
        i_data_bus[729]), .B2(n6619), .ZN(n6449) );
  AOI22D1BWP30P140LVT U9507 ( .A1(i_data_bus[697]), .A2(n6620), .B1(
        i_data_bus[665]), .B2(n6225), .ZN(n6448) );
  ND2D1BWP30P140LVT U9508 ( .A1(n6449), .A2(n6448), .ZN(N4400) );
  AOI22D1BWP30P140LVT U9509 ( .A1(i_data_bus[753]), .A2(n6618), .B1(
        i_data_bus[721]), .B2(n6619), .ZN(n6451) );
  AOI22D1BWP30P140LVT U9510 ( .A1(i_data_bus[689]), .A2(n6620), .B1(
        i_data_bus[657]), .B2(n6225), .ZN(n6450) );
  ND2D1BWP30P140LVT U9511 ( .A1(n6451), .A2(n6450), .ZN(N4392) );
  AOI22D1BWP30P140LVT U9512 ( .A1(i_data_bus[737]), .A2(n6618), .B1(
        i_data_bus[705]), .B2(n6619), .ZN(n6453) );
  AOI22D1BWP30P140LVT U9513 ( .A1(i_data_bus[673]), .A2(n6620), .B1(
        i_data_bus[641]), .B2(n6225), .ZN(n6452) );
  ND2D1BWP30P140LVT U9514 ( .A1(n6453), .A2(n6452), .ZN(N4376) );
  AOI22D1BWP30P140LVT U9515 ( .A1(i_data_bus[847]), .A2(n6760), .B1(
        i_data_bus[783]), .B2(n6758), .ZN(n6455) );
  AOI22D1BWP30P140LVT U9516 ( .A1(i_data_bus[815]), .A2(n6759), .B1(
        i_data_bus[879]), .B2(n6761), .ZN(n6454) );
  ND2D1BWP30P140LVT U9517 ( .A1(n6455), .A2(n6454), .ZN(N7330) );
  AOI22D1BWP30P140LVT U9518 ( .A1(i_data_bus[731]), .A2(n6876), .B1(
        i_data_bus[763]), .B2(n6879), .ZN(n6457) );
  AOI22D1BWP30P140LVT U9519 ( .A1(i_data_bus[667]), .A2(n6878), .B1(
        i_data_bus[699]), .B2(n6877), .ZN(n6456) );
  ND2D1BWP30P140LVT U9520 ( .A1(n6457), .A2(n6456), .ZN(N10956) );
  AOI22D1BWP30P140LVT U9521 ( .A1(i_data_bus[728]), .A2(n6876), .B1(
        i_data_bus[696]), .B2(n6877), .ZN(n6459) );
  AOI22D1BWP30P140LVT U9522 ( .A1(i_data_bus[664]), .A2(n6878), .B1(
        i_data_bus[760]), .B2(n6879), .ZN(n6458) );
  ND2D1BWP30P140LVT U9523 ( .A1(n6459), .A2(n6458), .ZN(N10953) );
  AOI22D1BWP30P140LVT U9524 ( .A1(i_data_bus[758]), .A2(n6879), .B1(
        i_data_bus[726]), .B2(n6876), .ZN(n6461) );
  AOI22D1BWP30P140LVT U9525 ( .A1(i_data_bus[662]), .A2(n6878), .B1(
        i_data_bus[694]), .B2(n6877), .ZN(n6460) );
  ND2D1BWP30P140LVT U9526 ( .A1(n6461), .A2(n6460), .ZN(N10951) );
  AOI22D1BWP30P140LVT U9527 ( .A1(i_data_bus[692]), .A2(n6877), .B1(
        i_data_bus[724]), .B2(n6876), .ZN(n6463) );
  AOI22D1BWP30P140LVT U9528 ( .A1(i_data_bus[660]), .A2(n6878), .B1(
        i_data_bus[756]), .B2(n6879), .ZN(n6462) );
  ND2D1BWP30P140LVT U9529 ( .A1(n6463), .A2(n6462), .ZN(N10949) );
  AOI22D1BWP30P140LVT U9530 ( .A1(i_data_bus[723]), .A2(n6876), .B1(
        i_data_bus[691]), .B2(n6877), .ZN(n6465) );
  AOI22D1BWP30P140LVT U9531 ( .A1(i_data_bus[659]), .A2(n6878), .B1(
        i_data_bus[755]), .B2(n6879), .ZN(n6464) );
  ND2D1BWP30P140LVT U9532 ( .A1(n6465), .A2(n6464), .ZN(N10948) );
  AOI22D1BWP30P140LVT U9533 ( .A1(i_data_bus[717]), .A2(n6876), .B1(
        i_data_bus[749]), .B2(n6879), .ZN(n6467) );
  AOI22D1BWP30P140LVT U9534 ( .A1(i_data_bus[653]), .A2(n6878), .B1(
        i_data_bus[685]), .B2(n6877), .ZN(n6466) );
  ND2D1BWP30P140LVT U9535 ( .A1(n6467), .A2(n6466), .ZN(N10942) );
  AOI22D1BWP30P140LVT U9536 ( .A1(i_data_bus[748]), .A2(n6879), .B1(
        i_data_bus[684]), .B2(n6877), .ZN(n6469) );
  AOI22D1BWP30P140LVT U9537 ( .A1(i_data_bus[652]), .A2(n6878), .B1(
        i_data_bus[716]), .B2(n6876), .ZN(n6468) );
  ND2D1BWP30P140LVT U9538 ( .A1(n6469), .A2(n6468), .ZN(N10941) );
  AOI22D1BWP30P140LVT U9539 ( .A1(i_data_bus[681]), .A2(n6877), .B1(
        i_data_bus[745]), .B2(n6879), .ZN(n6471) );
  AOI22D1BWP30P140LVT U9540 ( .A1(i_data_bus[649]), .A2(n6878), .B1(
        i_data_bus[713]), .B2(n6876), .ZN(n6470) );
  ND2D1BWP30P140LVT U9541 ( .A1(n6471), .A2(n6470), .ZN(N10938) );
  AOI22D1BWP30P140LVT U9542 ( .A1(i_data_bus[675]), .A2(n6877), .B1(
        i_data_bus[739]), .B2(n6879), .ZN(n6473) );
  AOI22D1BWP30P140LVT U9543 ( .A1(i_data_bus[643]), .A2(n6878), .B1(
        i_data_bus[707]), .B2(n6876), .ZN(n6472) );
  ND2D1BWP30P140LVT U9544 ( .A1(n6473), .A2(n6472), .ZN(N10932) );
  AOI22D1BWP30P140LVT U9545 ( .A1(i_data_bus[704]), .A2(n6876), .B1(
        i_data_bus[672]), .B2(n6877), .ZN(n6475) );
  AOI22D1BWP30P140LVT U9546 ( .A1(i_data_bus[640]), .A2(n6878), .B1(
        i_data_bus[736]), .B2(n6879), .ZN(n6474) );
  ND2D1BWP30P140LVT U9547 ( .A1(n6475), .A2(n6474), .ZN(N10929) );
  AOI22D1BWP30P140LVT U9548 ( .A1(i_data_bus[703]), .A2(n6882), .B1(
        i_data_bus[735]), .B2(n6883), .ZN(n6477) );
  AOI22D1BWP30P140LVT U9549 ( .A1(i_data_bus[671]), .A2(n6884), .B1(
        i_data_bus[767]), .B2(n6885), .ZN(n6476) );
  ND2D1BWP30P140LVT U9550 ( .A1(n6477), .A2(n6476), .ZN(N8236) );
  AOI22D1BWP30P140LVT U9551 ( .A1(i_data_bus[761]), .A2(n6885), .B1(
        i_data_bus[697]), .B2(n6882), .ZN(n6479) );
  AOI22D1BWP30P140LVT U9552 ( .A1(i_data_bus[665]), .A2(n6884), .B1(
        i_data_bus[729]), .B2(n6883), .ZN(n6478) );
  ND2D1BWP30P140LVT U9553 ( .A1(n6479), .A2(n6478), .ZN(N8230) );
  AOI22D1BWP30P140LVT U9554 ( .A1(i_data_bus[758]), .A2(n6885), .B1(
        i_data_bus[726]), .B2(n6883), .ZN(n6481) );
  AOI22D1BWP30P140LVT U9555 ( .A1(i_data_bus[662]), .A2(n6884), .B1(
        i_data_bus[694]), .B2(n6882), .ZN(n6480) );
  ND2D1BWP30P140LVT U9556 ( .A1(n6481), .A2(n6480), .ZN(N8227) );
  AOI22D1BWP30P140LVT U9557 ( .A1(i_data_bus[692]), .A2(n6882), .B1(
        i_data_bus[724]), .B2(n6883), .ZN(n6483) );
  AOI22D1BWP30P140LVT U9558 ( .A1(i_data_bus[660]), .A2(n6884), .B1(
        i_data_bus[756]), .B2(n6885), .ZN(n6482) );
  ND2D1BWP30P140LVT U9559 ( .A1(n6483), .A2(n6482), .ZN(N8225) );
  AOI22D1BWP30P140LVT U9560 ( .A1(i_data_bus[685]), .A2(n6882), .B1(
        i_data_bus[717]), .B2(n6883), .ZN(n6485) );
  AOI22D1BWP30P140LVT U9561 ( .A1(i_data_bus[653]), .A2(n6884), .B1(
        i_data_bus[749]), .B2(n6885), .ZN(n6484) );
  ND2D1BWP30P140LVT U9562 ( .A1(n6485), .A2(n6484), .ZN(N8218) );
  AOI22D1BWP30P140LVT U9563 ( .A1(i_data_bus[748]), .A2(n6885), .B1(
        i_data_bus[684]), .B2(n6882), .ZN(n6487) );
  AOI22D1BWP30P140LVT U9564 ( .A1(i_data_bus[652]), .A2(n6884), .B1(
        i_data_bus[716]), .B2(n6883), .ZN(n6486) );
  ND2D1BWP30P140LVT U9565 ( .A1(n6487), .A2(n6486), .ZN(N8217) );
  AOI22D1BWP30P140LVT U9566 ( .A1(i_data_bus[746]), .A2(n6885), .B1(
        i_data_bus[714]), .B2(n6883), .ZN(n6489) );
  AOI22D1BWP30P140LVT U9567 ( .A1(i_data_bus[650]), .A2(n6884), .B1(
        i_data_bus[682]), .B2(n6882), .ZN(n6488) );
  ND2D1BWP30P140LVT U9568 ( .A1(n6489), .A2(n6488), .ZN(N8215) );
  AOI22D1BWP30P140LVT U9569 ( .A1(i_data_bus[681]), .A2(n6882), .B1(
        i_data_bus[745]), .B2(n6885), .ZN(n6491) );
  AOI22D1BWP30P140LVT U9570 ( .A1(i_data_bus[649]), .A2(n6884), .B1(
        i_data_bus[713]), .B2(n6883), .ZN(n6490) );
  ND2D1BWP30P140LVT U9571 ( .A1(n6491), .A2(n6490), .ZN(N8214) );
  AOI22D1BWP30P140LVT U9572 ( .A1(i_data_bus[675]), .A2(n6882), .B1(
        i_data_bus[707]), .B2(n6883), .ZN(n6493) );
  AOI22D1BWP30P140LVT U9573 ( .A1(i_data_bus[643]), .A2(n6884), .B1(
        i_data_bus[739]), .B2(n6885), .ZN(n6492) );
  ND2D1BWP30P140LVT U9574 ( .A1(n6493), .A2(n6492), .ZN(N8208) );
  AOI22D1BWP30P140LVT U9575 ( .A1(i_data_bus[737]), .A2(n6885), .B1(
        i_data_bus[673]), .B2(n6882), .ZN(n6495) );
  AOI22D1BWP30P140LVT U9576 ( .A1(i_data_bus[641]), .A2(n6884), .B1(
        i_data_bus[705]), .B2(n6883), .ZN(n6494) );
  ND2D1BWP30P140LVT U9577 ( .A1(n6495), .A2(n6494), .ZN(N8206) );
  AOI22D1BWP30P140LVT U9578 ( .A1(i_data_bus[764]), .A2(n6908), .B1(
        i_data_bus[700]), .B2(n6909), .ZN(n6497) );
  AOI22D1BWP30P140LVT U9579 ( .A1(i_data_bus[668]), .A2(n6910), .B1(
        i_data_bus[732]), .B2(n6911), .ZN(n6496) );
  ND2D1BWP30P140LVT U9580 ( .A1(n6497), .A2(n6496), .ZN(N5509) );
  AOI22D1BWP30P140LVT U9581 ( .A1(i_data_bus[731]), .A2(n6911), .B1(
        i_data_bus[699]), .B2(n6909), .ZN(n6499) );
  AOI22D1BWP30P140LVT U9582 ( .A1(i_data_bus[667]), .A2(n6910), .B1(
        i_data_bus[763]), .B2(n6908), .ZN(n6498) );
  ND2D1BWP30P140LVT U9583 ( .A1(n6499), .A2(n6498), .ZN(N5508) );
  AOI22D1BWP30P140LVT U9584 ( .A1(i_data_bus[761]), .A2(n6908), .B1(
        i_data_bus[697]), .B2(n6909), .ZN(n6501) );
  AOI22D1BWP30P140LVT U9585 ( .A1(i_data_bus[665]), .A2(n6910), .B1(
        i_data_bus[729]), .B2(n6911), .ZN(n6500) );
  ND2D1BWP30P140LVT U9586 ( .A1(n6501), .A2(n6500), .ZN(N5506) );
  AOI22D1BWP30P140LVT U9587 ( .A1(i_data_bus[694]), .A2(n6909), .B1(
        i_data_bus[726]), .B2(n6911), .ZN(n6503) );
  AOI22D1BWP30P140LVT U9588 ( .A1(i_data_bus[662]), .A2(n6910), .B1(
        i_data_bus[758]), .B2(n6908), .ZN(n6502) );
  ND2D1BWP30P140LVT U9589 ( .A1(n6503), .A2(n6502), .ZN(N5503) );
  AOI22D1BWP30P140LVT U9590 ( .A1(i_data_bus[692]), .A2(n6909), .B1(
        i_data_bus[724]), .B2(n6911), .ZN(n6505) );
  AOI22D1BWP30P140LVT U9591 ( .A1(i_data_bus[660]), .A2(n6910), .B1(
        i_data_bus[756]), .B2(n6908), .ZN(n6504) );
  ND2D1BWP30P140LVT U9592 ( .A1(n6505), .A2(n6504), .ZN(N5501) );
  AOI22D1BWP30P140LVT U9593 ( .A1(i_data_bus[687]), .A2(n6909), .B1(
        i_data_bus[751]), .B2(n6908), .ZN(n6507) );
  AOI22D1BWP30P140LVT U9594 ( .A1(i_data_bus[655]), .A2(n6910), .B1(
        i_data_bus[719]), .B2(n6911), .ZN(n6506) );
  ND2D1BWP30P140LVT U9595 ( .A1(n6507), .A2(n6506), .ZN(N5496) );
  AOI22D1BWP30P140LVT U9596 ( .A1(i_data_bus[686]), .A2(n6909), .B1(
        i_data_bus[750]), .B2(n6908), .ZN(n6509) );
  AOI22D1BWP30P140LVT U9597 ( .A1(i_data_bus[654]), .A2(n6910), .B1(
        i_data_bus[718]), .B2(n6911), .ZN(n6508) );
  ND2D1BWP30P140LVT U9598 ( .A1(n6509), .A2(n6508), .ZN(N5495) );
  AOI22D1BWP30P140LVT U9599 ( .A1(i_data_bus[745]), .A2(n6908), .B1(
        i_data_bus[713]), .B2(n6911), .ZN(n6511) );
  AOI22D1BWP30P140LVT U9600 ( .A1(i_data_bus[649]), .A2(n6910), .B1(
        i_data_bus[681]), .B2(n6909), .ZN(n6510) );
  ND2D1BWP30P140LVT U9601 ( .A1(n6511), .A2(n6510), .ZN(N5490) );
  AOI22D1BWP30P140LVT U9602 ( .A1(i_data_bus[675]), .A2(n6909), .B1(
        i_data_bus[739]), .B2(n6908), .ZN(n6513) );
  AOI22D1BWP30P140LVT U9603 ( .A1(i_data_bus[643]), .A2(n6910), .B1(
        i_data_bus[707]), .B2(n6911), .ZN(n6512) );
  ND2D1BWP30P140LVT U9604 ( .A1(n6513), .A2(n6512), .ZN(N5484) );
  AOI22D1BWP30P140LVT U9605 ( .A1(i_data_bus[737]), .A2(n6908), .B1(
        i_data_bus[673]), .B2(n6909), .ZN(n6515) );
  AOI22D1BWP30P140LVT U9606 ( .A1(i_data_bus[641]), .A2(n6910), .B1(
        i_data_bus[705]), .B2(n6911), .ZN(n6514) );
  ND2D1BWP30P140LVT U9607 ( .A1(n6515), .A2(n6514), .ZN(N5482) );
  AOI22D1BWP30P140LVT U9608 ( .A1(i_data_bus[699]), .A2(n6923), .B1(
        i_data_bus[763]), .B2(n6925), .ZN(n6517) );
  AOI22D1BWP30P140LVT U9609 ( .A1(i_data_bus[667]), .A2(n6924), .B1(
        i_data_bus[731]), .B2(n6922), .ZN(n6516) );
  ND2D1BWP30P140LVT U9610 ( .A1(n6517), .A2(n6516), .ZN(N9850) );
  AOI22D1BWP30P140LVT U9611 ( .A1(i_data_bus[761]), .A2(n6925), .B1(
        i_data_bus[697]), .B2(n6923), .ZN(n6519) );
  AOI22D1BWP30P140LVT U9612 ( .A1(i_data_bus[665]), .A2(n6924), .B1(
        i_data_bus[729]), .B2(n6922), .ZN(n6518) );
  ND2D1BWP30P140LVT U9613 ( .A1(n6519), .A2(n6518), .ZN(N9848) );
  AOI22D1BWP30P140LVT U9614 ( .A1(i_data_bus[728]), .A2(n6922), .B1(
        i_data_bus[696]), .B2(n6923), .ZN(n6521) );
  AOI22D1BWP30P140LVT U9615 ( .A1(i_data_bus[664]), .A2(n6924), .B1(
        i_data_bus[760]), .B2(n6925), .ZN(n6520) );
  ND2D1BWP30P140LVT U9616 ( .A1(n6521), .A2(n6520), .ZN(N9847) );
  AOI22D1BWP30P140LVT U9617 ( .A1(i_data_bus[694]), .A2(n6923), .B1(
        i_data_bus[758]), .B2(n6925), .ZN(n6523) );
  AOI22D1BWP30P140LVT U9618 ( .A1(i_data_bus[662]), .A2(n6924), .B1(
        i_data_bus[726]), .B2(n6922), .ZN(n6522) );
  ND2D1BWP30P140LVT U9619 ( .A1(n6523), .A2(n6522), .ZN(N9845) );
  AOI22D1BWP30P140LVT U9620 ( .A1(i_data_bus[719]), .A2(n6922), .B1(
        i_data_bus[751]), .B2(n6925), .ZN(n6525) );
  AOI22D1BWP30P140LVT U9621 ( .A1(i_data_bus[655]), .A2(n6924), .B1(
        i_data_bus[687]), .B2(n6923), .ZN(n6524) );
  ND2D1BWP30P140LVT U9622 ( .A1(n6525), .A2(n6524), .ZN(N9838) );
  AOI22D1BWP30P140LVT U9623 ( .A1(i_data_bus[750]), .A2(n6925), .B1(
        i_data_bus[718]), .B2(n6922), .ZN(n6527) );
  AOI22D1BWP30P140LVT U9624 ( .A1(i_data_bus[654]), .A2(n6924), .B1(
        i_data_bus[686]), .B2(n6923), .ZN(n6526) );
  ND2D1BWP30P140LVT U9625 ( .A1(n6527), .A2(n6526), .ZN(N9837) );
  AOI22D1BWP30P140LVT U9626 ( .A1(i_data_bus[745]), .A2(n6925), .B1(
        i_data_bus[713]), .B2(n6922), .ZN(n6529) );
  AOI22D1BWP30P140LVT U9627 ( .A1(i_data_bus[649]), .A2(n6924), .B1(
        i_data_bus[681]), .B2(n6923), .ZN(n6528) );
  ND2D1BWP30P140LVT U9628 ( .A1(n6529), .A2(n6528), .ZN(N9832) );
  AOI22D1BWP30P140LVT U9629 ( .A1(i_data_bus[675]), .A2(n6923), .B1(
        i_data_bus[739]), .B2(n6925), .ZN(n6531) );
  AOI22D1BWP30P140LVT U9630 ( .A1(i_data_bus[643]), .A2(n6924), .B1(
        i_data_bus[707]), .B2(n6922), .ZN(n6530) );
  ND2D1BWP30P140LVT U9631 ( .A1(n6531), .A2(n6530), .ZN(N9826) );
  AOI22D1BWP30P140LVT U9632 ( .A1(i_data_bus[737]), .A2(n6925), .B1(
        i_data_bus[673]), .B2(n6923), .ZN(n6533) );
  AOI22D1BWP30P140LVT U9633 ( .A1(i_data_bus[641]), .A2(n6924), .B1(
        i_data_bus[705]), .B2(n6922), .ZN(n6532) );
  ND2D1BWP30P140LVT U9634 ( .A1(n6533), .A2(n6532), .ZN(N9824) );
  AOI22D1BWP30P140LVT U9635 ( .A1(i_data_bus[846]), .A2(n6722), .B1(
        i_data_bus[782]), .B2(n6720), .ZN(n6535) );
  AOI22D1BWP30P140LVT U9636 ( .A1(i_data_bus[814]), .A2(n6721), .B1(
        i_data_bus[878]), .B2(n6723), .ZN(n6534) );
  ND2D1BWP30P140LVT U9637 ( .A1(n6535), .A2(n6534), .ZN(N5583) );
  AOI22D1BWP30P140LVT U9638 ( .A1(i_data_bus[813]), .A2(n6721), .B1(
        i_data_bus[781]), .B2(n6720), .ZN(n6537) );
  AOI22D1BWP30P140LVT U9639 ( .A1(i_data_bus[845]), .A2(n6722), .B1(
        i_data_bus[877]), .B2(n6723), .ZN(n6536) );
  ND2D1BWP30P140LVT U9640 ( .A1(n6537), .A2(n6536), .ZN(N5582) );
  AOI22D1BWP30P140LVT U9641 ( .A1(i_data_bus[703]), .A2(n6620), .B1(
        i_data_bus[671]), .B2(n6225), .ZN(n6539) );
  AOI22D1BWP30P140LVT U9642 ( .A1(i_data_bus[735]), .A2(n6619), .B1(
        i_data_bus[767]), .B2(n6618), .ZN(n6538) );
  ND2D1BWP30P140LVT U9643 ( .A1(n6539), .A2(n6538), .ZN(N4406) );
  AOI22D1BWP30P140LVT U9644 ( .A1(i_data_bus[698]), .A2(n6620), .B1(
        i_data_bus[666]), .B2(n6225), .ZN(n6541) );
  AOI22D1BWP30P140LVT U9645 ( .A1(i_data_bus[730]), .A2(n6619), .B1(
        i_data_bus[762]), .B2(n6618), .ZN(n6540) );
  ND2D1BWP30P140LVT U9646 ( .A1(n6541), .A2(n6540), .ZN(N4401) );
  AOI22D1BWP30P140LVT U9647 ( .A1(i_data_bus[688]), .A2(n6620), .B1(
        i_data_bus[656]), .B2(n6225), .ZN(n6543) );
  AOI22D1BWP30P140LVT U9648 ( .A1(i_data_bus[720]), .A2(n6619), .B1(
        i_data_bus[752]), .B2(n6618), .ZN(n6542) );
  ND2D1BWP30P140LVT U9649 ( .A1(n6543), .A2(n6542), .ZN(N4391) );
  AOI22D1BWP30P140LVT U9650 ( .A1(i_data_bus[687]), .A2(n6620), .B1(
        i_data_bus[719]), .B2(n6619), .ZN(n6545) );
  AOI22D1BWP30P140LVT U9651 ( .A1(i_data_bus[655]), .A2(n6225), .B1(
        i_data_bus[751]), .B2(n6618), .ZN(n6544) );
  ND2D1BWP30P140LVT U9652 ( .A1(n6545), .A2(n6544), .ZN(N4390) );
  AOI22D1BWP30P140LVT U9653 ( .A1(i_data_bus[654]), .A2(n6225), .B1(
        i_data_bus[718]), .B2(n6619), .ZN(n6547) );
  AOI22D1BWP30P140LVT U9654 ( .A1(i_data_bus[686]), .A2(n6620), .B1(
        i_data_bus[750]), .B2(n6618), .ZN(n6546) );
  ND2D1BWP30P140LVT U9655 ( .A1(n6547), .A2(n6546), .ZN(N4389) );
  AOI22D1BWP30P140LVT U9656 ( .A1(i_data_bus[664]), .A2(n6942), .B1(
        i_data_bus[696]), .B2(n6943), .ZN(n6553) );
  AOI22D1BWP30P140LVT U9657 ( .A1(i_data_bus[728]), .A2(n6941), .B1(
        i_data_bus[760]), .B2(n6940), .ZN(n6552) );
  ND2D1BWP30P140LVT U9658 ( .A1(n6553), .A2(n6552), .ZN(N2781) );
  AOI22D1BWP30P140LVT U9659 ( .A1(i_data_bus[662]), .A2(n6942), .B1(
        i_data_bus[726]), .B2(n6941), .ZN(n6555) );
  AOI22D1BWP30P140LVT U9660 ( .A1(i_data_bus[694]), .A2(n6943), .B1(
        i_data_bus[758]), .B2(n6940), .ZN(n6554) );
  ND2D1BWP30P140LVT U9661 ( .A1(n6555), .A2(n6554), .ZN(N2779) );
  AOI22D1BWP30P140LVT U9662 ( .A1(i_data_bus[655]), .A2(n6942), .B1(
        i_data_bus[719]), .B2(n6941), .ZN(n6557) );
  AOI22D1BWP30P140LVT U9663 ( .A1(i_data_bus[687]), .A2(n6943), .B1(
        i_data_bus[751]), .B2(n6940), .ZN(n6556) );
  ND2D1BWP30P140LVT U9664 ( .A1(n6557), .A2(n6556), .ZN(N2772) );
  AOI22D1BWP30P140LVT U9665 ( .A1(i_data_bus[654]), .A2(n6942), .B1(
        i_data_bus[718]), .B2(n6941), .ZN(n6559) );
  AOI22D1BWP30P140LVT U9666 ( .A1(i_data_bus[686]), .A2(n6943), .B1(
        i_data_bus[750]), .B2(n6940), .ZN(n6558) );
  ND2D1BWP30P140LVT U9667 ( .A1(n6559), .A2(n6558), .ZN(N2771) );
  AOI22D1BWP30P140LVT U9668 ( .A1(i_data_bus[653]), .A2(n6942), .B1(
        i_data_bus[685]), .B2(n6943), .ZN(n6561) );
  AOI22D1BWP30P140LVT U9669 ( .A1(i_data_bus[717]), .A2(n6941), .B1(
        i_data_bus[749]), .B2(n6940), .ZN(n6560) );
  ND2D1BWP30P140LVT U9670 ( .A1(n6561), .A2(n6560), .ZN(N2770) );
  AOI22D1BWP30P140LVT U9671 ( .A1(i_data_bus[668]), .A2(n6225), .B1(
        i_data_bus[764]), .B2(n6618), .ZN(n6563) );
  AOI22D1BWP30P140LVT U9672 ( .A1(i_data_bus[732]), .A2(n6619), .B1(
        i_data_bus[700]), .B2(n6620), .ZN(n6562) );
  ND2D1BWP30P140LVT U9673 ( .A1(n6563), .A2(n6562), .ZN(N4403) );
  AOI22D1BWP30P140LVT U9674 ( .A1(i_data_bus[759]), .A2(n6618), .B1(
        i_data_bus[727]), .B2(n6619), .ZN(n6565) );
  AOI22D1BWP30P140LVT U9675 ( .A1(i_data_bus[663]), .A2(n6225), .B1(
        i_data_bus[695]), .B2(n6620), .ZN(n6564) );
  ND2D1BWP30P140LVT U9676 ( .A1(n6565), .A2(n6564), .ZN(N4398) );
  AOI22D1BWP30P140LVT U9677 ( .A1(i_data_bus[758]), .A2(n6618), .B1(
        i_data_bus[726]), .B2(n6619), .ZN(n6567) );
  AOI22D1BWP30P140LVT U9678 ( .A1(i_data_bus[662]), .A2(n6225), .B1(
        i_data_bus[694]), .B2(n6620), .ZN(n6566) );
  ND2D1BWP30P140LVT U9679 ( .A1(n6567), .A2(n6566), .ZN(N4397) );
  AOI22D1BWP30P140LVT U9680 ( .A1(i_data_bus[754]), .A2(n6618), .B1(
        i_data_bus[658]), .B2(n6225), .ZN(n6569) );
  AOI22D1BWP30P140LVT U9681 ( .A1(i_data_bus[722]), .A2(n6619), .B1(
        i_data_bus[690]), .B2(n6620), .ZN(n6568) );
  ND2D1BWP30P140LVT U9682 ( .A1(n6569), .A2(n6568), .ZN(N4393) );
  AOI22D1BWP30P140LVT U9683 ( .A1(i_data_bus[715]), .A2(n6619), .B1(
        i_data_bus[651]), .B2(n6225), .ZN(n6571) );
  AOI22D1BWP30P140LVT U9684 ( .A1(i_data_bus[747]), .A2(n6618), .B1(
        i_data_bus[683]), .B2(n6620), .ZN(n6570) );
  ND2D1BWP30P140LVT U9685 ( .A1(n6571), .A2(n6570), .ZN(N4386) );
  AOI22D1BWP30P140LVT U9686 ( .A1(i_data_bus[711]), .A2(n6619), .B1(
        i_data_bus[647]), .B2(n6225), .ZN(n6573) );
  AOI22D1BWP30P140LVT U9687 ( .A1(i_data_bus[743]), .A2(n6618), .B1(
        i_data_bus[679]), .B2(n6620), .ZN(n6572) );
  ND2D1BWP30P140LVT U9688 ( .A1(n6573), .A2(n6572), .ZN(N4382) );
  AOI22D1BWP30P140LVT U9689 ( .A1(i_data_bus[640]), .A2(n6225), .B1(
        i_data_bus[736]), .B2(n6618), .ZN(n6575) );
  AOI22D1BWP30P140LVT U9690 ( .A1(i_data_bus[704]), .A2(n6619), .B1(
        i_data_bus[672]), .B2(n6620), .ZN(n6574) );
  ND2D1BWP30P140LVT U9691 ( .A1(n6575), .A2(n6574), .ZN(N4375) );
  AOI22D1BWP30P140LVT U9692 ( .A1(i_data_bus[663]), .A2(n6942), .B1(
        i_data_bus[727]), .B2(n6941), .ZN(n6577) );
  AOI22D1BWP30P140LVT U9693 ( .A1(i_data_bus[759]), .A2(n6940), .B1(
        i_data_bus[695]), .B2(n6943), .ZN(n6576) );
  ND2D1BWP30P140LVT U9694 ( .A1(n6577), .A2(n6576), .ZN(N2780) );
  AOI22D1BWP30P140LVT U9695 ( .A1(i_data_bus[652]), .A2(n6942), .B1(
        i_data_bus[716]), .B2(n6941), .ZN(n6579) );
  AOI22D1BWP30P140LVT U9696 ( .A1(i_data_bus[748]), .A2(n6940), .B1(
        i_data_bus[684]), .B2(n6943), .ZN(n6578) );
  ND2D1BWP30P140LVT U9697 ( .A1(n6579), .A2(n6578), .ZN(N2769) );
  AOI22D1BWP30P140LVT U9698 ( .A1(i_data_bus[746]), .A2(n6940), .B1(
        i_data_bus[714]), .B2(n6941), .ZN(n6581) );
  AOI22D1BWP30P140LVT U9699 ( .A1(i_data_bus[650]), .A2(n6942), .B1(
        i_data_bus[682]), .B2(n6943), .ZN(n6580) );
  ND2D1BWP30P140LVT U9700 ( .A1(n6581), .A2(n6580), .ZN(N2767) );
  AOI22D1BWP30P140LVT U9701 ( .A1(i_data_bus[745]), .A2(n6940), .B1(
        i_data_bus[713]), .B2(n6941), .ZN(n6583) );
  AOI22D1BWP30P140LVT U9702 ( .A1(i_data_bus[649]), .A2(n6942), .B1(
        i_data_bus[681]), .B2(n6943), .ZN(n6582) );
  ND2D1BWP30P140LVT U9703 ( .A1(n6583), .A2(n6582), .ZN(N2766) );
  AOI22D1BWP30P140LVT U9704 ( .A1(i_data_bus[641]), .A2(n6942), .B1(
        i_data_bus[705]), .B2(n6941), .ZN(n6585) );
  AOI22D1BWP30P140LVT U9705 ( .A1(i_data_bus[737]), .A2(n6940), .B1(
        i_data_bus[673]), .B2(n6943), .ZN(n6584) );
  ND2D1BWP30P140LVT U9706 ( .A1(n6585), .A2(n6584), .ZN(N2758) );
  AOI22D1BWP30P140LVT U9707 ( .A1(i_data_bus[670]), .A2(n6942), .B1(
        i_data_bus[702]), .B2(n6943), .ZN(n6587) );
  AOI22D1BWP30P140LVT U9708 ( .A1(i_data_bus[766]), .A2(n6940), .B1(
        i_data_bus[734]), .B2(n6941), .ZN(n6586) );
  ND2D1BWP30P140LVT U9709 ( .A1(n6587), .A2(n6586), .ZN(N2787) );
  AOI22D1BWP30P140LVT U9710 ( .A1(i_data_bus[764]), .A2(n6940), .B1(
        i_data_bus[700]), .B2(n6943), .ZN(n6589) );
  AOI22D1BWP30P140LVT U9711 ( .A1(i_data_bus[668]), .A2(n6942), .B1(
        i_data_bus[732]), .B2(n6941), .ZN(n6588) );
  ND2D1BWP30P140LVT U9712 ( .A1(n6589), .A2(n6588), .ZN(N2785) );
  AOI22D1BWP30P140LVT U9713 ( .A1(i_data_bus[699]), .A2(n6943), .B1(
        i_data_bus[763]), .B2(n6940), .ZN(n6591) );
  AOI22D1BWP30P140LVT U9714 ( .A1(i_data_bus[667]), .A2(n6942), .B1(
        i_data_bus[731]), .B2(n6941), .ZN(n6590) );
  ND2D1BWP30P140LVT U9715 ( .A1(n6591), .A2(n6590), .ZN(N2784) );
  AOI22D1BWP30P140LVT U9716 ( .A1(i_data_bus[755]), .A2(n6940), .B1(
        i_data_bus[691]), .B2(n6943), .ZN(n6593) );
  AOI22D1BWP30P140LVT U9717 ( .A1(i_data_bus[659]), .A2(n6942), .B1(
        i_data_bus[723]), .B2(n6941), .ZN(n6592) );
  ND2D1BWP30P140LVT U9718 ( .A1(n6593), .A2(n6592), .ZN(N2776) );
  AOI22D1BWP30P140LVT U9719 ( .A1(i_data_bus[643]), .A2(n6942), .B1(
        i_data_bus[739]), .B2(n6940), .ZN(n6595) );
  AOI22D1BWP30P140LVT U9720 ( .A1(i_data_bus[675]), .A2(n6943), .B1(
        i_data_bus[707]), .B2(n6941), .ZN(n6594) );
  ND2D1BWP30P140LVT U9721 ( .A1(n6595), .A2(n6594), .ZN(N2760) );
  AOI22D1BWP30P140LVT U9722 ( .A1(i_data_bus[699]), .A2(n6620), .B1(
        i_data_bus[763]), .B2(n6618), .ZN(n6597) );
  AOI22D1BWP30P140LVT U9723 ( .A1(i_data_bus[667]), .A2(n6225), .B1(
        i_data_bus[731]), .B2(n6619), .ZN(n6596) );
  ND2D1BWP30P140LVT U9724 ( .A1(n6597), .A2(n6596), .ZN(N4402) );
  AOI22D1BWP30P140LVT U9725 ( .A1(i_data_bus[760]), .A2(n6618), .B1(
        i_data_bus[696]), .B2(n6620), .ZN(n6599) );
  AOI22D1BWP30P140LVT U9726 ( .A1(i_data_bus[664]), .A2(n6225), .B1(
        i_data_bus[728]), .B2(n6619), .ZN(n6598) );
  ND2D1BWP30P140LVT U9727 ( .A1(n6599), .A2(n6598), .ZN(N4399) );
  AOI22D1BWP30P140LVT U9728 ( .A1(i_data_bus[660]), .A2(n6225), .B1(
        i_data_bus[756]), .B2(n6618), .ZN(n6601) );
  AOI22D1BWP30P140LVT U9729 ( .A1(i_data_bus[692]), .A2(n6620), .B1(
        i_data_bus[724]), .B2(n6619), .ZN(n6600) );
  ND2D1BWP30P140LVT U9730 ( .A1(n6601), .A2(n6600), .ZN(N4395) );
  AOI22D1BWP30P140LVT U9731 ( .A1(i_data_bus[659]), .A2(n6225), .B1(
        i_data_bus[691]), .B2(n6620), .ZN(n6603) );
  AOI22D1BWP30P140LVT U9732 ( .A1(i_data_bus[755]), .A2(n6618), .B1(
        i_data_bus[723]), .B2(n6619), .ZN(n6602) );
  ND2D1BWP30P140LVT U9733 ( .A1(n6603), .A2(n6602), .ZN(N4394) );
  AOI22D1BWP30P140LVT U9734 ( .A1(i_data_bus[685]), .A2(n6620), .B1(
        i_data_bus[749]), .B2(n6618), .ZN(n6605) );
  AOI22D1BWP30P140LVT U9735 ( .A1(i_data_bus[653]), .A2(n6225), .B1(
        i_data_bus[717]), .B2(n6619), .ZN(n6604) );
  ND2D1BWP30P140LVT U9736 ( .A1(n6605), .A2(n6604), .ZN(N4388) );
  AOI22D1BWP30P140LVT U9737 ( .A1(i_data_bus[748]), .A2(n6618), .B1(
        i_data_bus[684]), .B2(n6620), .ZN(n6607) );
  AOI22D1BWP30P140LVT U9738 ( .A1(i_data_bus[652]), .A2(n6225), .B1(
        i_data_bus[716]), .B2(n6619), .ZN(n6606) );
  ND2D1BWP30P140LVT U9739 ( .A1(n6607), .A2(n6606), .ZN(N4387) );
  AOI22D1BWP30P140LVT U9740 ( .A1(i_data_bus[650]), .A2(n6225), .B1(
        i_data_bus[682]), .B2(n6620), .ZN(n6609) );
  AOI22D1BWP30P140LVT U9741 ( .A1(i_data_bus[746]), .A2(n6618), .B1(
        i_data_bus[714]), .B2(n6619), .ZN(n6608) );
  ND2D1BWP30P140LVT U9742 ( .A1(n6609), .A2(n6608), .ZN(N4385) );
  AOI22D1BWP30P140LVT U9743 ( .A1(i_data_bus[649]), .A2(n6225), .B1(
        i_data_bus[681]), .B2(n6620), .ZN(n6611) );
  AOI22D1BWP30P140LVT U9744 ( .A1(i_data_bus[745]), .A2(n6618), .B1(
        i_data_bus[713]), .B2(n6619), .ZN(n6610) );
  ND2D1BWP30P140LVT U9745 ( .A1(n6611), .A2(n6610), .ZN(N4384) );
  AOI22D1BWP30P140LVT U9746 ( .A1(i_data_bus[680]), .A2(n6620), .B1(
        i_data_bus[648]), .B2(n6225), .ZN(n6613) );
  AOI22D1BWP30P140LVT U9747 ( .A1(i_data_bus[744]), .A2(n6618), .B1(
        i_data_bus[712]), .B2(n6619), .ZN(n6612) );
  ND2D1BWP30P140LVT U9748 ( .A1(n6613), .A2(n6612), .ZN(N4383) );
  AOI22D1BWP30P140LVT U9749 ( .A1(i_data_bus[742]), .A2(n6618), .B1(
        i_data_bus[646]), .B2(n6225), .ZN(n6615) );
  AOI22D1BWP30P140LVT U9750 ( .A1(i_data_bus[678]), .A2(n6620), .B1(
        i_data_bus[710]), .B2(n6619), .ZN(n6614) );
  ND2D1BWP30P140LVT U9751 ( .A1(n6615), .A2(n6614), .ZN(N4381) );
  AOI22D1BWP30P140LVT U9752 ( .A1(i_data_bus[675]), .A2(n6620), .B1(
        i_data_bus[739]), .B2(n6618), .ZN(n6617) );
  AOI22D1BWP30P140LVT U9753 ( .A1(i_data_bus[643]), .A2(n6225), .B1(
        i_data_bus[707]), .B2(n6619), .ZN(n6616) );
  ND2D1BWP30P140LVT U9754 ( .A1(n6617), .A2(n6616), .ZN(N4378) );
  AOI22D1BWP30P140LVT U9755 ( .A1(i_data_bus[738]), .A2(n6618), .B1(
        i_data_bus[642]), .B2(n6225), .ZN(n6622) );
  AOI22D1BWP30P140LVT U9756 ( .A1(i_data_bus[674]), .A2(n6620), .B1(
        i_data_bus[706]), .B2(n6619), .ZN(n6621) );
  ND2D1BWP30P140LVT U9757 ( .A1(n6622), .A2(n6621), .ZN(N4377) );
  AOI22D1BWP30P140LVT U9758 ( .A1(i_data_bus[886]), .A2(n6723), .B1(
        i_data_bus[822]), .B2(n6721), .ZN(n6624) );
  AOI22D1BWP30P140LVT U9759 ( .A1(i_data_bus[854]), .A2(n6722), .B1(
        i_data_bus[790]), .B2(n6720), .ZN(n6623) );
  ND2D1BWP30P140LVT U9760 ( .A1(n6624), .A2(n6623), .ZN(N5591) );
  AOI22D1BWP30P140LVT U9761 ( .A1(i_data_bus[789]), .A2(n6720), .B1(
        i_data_bus[821]), .B2(n6721), .ZN(n6626) );
  AOI22D1BWP30P140LVT U9762 ( .A1(i_data_bus[853]), .A2(n6722), .B1(
        i_data_bus[885]), .B2(n6723), .ZN(n6625) );
  ND2D1BWP30P140LVT U9763 ( .A1(n6626), .A2(n6625), .ZN(N5590) );
  AOI22D1BWP30P140LVT U9764 ( .A1(i_data_bus[840]), .A2(n6722), .B1(
        i_data_bus[808]), .B2(n6721), .ZN(n6628) );
  AOI22D1BWP30P140LVT U9765 ( .A1(i_data_bus[776]), .A2(n6720), .B1(
        i_data_bus[872]), .B2(n6723), .ZN(n6627) );
  ND2D1BWP30P140LVT U9766 ( .A1(n6628), .A2(n6627), .ZN(N5577) );
  AOI22D1BWP30P140LVT U9767 ( .A1(i_data_bus[834]), .A2(n6722), .B1(
        i_data_bus[802]), .B2(n6721), .ZN(n6630) );
  AOI22D1BWP30P140LVT U9768 ( .A1(i_data_bus[770]), .A2(n6720), .B1(
        i_data_bus[866]), .B2(n6723), .ZN(n6629) );
  ND2D1BWP30P140LVT U9769 ( .A1(n6630), .A2(n6629), .ZN(N5571) );
  AOI22D1BWP30P140LVT U9770 ( .A1(i_data_bus[832]), .A2(n6722), .B1(
        i_data_bus[800]), .B2(n6721), .ZN(n6632) );
  AOI22D1BWP30P140LVT U9771 ( .A1(i_data_bus[768]), .A2(n6720), .B1(
        i_data_bus[864]), .B2(n6723), .ZN(n6631) );
  ND2D1BWP30P140LVT U9772 ( .A1(n6632), .A2(n6631), .ZN(N5569) );
  AOI22D1BWP30P140LVT U9773 ( .A1(i_data_bus[817]), .A2(n6721), .B1(
        i_data_bus[849]), .B2(n6722), .ZN(n6634) );
  AOI22D1BWP30P140LVT U9774 ( .A1(i_data_bus[881]), .A2(n6723), .B1(
        i_data_bus[785]), .B2(n6720), .ZN(n6633) );
  ND2D1BWP30P140LVT U9775 ( .A1(n6634), .A2(n6633), .ZN(N5586) );
  AOI22D1BWP30P140LVT U9776 ( .A1(i_data_bus[880]), .A2(n6723), .B1(
        i_data_bus[848]), .B2(n6722), .ZN(n6636) );
  AOI22D1BWP30P140LVT U9777 ( .A1(i_data_bus[816]), .A2(n6721), .B1(
        i_data_bus[784]), .B2(n6720), .ZN(n6635) );
  ND2D1BWP30P140LVT U9778 ( .A1(n6636), .A2(n6635), .ZN(N5585) );
  AOI22D1BWP30P140LVT U9779 ( .A1(i_data_bus[870]), .A2(n6723), .B1(
        i_data_bus[838]), .B2(n6722), .ZN(n6638) );
  AOI22D1BWP30P140LVT U9780 ( .A1(i_data_bus[806]), .A2(n6721), .B1(
        i_data_bus[774]), .B2(n6720), .ZN(n6637) );
  ND2D1BWP30P140LVT U9781 ( .A1(n6638), .A2(n6637), .ZN(N5575) );
  AOI22D1BWP30P140LVT U9782 ( .A1(i_data_bus[810]), .A2(n6721), .B1(
        i_data_bus[842]), .B2(n6722), .ZN(n6640) );
  AOI22D1BWP30P140LVT U9783 ( .A1(i_data_bus[778]), .A2(n6720), .B1(
        i_data_bus[874]), .B2(n6723), .ZN(n6639) );
  ND2D1BWP30P140LVT U9784 ( .A1(n6640), .A2(n6639), .ZN(N5579) );
  AOI22D1BWP30P140LVT U9785 ( .A1(i_data_bus[803]), .A2(n6721), .B1(
        i_data_bus[835]), .B2(n6722), .ZN(n6642) );
  AOI22D1BWP30P140LVT U9786 ( .A1(i_data_bus[771]), .A2(n6720), .B1(
        i_data_bus[867]), .B2(n6723), .ZN(n6641) );
  ND2D1BWP30P140LVT U9787 ( .A1(n6642), .A2(n6641), .ZN(N5572) );
  AOI22D1BWP30P140LVT U9788 ( .A1(i_data_bus[841]), .A2(n6760), .B1(
        i_data_bus[809]), .B2(n6759), .ZN(n6644) );
  AOI22D1BWP30P140LVT U9789 ( .A1(i_data_bus[873]), .A2(n6761), .B1(
        i_data_bus[777]), .B2(n6758), .ZN(n6643) );
  ND2D1BWP30P140LVT U9790 ( .A1(n6644), .A2(n6643), .ZN(N7324) );
  AOI22D1BWP30P140LVT U9791 ( .A1(i_data_bus[779]), .A2(n6758), .B1(
        i_data_bus[811]), .B2(n6759), .ZN(n6646) );
  AOI22D1BWP30P140LVT U9792 ( .A1(i_data_bus[843]), .A2(n6760), .B1(
        i_data_bus[875]), .B2(n6761), .ZN(n6645) );
  ND2D1BWP30P140LVT U9793 ( .A1(n6646), .A2(n6645), .ZN(N7326) );
  AOI22D1BWP30P140LVT U9794 ( .A1(i_data_bus[834]), .A2(n6760), .B1(
        i_data_bus[802]), .B2(n6759), .ZN(n6648) );
  AOI22D1BWP30P140LVT U9795 ( .A1(i_data_bus[770]), .A2(n6758), .B1(
        i_data_bus[866]), .B2(n6761), .ZN(n6647) );
  ND2D1BWP30P140LVT U9796 ( .A1(n6648), .A2(n6647), .ZN(N7317) );
  AOI22D1BWP30P140LVT U9797 ( .A1(i_data_bus[832]), .A2(n6760), .B1(
        i_data_bus[800]), .B2(n6759), .ZN(n6650) );
  AOI22D1BWP30P140LVT U9798 ( .A1(i_data_bus[768]), .A2(n6758), .B1(
        i_data_bus[864]), .B2(n6761), .ZN(n6649) );
  ND2D1BWP30P140LVT U9799 ( .A1(n6650), .A2(n6649), .ZN(N7315) );
  AOI22D1BWP30P140LVT U9800 ( .A1(i_data_bus[830]), .A2(n6759), .B1(
        i_data_bus[862]), .B2(n6760), .ZN(n6652) );
  AOI22D1BWP30P140LVT U9801 ( .A1(i_data_bus[894]), .A2(n6761), .B1(
        i_data_bus[798]), .B2(n6758), .ZN(n6651) );
  ND2D1BWP30P140LVT U9802 ( .A1(n6652), .A2(n6651), .ZN(N7345) );
  AOI22D1BWP30P140LVT U9803 ( .A1(i_data_bus[814]), .A2(n6759), .B1(
        i_data_bus[846]), .B2(n6760), .ZN(n6654) );
  AOI22D1BWP30P140LVT U9804 ( .A1(i_data_bus[878]), .A2(n6761), .B1(
        i_data_bus[782]), .B2(n6758), .ZN(n6653) );
  ND2D1BWP30P140LVT U9805 ( .A1(n6654), .A2(n6653), .ZN(N7329) );
  AOI22D1BWP30P140LVT U9806 ( .A1(i_data_bus[806]), .A2(n6759), .B1(
        i_data_bus[838]), .B2(n6760), .ZN(n6656) );
  AOI22D1BWP30P140LVT U9807 ( .A1(i_data_bus[870]), .A2(n6761), .B1(
        i_data_bus[774]), .B2(n6758), .ZN(n6655) );
  ND2D1BWP30P140LVT U9808 ( .A1(n6656), .A2(n6655), .ZN(N7321) );
  AOI22D1BWP30P140LVT U9809 ( .A1(i_data_bus[880]), .A2(n6761), .B1(
        i_data_bus[848]), .B2(n6760), .ZN(n6658) );
  AOI22D1BWP30P140LVT U9810 ( .A1(i_data_bus[816]), .A2(n6759), .B1(
        i_data_bus[784]), .B2(n6758), .ZN(n6657) );
  ND2D1BWP30P140LVT U9811 ( .A1(n6658), .A2(n6657), .ZN(N7331) );
  AOI22D1BWP30P140LVT U9812 ( .A1(i_data_bus[825]), .A2(n6759), .B1(
        i_data_bus[857]), .B2(n6760), .ZN(n6660) );
  AOI22D1BWP30P140LVT U9813 ( .A1(i_data_bus[793]), .A2(n6758), .B1(
        i_data_bus[889]), .B2(n6761), .ZN(n6659) );
  ND2D1BWP30P140LVT U9814 ( .A1(n6660), .A2(n6659), .ZN(N7340) );
  AOI22D1BWP30P140LVT U9815 ( .A1(i_data_bus[786]), .A2(n6758), .B1(
        i_data_bus[850]), .B2(n6760), .ZN(n6662) );
  AOI22D1BWP30P140LVT U9816 ( .A1(i_data_bus[818]), .A2(n6759), .B1(
        i_data_bus[882]), .B2(n6761), .ZN(n6661) );
  ND2D1BWP30P140LVT U9817 ( .A1(n6662), .A2(n6661), .ZN(N7333) );
  AOI22D1BWP30P140LVT U9818 ( .A1(i_data_bus[771]), .A2(n6758), .B1(
        i_data_bus[835]), .B2(n6760), .ZN(n6664) );
  AOI22D1BWP30P140LVT U9819 ( .A1(i_data_bus[803]), .A2(n6759), .B1(
        i_data_bus[867]), .B2(n6761), .ZN(n6663) );
  ND2D1BWP30P140LVT U9820 ( .A1(n6664), .A2(n6663), .ZN(N7318) );
  AOI22D1BWP30P140LVT U9821 ( .A1(i_data_bus[799]), .A2(n6720), .B1(
        i_data_bus[863]), .B2(n6722), .ZN(n6666) );
  AOI22D1BWP30P140LVT U9822 ( .A1(i_data_bus[895]), .A2(n6723), .B1(
        i_data_bus[831]), .B2(n6721), .ZN(n6665) );
  ND2D1BWP30P140LVT U9823 ( .A1(n6666), .A2(n6665), .ZN(N5600) );
  AOI22D1BWP30P140LVT U9824 ( .A1(i_data_bus[798]), .A2(n6720), .B1(
        i_data_bus[862]), .B2(n6722), .ZN(n6668) );
  AOI22D1BWP30P140LVT U9825 ( .A1(i_data_bus[894]), .A2(n6723), .B1(
        i_data_bus[830]), .B2(n6721), .ZN(n6667) );
  ND2D1BWP30P140LVT U9826 ( .A1(n6668), .A2(n6667), .ZN(N5599) );
  AOI22D1BWP30P140LVT U9827 ( .A1(i_data_bus[860]), .A2(n6722), .B1(
        i_data_bus[796]), .B2(n6720), .ZN(n6670) );
  AOI22D1BWP30P140LVT U9828 ( .A1(i_data_bus[892]), .A2(n6723), .B1(
        i_data_bus[828]), .B2(n6721), .ZN(n6669) );
  ND2D1BWP30P140LVT U9829 ( .A1(n6670), .A2(n6669), .ZN(N5597) );
  AOI22D1BWP30P140LVT U9830 ( .A1(i_data_bus[891]), .A2(n6723), .B1(
        i_data_bus[859]), .B2(n6722), .ZN(n6672) );
  AOI22D1BWP30P140LVT U9831 ( .A1(i_data_bus[795]), .A2(n6720), .B1(
        i_data_bus[827]), .B2(n6721), .ZN(n6671) );
  ND2D1BWP30P140LVT U9832 ( .A1(n6672), .A2(n6671), .ZN(N5596) );
  AOI22D1BWP30P140LVT U9833 ( .A1(i_data_bus[858]), .A2(n6722), .B1(
        i_data_bus[890]), .B2(n6723), .ZN(n6674) );
  AOI22D1BWP30P140LVT U9834 ( .A1(i_data_bus[794]), .A2(n6720), .B1(
        i_data_bus[826]), .B2(n6721), .ZN(n6673) );
  ND2D1BWP30P140LVT U9835 ( .A1(n6674), .A2(n6673), .ZN(N5595) );
  AOI22D1BWP30P140LVT U9836 ( .A1(i_data_bus[889]), .A2(n6723), .B1(
        i_data_bus[857]), .B2(n6722), .ZN(n6676) );
  AOI22D1BWP30P140LVT U9837 ( .A1(i_data_bus[793]), .A2(n6720), .B1(
        i_data_bus[825]), .B2(n6721), .ZN(n6675) );
  ND2D1BWP30P140LVT U9838 ( .A1(n6676), .A2(n6675), .ZN(N5594) );
  AOI22D1BWP30P140LVT U9839 ( .A1(i_data_bus[888]), .A2(n6723), .B1(
        i_data_bus[856]), .B2(n6722), .ZN(n6678) );
  AOI22D1BWP30P140LVT U9840 ( .A1(i_data_bus[792]), .A2(n6720), .B1(
        i_data_bus[824]), .B2(n6721), .ZN(n6677) );
  ND2D1BWP30P140LVT U9841 ( .A1(n6678), .A2(n6677), .ZN(N5593) );
  AOI22D1BWP30P140LVT U9842 ( .A1(i_data_bus[791]), .A2(n6720), .B1(
        i_data_bus[855]), .B2(n6722), .ZN(n6680) );
  AOI22D1BWP30P140LVT U9843 ( .A1(i_data_bus[887]), .A2(n6723), .B1(
        i_data_bus[823]), .B2(n6721), .ZN(n6679) );
  ND2D1BWP30P140LVT U9844 ( .A1(n6680), .A2(n6679), .ZN(N5592) );
  AOI22D1BWP30P140LVT U9845 ( .A1(i_data_bus[787]), .A2(n6720), .B1(
        i_data_bus[851]), .B2(n6722), .ZN(n6682) );
  AOI22D1BWP30P140LVT U9846 ( .A1(i_data_bus[883]), .A2(n6723), .B1(
        i_data_bus[819]), .B2(n6721), .ZN(n6681) );
  ND2D1BWP30P140LVT U9847 ( .A1(n6682), .A2(n6681), .ZN(N5588) );
  AOI22D1BWP30P140LVT U9848 ( .A1(i_data_bus[779]), .A2(n6720), .B1(
        i_data_bus[875]), .B2(n6723), .ZN(n6684) );
  AOI22D1BWP30P140LVT U9849 ( .A1(i_data_bus[843]), .A2(n6722), .B1(
        i_data_bus[811]), .B2(n6721), .ZN(n6683) );
  ND2D1BWP30P140LVT U9850 ( .A1(n6684), .A2(n6683), .ZN(N5580) );
  AOI22D1BWP30P140LVT U9851 ( .A1(i_data_bus[873]), .A2(n6723), .B1(
        i_data_bus[777]), .B2(n6720), .ZN(n6686) );
  AOI22D1BWP30P140LVT U9852 ( .A1(i_data_bus[841]), .A2(n6722), .B1(
        i_data_bus[809]), .B2(n6721), .ZN(n6685) );
  ND2D1BWP30P140LVT U9853 ( .A1(n6686), .A2(n6685), .ZN(N5578) );
  AOI22D1BWP30P140LVT U9854 ( .A1(i_data_bus[772]), .A2(n6720), .B1(
        i_data_bus[836]), .B2(n6722), .ZN(n6688) );
  AOI22D1BWP30P140LVT U9855 ( .A1(i_data_bus[868]), .A2(n6723), .B1(
        i_data_bus[804]), .B2(n6721), .ZN(n6687) );
  ND2D1BWP30P140LVT U9856 ( .A1(n6688), .A2(n6687), .ZN(N5573) );
  NR3D0P7BWP30P140LVT U9857 ( .A1(i_cmd[176]), .A2(i_cmd[168]), .A3(i_cmd[184]), .ZN(n11156) );
  INR4D1BWP30P140LVT U9858 ( .A1(i_cmd[184]), .B1(i_cmd[168]), .B2(n6692), 
        .B3(n6690), .ZN(n6984) );
  AOI22D1BWP30P140LVT U9859 ( .A1(i_data_bus[640]), .A2(n6986), .B1(
        i_data_bus[736]), .B2(n6984), .ZN(n6695) );
  OR2D1BWP30P140LVT U9860 ( .A1(i_cmd[184]), .A2(i_cmd[168]), .Z(n11160) );
  INR4D1BWP30P140LVT U9861 ( .A1(i_cmd[176]), .B1(i_cmd[160]), .B2(n6691), 
        .B3(n11160), .ZN(n6985) );
  INR4D1BWP30P140LVT U9862 ( .A1(i_cmd[168]), .B1(i_cmd[184]), .B2(n6693), 
        .B3(n6692), .ZN(n6987) );
  AOI22D1BWP30P140LVT U9863 ( .A1(i_data_bus[704]), .A2(n6985), .B1(
        i_data_bus[672]), .B2(n6987), .ZN(n6694) );
  ND2D1BWP30P140LVT U9864 ( .A1(n6695), .A2(n6694), .ZN(N1643) );
  AOI22D1BWP30P140LVT U9865 ( .A1(n6986), .A2(i_data_bus[671]), .B1(n6984), 
        .B2(i_data_bus[767]), .ZN(n6697) );
  AOI22D1BWP30P140LVT U9866 ( .A1(n6985), .A2(i_data_bus[735]), .B1(n6987), 
        .B2(i_data_bus[703]), .ZN(n6696) );
  ND2D1BWP30P140LVT U9867 ( .A1(n6697), .A2(n6696), .ZN(N1674) );
  AOI22D1BWP30P140LVT U9868 ( .A1(n6986), .A2(i_data_bus[661]), .B1(n6984), 
        .B2(i_data_bus[757]), .ZN(n6699) );
  AOI22D1BWP30P140LVT U9869 ( .A1(n6985), .A2(i_data_bus[725]), .B1(n6987), 
        .B2(i_data_bus[693]), .ZN(n6698) );
  ND2D1BWP30P140LVT U9870 ( .A1(n6699), .A2(n6698), .ZN(N1664) );
  AOI22D1BWP30P140LVT U9871 ( .A1(n6986), .A2(i_data_bus[660]), .B1(n6984), 
        .B2(i_data_bus[756]), .ZN(n6701) );
  AOI22D1BWP30P140LVT U9872 ( .A1(n6985), .A2(i_data_bus[724]), .B1(n6987), 
        .B2(i_data_bus[692]), .ZN(n6700) );
  ND2D1BWP30P140LVT U9873 ( .A1(n6701), .A2(n6700), .ZN(N1663) );
  AOI22D1BWP30P140LVT U9874 ( .A1(n6986), .A2(i_data_bus[658]), .B1(n6984), 
        .B2(i_data_bus[754]), .ZN(n6703) );
  AOI22D1BWP30P140LVT U9875 ( .A1(n6985), .A2(i_data_bus[722]), .B1(n6987), 
        .B2(i_data_bus[690]), .ZN(n6702) );
  ND2D1BWP30P140LVT U9876 ( .A1(n6703), .A2(n6702), .ZN(N1661) );
  AOI22D1BWP30P140LVT U9877 ( .A1(n6986), .A2(i_data_bus[656]), .B1(n6984), 
        .B2(i_data_bus[752]), .ZN(n6705) );
  AOI22D1BWP30P140LVT U9878 ( .A1(n6985), .A2(i_data_bus[720]), .B1(n6987), 
        .B2(i_data_bus[688]), .ZN(n6704) );
  ND2D1BWP30P140LVT U9879 ( .A1(n6705), .A2(n6704), .ZN(N1659) );
  AOI22D1BWP30P140LVT U9880 ( .A1(n6986), .A2(i_data_bus[646]), .B1(n6984), 
        .B2(i_data_bus[742]), .ZN(n6707) );
  AOI22D1BWP30P140LVT U9881 ( .A1(n6985), .A2(i_data_bus[710]), .B1(n6987), 
        .B2(i_data_bus[678]), .ZN(n6706) );
  ND2D1BWP30P140LVT U9882 ( .A1(n6707), .A2(n6706), .ZN(N1649) );
  AOI22D1BWP30P140LVT U9883 ( .A1(n6986), .A2(i_data_bus[645]), .B1(n6984), 
        .B2(i_data_bus[741]), .ZN(n6709) );
  AOI22D1BWP30P140LVT U9884 ( .A1(n6985), .A2(i_data_bus[709]), .B1(n6987), 
        .B2(i_data_bus[677]), .ZN(n6708) );
  ND2D1BWP30P140LVT U9885 ( .A1(n6709), .A2(n6708), .ZN(N1648) );
  AOI22D1BWP30P140LVT U9886 ( .A1(i_data_bus[893]), .A2(n6723), .B1(
        i_data_bus[829]), .B2(n6721), .ZN(n6711) );
  AOI22D1BWP30P140LVT U9887 ( .A1(i_data_bus[797]), .A2(n6720), .B1(
        i_data_bus[861]), .B2(n6722), .ZN(n6710) );
  ND2D1BWP30P140LVT U9888 ( .A1(n6711), .A2(n6710), .ZN(N5598) );
  AOI22D1BWP30P140LVT U9889 ( .A1(i_data_bus[818]), .A2(n6721), .B1(
        i_data_bus[882]), .B2(n6723), .ZN(n6713) );
  AOI22D1BWP30P140LVT U9890 ( .A1(i_data_bus[786]), .A2(n6720), .B1(
        i_data_bus[850]), .B2(n6722), .ZN(n6712) );
  ND2D1BWP30P140LVT U9891 ( .A1(n6713), .A2(n6712), .ZN(N5587) );
  AOI22D1BWP30P140LVT U9892 ( .A1(i_data_bus[879]), .A2(n6723), .B1(
        i_data_bus[783]), .B2(n6720), .ZN(n6715) );
  AOI22D1BWP30P140LVT U9893 ( .A1(i_data_bus[815]), .A2(n6721), .B1(
        i_data_bus[847]), .B2(n6722), .ZN(n6714) );
  ND2D1BWP30P140LVT U9894 ( .A1(n6715), .A2(n6714), .ZN(N5584) );
  AOI22D1BWP30P140LVT U9895 ( .A1(i_data_bus[775]), .A2(n6720), .B1(
        i_data_bus[807]), .B2(n6721), .ZN(n6717) );
  AOI22D1BWP30P140LVT U9896 ( .A1(i_data_bus[871]), .A2(n6723), .B1(
        i_data_bus[839]), .B2(n6722), .ZN(n6716) );
  ND2D1BWP30P140LVT U9897 ( .A1(n6717), .A2(n6716), .ZN(N5576) );
  AOI22D1BWP30P140LVT U9898 ( .A1(i_data_bus[869]), .A2(n6723), .B1(
        i_data_bus[773]), .B2(n6720), .ZN(n6719) );
  AOI22D1BWP30P140LVT U9899 ( .A1(i_data_bus[805]), .A2(n6721), .B1(
        i_data_bus[837]), .B2(n6722), .ZN(n6718) );
  ND2D1BWP30P140LVT U9900 ( .A1(n6719), .A2(n6718), .ZN(N5574) );
  AOI22D1BWP30P140LVT U9901 ( .A1(i_data_bus[801]), .A2(n6721), .B1(
        i_data_bus[769]), .B2(n6720), .ZN(n6725) );
  AOI22D1BWP30P140LVT U9902 ( .A1(i_data_bus[865]), .A2(n6723), .B1(
        i_data_bus[833]), .B2(n6722), .ZN(n6724) );
  ND2D1BWP30P140LVT U9903 ( .A1(n6725), .A2(n6724), .ZN(N5570) );
  AOI22D1BWP30P140LVT U9904 ( .A1(i_data_bus[797]), .A2(n6758), .B1(
        i_data_bus[861]), .B2(n6760), .ZN(n6727) );
  AOI22D1BWP30P140LVT U9905 ( .A1(i_data_bus[893]), .A2(n6761), .B1(
        i_data_bus[829]), .B2(n6759), .ZN(n6726) );
  ND2D1BWP30P140LVT U9906 ( .A1(n6727), .A2(n6726), .ZN(N7344) );
  AOI22D1BWP30P140LVT U9907 ( .A1(i_data_bus[892]), .A2(n6761), .B1(
        i_data_bus[860]), .B2(n6760), .ZN(n6729) );
  AOI22D1BWP30P140LVT U9908 ( .A1(i_data_bus[796]), .A2(n6758), .B1(
        i_data_bus[828]), .B2(n6759), .ZN(n6728) );
  ND2D1BWP30P140LVT U9909 ( .A1(n6729), .A2(n6728), .ZN(N7343) );
  AOI22D1BWP30P140LVT U9910 ( .A1(i_data_bus[890]), .A2(n6761), .B1(
        i_data_bus[794]), .B2(n6758), .ZN(n6731) );
  AOI22D1BWP30P140LVT U9911 ( .A1(i_data_bus[858]), .A2(n6760), .B1(
        i_data_bus[826]), .B2(n6759), .ZN(n6730) );
  ND2D1BWP30P140LVT U9912 ( .A1(n6731), .A2(n6730), .ZN(N7341) );
  AOI22D1BWP30P140LVT U9913 ( .A1(i_data_bus[888]), .A2(n6761), .B1(
        i_data_bus[856]), .B2(n6760), .ZN(n6733) );
  AOI22D1BWP30P140LVT U9914 ( .A1(i_data_bus[792]), .A2(n6758), .B1(
        i_data_bus[824]), .B2(n6759), .ZN(n6732) );
  ND2D1BWP30P140LVT U9915 ( .A1(n6733), .A2(n6732), .ZN(N7339) );
  AOI22D1BWP30P140LVT U9916 ( .A1(i_data_bus[854]), .A2(n6760), .B1(
        i_data_bus[790]), .B2(n6758), .ZN(n6735) );
  AOI22D1BWP30P140LVT U9917 ( .A1(i_data_bus[886]), .A2(n6761), .B1(
        i_data_bus[822]), .B2(n6759), .ZN(n6734) );
  ND2D1BWP30P140LVT U9918 ( .A1(n6735), .A2(n6734), .ZN(N7337) );
  AOI22D1BWP30P140LVT U9919 ( .A1(i_data_bus[789]), .A2(n6758), .B1(
        i_data_bus[885]), .B2(n6761), .ZN(n6737) );
  AOI22D1BWP30P140LVT U9920 ( .A1(i_data_bus[853]), .A2(n6760), .B1(
        i_data_bus[821]), .B2(n6759), .ZN(n6736) );
  ND2D1BWP30P140LVT U9921 ( .A1(n6737), .A2(n6736), .ZN(N7336) );
  AOI22D1BWP30P140LVT U9922 ( .A1(i_data_bus[787]), .A2(n6758), .B1(
        i_data_bus[851]), .B2(n6760), .ZN(n6739) );
  AOI22D1BWP30P140LVT U9923 ( .A1(i_data_bus[883]), .A2(n6761), .B1(
        i_data_bus[819]), .B2(n6759), .ZN(n6738) );
  ND2D1BWP30P140LVT U9924 ( .A1(n6739), .A2(n6738), .ZN(N7334) );
  AOI22D1BWP30P140LVT U9925 ( .A1(i_data_bus[776]), .A2(n6758), .B1(
        i_data_bus[872]), .B2(n6761), .ZN(n6741) );
  AOI22D1BWP30P140LVT U9926 ( .A1(i_data_bus[840]), .A2(n6760), .B1(
        i_data_bus[808]), .B2(n6759), .ZN(n6740) );
  ND2D1BWP30P140LVT U9927 ( .A1(n6741), .A2(n6740), .ZN(N7323) );
  AOI22D1BWP30P140LVT U9928 ( .A1(i_data_bus[895]), .A2(n6761), .B1(
        i_data_bus[831]), .B2(n6759), .ZN(n6743) );
  AOI22D1BWP30P140LVT U9929 ( .A1(i_data_bus[799]), .A2(n6758), .B1(
        i_data_bus[863]), .B2(n6760), .ZN(n6742) );
  ND2D1BWP30P140LVT U9930 ( .A1(n6743), .A2(n6742), .ZN(N7346) );
  AOI22D1BWP30P140LVT U9931 ( .A1(i_data_bus[795]), .A2(n6758), .B1(
        i_data_bus[827]), .B2(n6759), .ZN(n6745) );
  AOI22D1BWP30P140LVT U9932 ( .A1(i_data_bus[891]), .A2(n6761), .B1(
        i_data_bus[859]), .B2(n6760), .ZN(n6744) );
  ND2D1BWP30P140LVT U9933 ( .A1(n6745), .A2(n6744), .ZN(N7342) );
  AOI22D1BWP30P140LVT U9934 ( .A1(i_data_bus[823]), .A2(n6759), .B1(
        i_data_bus[791]), .B2(n6758), .ZN(n6747) );
  AOI22D1BWP30P140LVT U9935 ( .A1(i_data_bus[887]), .A2(n6761), .B1(
        i_data_bus[855]), .B2(n6760), .ZN(n6746) );
  ND2D1BWP30P140LVT U9936 ( .A1(n6747), .A2(n6746), .ZN(N7338) );
  AOI22D1BWP30P140LVT U9937 ( .A1(i_data_bus[881]), .A2(n6761), .B1(
        i_data_bus[817]), .B2(n6759), .ZN(n6749) );
  AOI22D1BWP30P140LVT U9938 ( .A1(i_data_bus[785]), .A2(n6758), .B1(
        i_data_bus[849]), .B2(n6760), .ZN(n6748) );
  ND2D1BWP30P140LVT U9939 ( .A1(n6749), .A2(n6748), .ZN(N7332) );
  AOI22D1BWP30P140LVT U9940 ( .A1(i_data_bus[874]), .A2(n6761), .B1(
        i_data_bus[810]), .B2(n6759), .ZN(n6751) );
  AOI22D1BWP30P140LVT U9941 ( .A1(i_data_bus[778]), .A2(n6758), .B1(
        i_data_bus[842]), .B2(n6760), .ZN(n6750) );
  ND2D1BWP30P140LVT U9942 ( .A1(n6751), .A2(n6750), .ZN(N7325) );
  AOI22D1BWP30P140LVT U9943 ( .A1(i_data_bus[871]), .A2(n6761), .B1(
        i_data_bus[807]), .B2(n6759), .ZN(n6753) );
  AOI22D1BWP30P140LVT U9944 ( .A1(i_data_bus[775]), .A2(n6758), .B1(
        i_data_bus[839]), .B2(n6760), .ZN(n6752) );
  ND2D1BWP30P140LVT U9945 ( .A1(n6753), .A2(n6752), .ZN(N7322) );
  AOI22D1BWP30P140LVT U9946 ( .A1(i_data_bus[805]), .A2(n6759), .B1(
        i_data_bus[773]), .B2(n6758), .ZN(n6755) );
  AOI22D1BWP30P140LVT U9947 ( .A1(i_data_bus[869]), .A2(n6761), .B1(
        i_data_bus[837]), .B2(n6760), .ZN(n6754) );
  ND2D1BWP30P140LVT U9948 ( .A1(n6755), .A2(n6754), .ZN(N7320) );
  AOI22D1BWP30P140LVT U9949 ( .A1(i_data_bus[772]), .A2(n6758), .B1(
        i_data_bus[804]), .B2(n6759), .ZN(n6757) );
  AOI22D1BWP30P140LVT U9950 ( .A1(i_data_bus[868]), .A2(n6761), .B1(
        i_data_bus[836]), .B2(n6760), .ZN(n6756) );
  ND2D1BWP30P140LVT U9951 ( .A1(n6757), .A2(n6756), .ZN(N7319) );
  AOI22D1BWP30P140LVT U9952 ( .A1(i_data_bus[801]), .A2(n6759), .B1(
        i_data_bus[769]), .B2(n6758), .ZN(n6763) );
  AOI22D1BWP30P140LVT U9953 ( .A1(i_data_bus[865]), .A2(n6761), .B1(
        i_data_bus[833]), .B2(n6760), .ZN(n6762) );
  ND2D1BWP30P140LVT U9954 ( .A1(n6763), .A2(n6762), .ZN(N7316) );
  AOI22D1BWP30P140LVT U9955 ( .A1(i_data_bus[688]), .A2(n6877), .B1(
        i_data_bus[656]), .B2(n6878), .ZN(n6765) );
  AOI22D1BWP30P140LVT U9956 ( .A1(i_data_bus[720]), .A2(n6876), .B1(
        i_data_bus[752]), .B2(n6879), .ZN(n6764) );
  ND2D1BWP30P140LVT U9957 ( .A1(n6765), .A2(n6764), .ZN(N10945) );
  AOI22D1BWP30P140LVT U9958 ( .A1(i_data_bus[754]), .A2(n6879), .B1(
        i_data_bus[658]), .B2(n6878), .ZN(n6767) );
  AOI22D1BWP30P140LVT U9959 ( .A1(i_data_bus[722]), .A2(n6876), .B1(
        i_data_bus[690]), .B2(n6877), .ZN(n6766) );
  ND2D1BWP30P140LVT U9960 ( .A1(n6767), .A2(n6766), .ZN(N10947) );
  AOI22D1BWP30P140LVT U9961 ( .A1(i_data_bus[743]), .A2(n6879), .B1(
        i_data_bus[647]), .B2(n6878), .ZN(n6769) );
  AOI22D1BWP30P140LVT U9962 ( .A1(i_data_bus[711]), .A2(n6876), .B1(
        i_data_bus[679]), .B2(n6877), .ZN(n6768) );
  ND2D1BWP30P140LVT U9963 ( .A1(n6769), .A2(n6768), .ZN(N10936) );
  AOI22D1BWP30P140LVT U9964 ( .A1(n6985), .A2(i_data_bus[732]), .B1(n6987), 
        .B2(i_data_bus[700]), .ZN(n6771) );
  AOI22D1BWP30P140LVT U9965 ( .A1(n6986), .A2(i_data_bus[668]), .B1(n6984), 
        .B2(i_data_bus[764]), .ZN(n6770) );
  ND2D1BWP30P140LVT U9966 ( .A1(n6771), .A2(n6770), .ZN(N1671) );
  AOI22D1BWP30P140LVT U9967 ( .A1(n6985), .A2(i_data_bus[727]), .B1(n6987), 
        .B2(i_data_bus[695]), .ZN(n6773) );
  AOI22D1BWP30P140LVT U9968 ( .A1(n6986), .A2(i_data_bus[663]), .B1(n6984), 
        .B2(i_data_bus[759]), .ZN(n6772) );
  ND2D1BWP30P140LVT U9969 ( .A1(n6773), .A2(n6772), .ZN(N1666) );
  AOI22D1BWP30P140LVT U9970 ( .A1(n6985), .A2(i_data_bus[723]), .B1(n6987), 
        .B2(i_data_bus[691]), .ZN(n6775) );
  AOI22D1BWP30P140LVT U9971 ( .A1(n6986), .A2(i_data_bus[659]), .B1(n6984), 
        .B2(i_data_bus[755]), .ZN(n6774) );
  ND2D1BWP30P140LVT U9972 ( .A1(n6775), .A2(n6774), .ZN(N1662) );
  AOI22D1BWP30P140LVT U9973 ( .A1(n6985), .A2(i_data_bus[714]), .B1(n6987), 
        .B2(i_data_bus[682]), .ZN(n6777) );
  AOI22D1BWP30P140LVT U9974 ( .A1(n6986), .A2(i_data_bus[650]), .B1(n6984), 
        .B2(i_data_bus[746]), .ZN(n6776) );
  ND2D1BWP30P140LVT U9975 ( .A1(n6777), .A2(n6776), .ZN(N1653) );
  AOI22D1BWP30P140LVT U9976 ( .A1(i_data_bus[697]), .A2(n6877), .B1(
        i_data_bus[665]), .B2(n6878), .ZN(n6779) );
  AOI22D1BWP30P140LVT U9977 ( .A1(i_data_bus[761]), .A2(n6879), .B1(
        i_data_bus[729]), .B2(n6876), .ZN(n6778) );
  ND2D1BWP30P140LVT U9978 ( .A1(n6779), .A2(n6778), .ZN(N10954) );
  AOI22D1BWP30P140LVT U9979 ( .A1(i_data_bus[766]), .A2(n6885), .B1(
        i_data_bus[670]), .B2(n6884), .ZN(n6781) );
  AOI22D1BWP30P140LVT U9980 ( .A1(i_data_bus[734]), .A2(n6883), .B1(
        i_data_bus[702]), .B2(n6882), .ZN(n6780) );
  ND2D1BWP30P140LVT U9981 ( .A1(n6781), .A2(n6780), .ZN(N8235) );
  AOI22D1BWP30P140LVT U9982 ( .A1(i_data_bus[733]), .A2(n6883), .B1(
        i_data_bus[669]), .B2(n6884), .ZN(n6783) );
  AOI22D1BWP30P140LVT U9983 ( .A1(i_data_bus[765]), .A2(n6885), .B1(
        i_data_bus[701]), .B2(n6882), .ZN(n6782) );
  ND2D1BWP30P140LVT U9984 ( .A1(n6783), .A2(n6782), .ZN(N8234) );
  AOI22D1BWP30P140LVT U9985 ( .A1(i_data_bus[762]), .A2(n6885), .B1(
        i_data_bus[666]), .B2(n6884), .ZN(n6785) );
  AOI22D1BWP30P140LVT U9986 ( .A1(i_data_bus[730]), .A2(n6883), .B1(
        i_data_bus[698]), .B2(n6882), .ZN(n6784) );
  ND2D1BWP30P140LVT U9987 ( .A1(n6785), .A2(n6784), .ZN(N8231) );
  AOI22D1BWP30P140LVT U9988 ( .A1(i_data_bus[747]), .A2(n6885), .B1(
        i_data_bus[651]), .B2(n6884), .ZN(n6787) );
  AOI22D1BWP30P140LVT U9989 ( .A1(i_data_bus[715]), .A2(n6883), .B1(
        i_data_bus[683]), .B2(n6882), .ZN(n6786) );
  ND2D1BWP30P140LVT U9990 ( .A1(n6787), .A2(n6786), .ZN(N8216) );
  AOI22D1BWP30P140LVT U9991 ( .A1(i_data_bus[711]), .A2(n6883), .B1(
        i_data_bus[647]), .B2(n6884), .ZN(n6789) );
  AOI22D1BWP30P140LVT U9992 ( .A1(i_data_bus[743]), .A2(n6885), .B1(
        i_data_bus[679]), .B2(n6882), .ZN(n6788) );
  ND2D1BWP30P140LVT U9993 ( .A1(n6789), .A2(n6788), .ZN(N8212) );
  AOI22D1BWP30P140LVT U9994 ( .A1(i_data_bus[708]), .A2(n6883), .B1(
        i_data_bus[644]), .B2(n6884), .ZN(n6791) );
  AOI22D1BWP30P140LVT U9995 ( .A1(i_data_bus[740]), .A2(n6885), .B1(
        i_data_bus[676]), .B2(n6882), .ZN(n6790) );
  ND2D1BWP30P140LVT U9996 ( .A1(n6791), .A2(n6790), .ZN(N8209) );
  AOI22D1BWP30P140LVT U9997 ( .A1(i_data_bus[725]), .A2(n6883), .B1(
        i_data_bus[661]), .B2(n6884), .ZN(n6793) );
  AOI22D1BWP30P140LVT U9998 ( .A1(i_data_bus[693]), .A2(n6882), .B1(
        i_data_bus[757]), .B2(n6885), .ZN(n6792) );
  ND2D1BWP30P140LVT U9999 ( .A1(n6793), .A2(n6792), .ZN(N8226) );
  AOI22D1BWP30P140LVT U10000 ( .A1(i_data_bus[690]), .A2(n6882), .B1(
        i_data_bus[658]), .B2(n6884), .ZN(n6795) );
  AOI22D1BWP30P140LVT U10001 ( .A1(i_data_bus[722]), .A2(n6883), .B1(
        i_data_bus[754]), .B2(n6885), .ZN(n6794) );
  ND2D1BWP30P140LVT U10002 ( .A1(n6795), .A2(n6794), .ZN(N8223) );
  AOI22D1BWP30P140LVT U10003 ( .A1(i_data_bus[688]), .A2(n6882), .B1(
        i_data_bus[656]), .B2(n6884), .ZN(n6797) );
  AOI22D1BWP30P140LVT U10004 ( .A1(i_data_bus[720]), .A2(n6883), .B1(
        i_data_bus[752]), .B2(n6885), .ZN(n6796) );
  ND2D1BWP30P140LVT U10005 ( .A1(n6797), .A2(n6796), .ZN(N8221) );
  AOI22D1BWP30P140LVT U10006 ( .A1(i_data_bus[710]), .A2(n6883), .B1(
        i_data_bus[646]), .B2(n6884), .ZN(n6799) );
  AOI22D1BWP30P140LVT U10007 ( .A1(i_data_bus[678]), .A2(n6882), .B1(
        i_data_bus[742]), .B2(n6885), .ZN(n6798) );
  ND2D1BWP30P140LVT U10008 ( .A1(n6799), .A2(n6798), .ZN(N8211) );
  AOI22D1BWP30P140LVT U10009 ( .A1(i_data_bus[672]), .A2(n6882), .B1(
        i_data_bus[640]), .B2(n6884), .ZN(n6801) );
  AOI22D1BWP30P140LVT U10010 ( .A1(i_data_bus[704]), .A2(n6883), .B1(
        i_data_bus[736]), .B2(n6885), .ZN(n6800) );
  ND2D1BWP30P140LVT U10011 ( .A1(n6801), .A2(n6800), .ZN(N8205) );
  AOI22D1BWP30P140LVT U10012 ( .A1(i_data_bus[689]), .A2(n6882), .B1(
        i_data_bus[657]), .B2(n6884), .ZN(n6803) );
  AOI22D1BWP30P140LVT U10013 ( .A1(i_data_bus[753]), .A2(n6885), .B1(
        i_data_bus[721]), .B2(n6883), .ZN(n6802) );
  ND2D1BWP30P140LVT U10014 ( .A1(n6803), .A2(n6802), .ZN(N8222) );
  AOI22D1BWP30P140LVT U10015 ( .A1(i_data_bus[680]), .A2(n6882), .B1(
        i_data_bus[648]), .B2(n6884), .ZN(n6805) );
  AOI22D1BWP30P140LVT U10016 ( .A1(i_data_bus[744]), .A2(n6885), .B1(
        i_data_bus[712]), .B2(n6883), .ZN(n6804) );
  ND2D1BWP30P140LVT U10017 ( .A1(n6805), .A2(n6804), .ZN(N8213) );
  AOI22D1BWP30P140LVT U10018 ( .A1(i_data_bus[674]), .A2(n6882), .B1(
        i_data_bus[642]), .B2(n6884), .ZN(n6807) );
  AOI22D1BWP30P140LVT U10019 ( .A1(i_data_bus[738]), .A2(n6885), .B1(
        i_data_bus[706]), .B2(n6883), .ZN(n6806) );
  ND2D1BWP30P140LVT U10020 ( .A1(n6807), .A2(n6806), .ZN(N8207) );
  AOI22D1BWP30P140LVT U10021 ( .A1(i_data_bus[703]), .A2(n6909), .B1(
        i_data_bus[671]), .B2(n6910), .ZN(n6809) );
  AOI22D1BWP30P140LVT U10022 ( .A1(i_data_bus[735]), .A2(n6911), .B1(
        i_data_bus[767]), .B2(n6908), .ZN(n6808) );
  ND2D1BWP30P140LVT U10023 ( .A1(n6809), .A2(n6808), .ZN(N5512) );
  AOI22D1BWP30P140LVT U10024 ( .A1(i_data_bus[766]), .A2(n6908), .B1(
        i_data_bus[670]), .B2(n6910), .ZN(n6811) );
  AOI22D1BWP30P140LVT U10025 ( .A1(i_data_bus[734]), .A2(n6911), .B1(
        i_data_bus[702]), .B2(n6909), .ZN(n6810) );
  ND2D1BWP30P140LVT U10026 ( .A1(n6811), .A2(n6810), .ZN(N5511) );
  AOI22D1BWP30P140LVT U10027 ( .A1(i_data_bus[762]), .A2(n6908), .B1(
        i_data_bus[666]), .B2(n6910), .ZN(n6813) );
  AOI22D1BWP30P140LVT U10028 ( .A1(i_data_bus[730]), .A2(n6911), .B1(
        i_data_bus[698]), .B2(n6909), .ZN(n6812) );
  ND2D1BWP30P140LVT U10029 ( .A1(n6813), .A2(n6812), .ZN(N5507) );
  AOI22D1BWP30P140LVT U10030 ( .A1(i_data_bus[754]), .A2(n6908), .B1(
        i_data_bus[658]), .B2(n6910), .ZN(n6815) );
  AOI22D1BWP30P140LVT U10031 ( .A1(i_data_bus[722]), .A2(n6911), .B1(
        i_data_bus[690]), .B2(n6909), .ZN(n6814) );
  ND2D1BWP30P140LVT U10032 ( .A1(n6815), .A2(n6814), .ZN(N5499) );
  AOI22D1BWP30P140LVT U10033 ( .A1(i_data_bus[742]), .A2(n6925), .B1(
        i_data_bus[646]), .B2(n6924), .ZN(n6817) );
  AOI22D1BWP30P140LVT U10034 ( .A1(i_data_bus[678]), .A2(n6923), .B1(
        i_data_bus[710]), .B2(n6922), .ZN(n6816) );
  ND2D1BWP30P140LVT U10035 ( .A1(n6817), .A2(n6816), .ZN(N9829) );
  AOI22D1BWP30P140LVT U10036 ( .A1(i_data_bus[693]), .A2(n6923), .B1(
        i_data_bus[661]), .B2(n6924), .ZN(n6819) );
  AOI22D1BWP30P140LVT U10037 ( .A1(i_data_bus[725]), .A2(n6922), .B1(
        i_data_bus[757]), .B2(n6925), .ZN(n6818) );
  ND2D1BWP30P140LVT U10038 ( .A1(n6819), .A2(n6818), .ZN(N9844) );
  AOI22D1BWP30P140LVT U10039 ( .A1(i_data_bus[724]), .A2(n6922), .B1(
        i_data_bus[660]), .B2(n6924), .ZN(n6821) );
  AOI22D1BWP30P140LVT U10040 ( .A1(i_data_bus[692]), .A2(n6923), .B1(
        i_data_bus[756]), .B2(n6925), .ZN(n6820) );
  ND2D1BWP30P140LVT U10041 ( .A1(n6821), .A2(n6820), .ZN(N9843) );
  AOI22D1BWP30P140LVT U10042 ( .A1(i_data_bus[722]), .A2(n6922), .B1(
        i_data_bus[658]), .B2(n6924), .ZN(n6823) );
  AOI22D1BWP30P140LVT U10043 ( .A1(i_data_bus[690]), .A2(n6923), .B1(
        i_data_bus[754]), .B2(n6925), .ZN(n6822) );
  ND2D1BWP30P140LVT U10044 ( .A1(n6823), .A2(n6822), .ZN(N9841) );
  AOI22D1BWP30P140LVT U10045 ( .A1(i_data_bus[688]), .A2(n6923), .B1(
        i_data_bus[656]), .B2(n6924), .ZN(n6825) );
  AOI22D1BWP30P140LVT U10046 ( .A1(i_data_bus[720]), .A2(n6922), .B1(
        i_data_bus[752]), .B2(n6925), .ZN(n6824) );
  ND2D1BWP30P140LVT U10047 ( .A1(n6825), .A2(n6824), .ZN(N9839) );
  AOI22D1BWP30P140LVT U10048 ( .A1(i_data_bus[677]), .A2(n6923), .B1(
        i_data_bus[645]), .B2(n6924), .ZN(n6827) );
  AOI22D1BWP30P140LVT U10049 ( .A1(i_data_bus[709]), .A2(n6922), .B1(
        i_data_bus[741]), .B2(n6925), .ZN(n6826) );
  ND2D1BWP30P140LVT U10050 ( .A1(n6827), .A2(n6826), .ZN(N9828) );
  AOI22D1BWP30P140LVT U10051 ( .A1(i_data_bus[704]), .A2(n6922), .B1(
        i_data_bus[640]), .B2(n6924), .ZN(n6829) );
  AOI22D1BWP30P140LVT U10052 ( .A1(i_data_bus[672]), .A2(n6923), .B1(
        i_data_bus[736]), .B2(n6925), .ZN(n6828) );
  ND2D1BWP30P140LVT U10053 ( .A1(n6829), .A2(n6828), .ZN(N9823) );
  AOI22D1BWP30P140LVT U10054 ( .A1(i_data_bus[730]), .A2(n6922), .B1(
        i_data_bus[666]), .B2(n6924), .ZN(n6831) );
  AOI22D1BWP30P140LVT U10055 ( .A1(i_data_bus[762]), .A2(n6925), .B1(
        i_data_bus[698]), .B2(n6923), .ZN(n6830) );
  ND2D1BWP30P140LVT U10056 ( .A1(n6831), .A2(n6830), .ZN(N9849) );
  AOI22D1BWP30P140LVT U10057 ( .A1(i_data_bus[721]), .A2(n6922), .B1(
        i_data_bus[657]), .B2(n6924), .ZN(n6833) );
  AOI22D1BWP30P140LVT U10058 ( .A1(i_data_bus[753]), .A2(n6925), .B1(
        i_data_bus[689]), .B2(n6923), .ZN(n6832) );
  ND2D1BWP30P140LVT U10059 ( .A1(n6833), .A2(n6832), .ZN(N9840) );
  AOI22D1BWP30P140LVT U10060 ( .A1(i_data_bus[715]), .A2(n6922), .B1(
        i_data_bus[651]), .B2(n6924), .ZN(n6835) );
  AOI22D1BWP30P140LVT U10061 ( .A1(i_data_bus[747]), .A2(n6925), .B1(
        i_data_bus[683]), .B2(n6923), .ZN(n6834) );
  ND2D1BWP30P140LVT U10062 ( .A1(n6835), .A2(n6834), .ZN(N9834) );
  AOI22D1BWP30P140LVT U10063 ( .A1(i_data_bus[712]), .A2(n6922), .B1(
        i_data_bus[648]), .B2(n6924), .ZN(n6837) );
  AOI22D1BWP30P140LVT U10064 ( .A1(i_data_bus[744]), .A2(n6925), .B1(
        i_data_bus[680]), .B2(n6923), .ZN(n6836) );
  ND2D1BWP30P140LVT U10065 ( .A1(n6837), .A2(n6836), .ZN(N9831) );
  AOI22D1BWP30P140LVT U10066 ( .A1(i_data_bus[698]), .A2(n6943), .B1(
        i_data_bus[666]), .B2(n6942), .ZN(n6839) );
  AOI22D1BWP30P140LVT U10067 ( .A1(i_data_bus[730]), .A2(n6941), .B1(
        i_data_bus[762]), .B2(n6940), .ZN(n6838) );
  ND2D1BWP30P140LVT U10068 ( .A1(n6839), .A2(n6838), .ZN(N2783) );
  AOI22D1BWP30P140LVT U10069 ( .A1(i_data_bus[693]), .A2(n6943), .B1(
        i_data_bus[661]), .B2(n6942), .ZN(n6841) );
  AOI22D1BWP30P140LVT U10070 ( .A1(i_data_bus[725]), .A2(n6941), .B1(
        i_data_bus[757]), .B2(n6940), .ZN(n6840) );
  ND2D1BWP30P140LVT U10071 ( .A1(n6841), .A2(n6840), .ZN(N2778) );
  AOI22D1BWP30P140LVT U10072 ( .A1(i_data_bus[692]), .A2(n6943), .B1(
        i_data_bus[660]), .B2(n6942), .ZN(n6843) );
  AOI22D1BWP30P140LVT U10073 ( .A1(i_data_bus[724]), .A2(n6941), .B1(
        i_data_bus[756]), .B2(n6940), .ZN(n6842) );
  ND2D1BWP30P140LVT U10074 ( .A1(n6843), .A2(n6842), .ZN(N2777) );
  AOI22D1BWP30P140LVT U10075 ( .A1(i_data_bus[722]), .A2(n6941), .B1(
        i_data_bus[658]), .B2(n6942), .ZN(n6845) );
  AOI22D1BWP30P140LVT U10076 ( .A1(i_data_bus[690]), .A2(n6943), .B1(
        i_data_bus[754]), .B2(n6940), .ZN(n6844) );
  ND2D1BWP30P140LVT U10077 ( .A1(n6845), .A2(n6844), .ZN(N2775) );
  AOI22D1BWP30P140LVT U10078 ( .A1(i_data_bus[720]), .A2(n6941), .B1(
        i_data_bus[656]), .B2(n6942), .ZN(n6847) );
  AOI22D1BWP30P140LVT U10079 ( .A1(i_data_bus[688]), .A2(n6943), .B1(
        i_data_bus[752]), .B2(n6940), .ZN(n6846) );
  ND2D1BWP30P140LVT U10080 ( .A1(n6847), .A2(n6846), .ZN(N2773) );
  AOI22D1BWP30P140LVT U10081 ( .A1(i_data_bus[715]), .A2(n6941), .B1(
        i_data_bus[651]), .B2(n6942), .ZN(n6849) );
  AOI22D1BWP30P140LVT U10082 ( .A1(i_data_bus[747]), .A2(n6940), .B1(
        i_data_bus[683]), .B2(n6943), .ZN(n6848) );
  ND2D1BWP30P140LVT U10083 ( .A1(n6849), .A2(n6848), .ZN(N2768) );
  AOI22D1BWP30P140LVT U10084 ( .A1(i_data_bus[741]), .A2(n6940), .B1(
        i_data_bus[645]), .B2(n6942), .ZN(n6851) );
  AOI22D1BWP30P140LVT U10085 ( .A1(i_data_bus[709]), .A2(n6941), .B1(
        i_data_bus[677]), .B2(n6943), .ZN(n6850) );
  ND2D1BWP30P140LVT U10086 ( .A1(n6851), .A2(n6850), .ZN(N2762) );
  AOI22D1BWP30P140LVT U10087 ( .A1(i_data_bus[708]), .A2(n6941), .B1(
        i_data_bus[644]), .B2(n6942), .ZN(n6853) );
  AOI22D1BWP30P140LVT U10088 ( .A1(i_data_bus[740]), .A2(n6940), .B1(
        i_data_bus[676]), .B2(n6943), .ZN(n6852) );
  ND2D1BWP30P140LVT U10089 ( .A1(n6853), .A2(n6852), .ZN(N2761) );
  AOI22D1BWP30P140LVT U10090 ( .A1(i_data_bus[680]), .A2(n6943), .B1(
        i_data_bus[648]), .B2(n6942), .ZN(n6855) );
  AOI22D1BWP30P140LVT U10091 ( .A1(i_data_bus[744]), .A2(n6940), .B1(
        i_data_bus[712]), .B2(n6941), .ZN(n6854) );
  ND2D1BWP30P140LVT U10092 ( .A1(n6855), .A2(n6854), .ZN(N2765) );
  AOI22D1BWP30P140LVT U10093 ( .A1(i_data_bus[738]), .A2(n6940), .B1(
        i_data_bus[642]), .B2(n6942), .ZN(n6857) );
  AOI22D1BWP30P140LVT U10094 ( .A1(i_data_bus[674]), .A2(n6943), .B1(
        i_data_bus[706]), .B2(n6941), .ZN(n6856) );
  ND2D1BWP30P140LVT U10095 ( .A1(n6857), .A2(n6856), .ZN(N2759) );
  AOI22D1BWP30P140LVT U10096 ( .A1(i_data_bus[735]), .A2(n6876), .B1(
        i_data_bus[767]), .B2(n6879), .ZN(n6859) );
  AOI22D1BWP30P140LVT U10097 ( .A1(i_data_bus[703]), .A2(n6877), .B1(
        i_data_bus[671]), .B2(n6878), .ZN(n6858) );
  ND2D1BWP30P140LVT U10098 ( .A1(n6859), .A2(n6858), .ZN(N10960) );
  AOI22D1BWP30P140LVT U10099 ( .A1(i_data_bus[765]), .A2(n6879), .B1(
        i_data_bus[701]), .B2(n6877), .ZN(n6861) );
  AOI22D1BWP30P140LVT U10100 ( .A1(i_data_bus[733]), .A2(n6876), .B1(
        i_data_bus[669]), .B2(n6878), .ZN(n6860) );
  ND2D1BWP30P140LVT U10101 ( .A1(n6861), .A2(n6860), .ZN(N10958) );
  AOI22D1BWP30P140LVT U10102 ( .A1(i_data_bus[730]), .A2(n6876), .B1(
        i_data_bus[762]), .B2(n6879), .ZN(n6863) );
  AOI22D1BWP30P140LVT U10103 ( .A1(i_data_bus[698]), .A2(n6877), .B1(
        i_data_bus[666]), .B2(n6878), .ZN(n6862) );
  ND2D1BWP30P140LVT U10104 ( .A1(n6863), .A2(n6862), .ZN(N10955) );
  AOI22D1BWP30P140LVT U10105 ( .A1(i_data_bus[753]), .A2(n6879), .B1(
        i_data_bus[721]), .B2(n6876), .ZN(n6865) );
  AOI22D1BWP30P140LVT U10106 ( .A1(i_data_bus[689]), .A2(n6877), .B1(
        i_data_bus[657]), .B2(n6878), .ZN(n6864) );
  ND2D1BWP30P140LVT U10107 ( .A1(n6865), .A2(n6864), .ZN(N10946) );
  AOI22D1BWP30P140LVT U10108 ( .A1(i_data_bus[747]), .A2(n6879), .B1(
        i_data_bus[683]), .B2(n6877), .ZN(n6867) );
  AOI22D1BWP30P140LVT U10109 ( .A1(i_data_bus[715]), .A2(n6876), .B1(
        i_data_bus[651]), .B2(n6878), .ZN(n6866) );
  ND2D1BWP30P140LVT U10110 ( .A1(n6867), .A2(n6866), .ZN(N10940) );
  AOI22D1BWP30P140LVT U10111 ( .A1(i_data_bus[744]), .A2(n6879), .B1(
        i_data_bus[680]), .B2(n6877), .ZN(n6869) );
  AOI22D1BWP30P140LVT U10112 ( .A1(i_data_bus[712]), .A2(n6876), .B1(
        i_data_bus[648]), .B2(n6878), .ZN(n6868) );
  ND2D1BWP30P140LVT U10113 ( .A1(n6869), .A2(n6868), .ZN(N10937) );
  AOI22D1BWP30P140LVT U10114 ( .A1(i_data_bus[678]), .A2(n6877), .B1(
        i_data_bus[710]), .B2(n6876), .ZN(n6871) );
  AOI22D1BWP30P140LVT U10115 ( .A1(i_data_bus[742]), .A2(n6879), .B1(
        i_data_bus[646]), .B2(n6878), .ZN(n6870) );
  ND2D1BWP30P140LVT U10116 ( .A1(n6871), .A2(n6870), .ZN(N10935) );
  AOI22D1BWP30P140LVT U10117 ( .A1(i_data_bus[709]), .A2(n6876), .B1(
        i_data_bus[741]), .B2(n6879), .ZN(n6873) );
  AOI22D1BWP30P140LVT U10118 ( .A1(i_data_bus[677]), .A2(n6877), .B1(
        i_data_bus[645]), .B2(n6878), .ZN(n6872) );
  ND2D1BWP30P140LVT U10119 ( .A1(n6873), .A2(n6872), .ZN(N10934) );
  AOI22D1BWP30P140LVT U10120 ( .A1(i_data_bus[740]), .A2(n6879), .B1(
        i_data_bus[676]), .B2(n6877), .ZN(n6875) );
  AOI22D1BWP30P140LVT U10121 ( .A1(i_data_bus[708]), .A2(n6876), .B1(
        i_data_bus[644]), .B2(n6878), .ZN(n6874) );
  ND2D1BWP30P140LVT U10122 ( .A1(n6875), .A2(n6874), .ZN(N10933) );
  AOI22D1BWP30P140LVT U10123 ( .A1(i_data_bus[674]), .A2(n6877), .B1(
        i_data_bus[706]), .B2(n6876), .ZN(n6881) );
  AOI22D1BWP30P140LVT U10124 ( .A1(i_data_bus[738]), .A2(n6879), .B1(
        i_data_bus[642]), .B2(n6878), .ZN(n6880) );
  ND2D1BWP30P140LVT U10125 ( .A1(n6881), .A2(n6880), .ZN(N10931) );
  AOI22D1BWP30P140LVT U10126 ( .A1(i_data_bus[709]), .A2(n6883), .B1(
        i_data_bus[677]), .B2(n6882), .ZN(n6887) );
  AOI22D1BWP30P140LVT U10127 ( .A1(i_data_bus[741]), .A2(n6885), .B1(
        i_data_bus[645]), .B2(n6884), .ZN(n6886) );
  ND2D1BWP30P140LVT U10128 ( .A1(n6887), .A2(n6886), .ZN(N8210) );
  AOI22D1BWP30P140LVT U10129 ( .A1(i_data_bus[733]), .A2(n6911), .B1(
        i_data_bus[765]), .B2(n6908), .ZN(n6889) );
  AOI22D1BWP30P140LVT U10130 ( .A1(i_data_bus[701]), .A2(n6909), .B1(
        i_data_bus[669]), .B2(n6910), .ZN(n6888) );
  ND2D1BWP30P140LVT U10131 ( .A1(n6889), .A2(n6888), .ZN(N5510) );
  AOI22D1BWP30P140LVT U10132 ( .A1(i_data_bus[693]), .A2(n6909), .B1(
        i_data_bus[757]), .B2(n6908), .ZN(n6891) );
  AOI22D1BWP30P140LVT U10133 ( .A1(i_data_bus[725]), .A2(n6911), .B1(
        i_data_bus[661]), .B2(n6910), .ZN(n6890) );
  ND2D1BWP30P140LVT U10134 ( .A1(n6891), .A2(n6890), .ZN(N5502) );
  AOI22D1BWP30P140LVT U10135 ( .A1(i_data_bus[721]), .A2(n6911), .B1(
        i_data_bus[689]), .B2(n6909), .ZN(n6893) );
  AOI22D1BWP30P140LVT U10136 ( .A1(i_data_bus[753]), .A2(n6908), .B1(
        i_data_bus[657]), .B2(n6910), .ZN(n6892) );
  ND2D1BWP30P140LVT U10137 ( .A1(n6893), .A2(n6892), .ZN(N5498) );
  AOI22D1BWP30P140LVT U10138 ( .A1(i_data_bus[720]), .A2(n6911), .B1(
        i_data_bus[752]), .B2(n6908), .ZN(n6895) );
  AOI22D1BWP30P140LVT U10139 ( .A1(i_data_bus[688]), .A2(n6909), .B1(
        i_data_bus[656]), .B2(n6910), .ZN(n6894) );
  ND2D1BWP30P140LVT U10140 ( .A1(n6895), .A2(n6894), .ZN(N5497) );
  AOI22D1BWP30P140LVT U10141 ( .A1(i_data_bus[744]), .A2(n6908), .B1(
        i_data_bus[712]), .B2(n6911), .ZN(n6897) );
  AOI22D1BWP30P140LVT U10142 ( .A1(i_data_bus[680]), .A2(n6909), .B1(
        i_data_bus[648]), .B2(n6910), .ZN(n6896) );
  ND2D1BWP30P140LVT U10143 ( .A1(n6897), .A2(n6896), .ZN(N5489) );
  AOI22D1BWP30P140LVT U10144 ( .A1(i_data_bus[711]), .A2(n6911), .B1(
        i_data_bus[743]), .B2(n6908), .ZN(n6899) );
  AOI22D1BWP30P140LVT U10145 ( .A1(i_data_bus[679]), .A2(n6909), .B1(
        i_data_bus[647]), .B2(n6910), .ZN(n6898) );
  ND2D1BWP30P140LVT U10146 ( .A1(n6899), .A2(n6898), .ZN(N5488) );
  AOI22D1BWP30P140LVT U10147 ( .A1(i_data_bus[710]), .A2(n6911), .B1(
        i_data_bus[742]), .B2(n6908), .ZN(n6901) );
  AOI22D1BWP30P140LVT U10148 ( .A1(i_data_bus[678]), .A2(n6909), .B1(
        i_data_bus[646]), .B2(n6910), .ZN(n6900) );
  ND2D1BWP30P140LVT U10149 ( .A1(n6901), .A2(n6900), .ZN(N5487) );
  AOI22D1BWP30P140LVT U10150 ( .A1(i_data_bus[709]), .A2(n6911), .B1(
        i_data_bus[741]), .B2(n6908), .ZN(n6903) );
  AOI22D1BWP30P140LVT U10151 ( .A1(i_data_bus[677]), .A2(n6909), .B1(
        i_data_bus[645]), .B2(n6910), .ZN(n6902) );
  ND2D1BWP30P140LVT U10152 ( .A1(n6903), .A2(n6902), .ZN(N5486) );
  AOI22D1BWP30P140LVT U10153 ( .A1(i_data_bus[740]), .A2(n6908), .B1(
        i_data_bus[676]), .B2(n6909), .ZN(n6905) );
  AOI22D1BWP30P140LVT U10154 ( .A1(i_data_bus[708]), .A2(n6911), .B1(
        i_data_bus[644]), .B2(n6910), .ZN(n6904) );
  ND2D1BWP30P140LVT U10155 ( .A1(n6905), .A2(n6904), .ZN(N5485) );
  AOI22D1BWP30P140LVT U10156 ( .A1(i_data_bus[674]), .A2(n6909), .B1(
        i_data_bus[706]), .B2(n6911), .ZN(n6907) );
  AOI22D1BWP30P140LVT U10157 ( .A1(i_data_bus[738]), .A2(n6908), .B1(
        i_data_bus[642]), .B2(n6910), .ZN(n6906) );
  ND2D1BWP30P140LVT U10158 ( .A1(n6907), .A2(n6906), .ZN(N5483) );
  AOI22D1BWP30P140LVT U10159 ( .A1(i_data_bus[672]), .A2(n6909), .B1(
        i_data_bus[736]), .B2(n6908), .ZN(n6913) );
  AOI22D1BWP30P140LVT U10160 ( .A1(i_data_bus[704]), .A2(n6911), .B1(
        i_data_bus[640]), .B2(n6910), .ZN(n6912) );
  ND2D1BWP30P140LVT U10161 ( .A1(n6913), .A2(n6912), .ZN(N5481) );
  AOI22D1BWP30P140LVT U10162 ( .A1(i_data_bus[703]), .A2(n6923), .B1(
        i_data_bus[767]), .B2(n6925), .ZN(n6915) );
  AOI22D1BWP30P140LVT U10163 ( .A1(i_data_bus[735]), .A2(n6922), .B1(
        i_data_bus[671]), .B2(n6924), .ZN(n6914) );
  ND2D1BWP30P140LVT U10164 ( .A1(n6915), .A2(n6914), .ZN(N9854) );
  AOI22D1BWP30P140LVT U10165 ( .A1(i_data_bus[733]), .A2(n6922), .B1(
        i_data_bus[765]), .B2(n6925), .ZN(n6917) );
  AOI22D1BWP30P140LVT U10166 ( .A1(i_data_bus[701]), .A2(n6923), .B1(
        i_data_bus[669]), .B2(n6924), .ZN(n6916) );
  ND2D1BWP30P140LVT U10167 ( .A1(n6917), .A2(n6916), .ZN(N9852) );
  AOI22D1BWP30P140LVT U10168 ( .A1(i_data_bus[711]), .A2(n6922), .B1(
        i_data_bus[679]), .B2(n6923), .ZN(n6919) );
  AOI22D1BWP30P140LVT U10169 ( .A1(i_data_bus[743]), .A2(n6925), .B1(
        i_data_bus[647]), .B2(n6924), .ZN(n6918) );
  ND2D1BWP30P140LVT U10170 ( .A1(n6919), .A2(n6918), .ZN(N9830) );
  AOI22D1BWP30P140LVT U10171 ( .A1(i_data_bus[708]), .A2(n6922), .B1(
        i_data_bus[676]), .B2(n6923), .ZN(n6921) );
  AOI22D1BWP30P140LVT U10172 ( .A1(i_data_bus[740]), .A2(n6925), .B1(
        i_data_bus[644]), .B2(n6924), .ZN(n6920) );
  ND2D1BWP30P140LVT U10173 ( .A1(n6921), .A2(n6920), .ZN(N9827) );
  AOI22D1BWP30P140LVT U10174 ( .A1(i_data_bus[674]), .A2(n6923), .B1(
        i_data_bus[706]), .B2(n6922), .ZN(n6927) );
  AOI22D1BWP30P140LVT U10175 ( .A1(i_data_bus[738]), .A2(n6925), .B1(
        i_data_bus[642]), .B2(n6924), .ZN(n6926) );
  ND2D1BWP30P140LVT U10176 ( .A1(n6927), .A2(n6926), .ZN(N9825) );
  AOI22D1BWP30P140LVT U10177 ( .A1(i_data_bus[735]), .A2(n6941), .B1(
        i_data_bus[767]), .B2(n6940), .ZN(n6929) );
  AOI22D1BWP30P140LVT U10178 ( .A1(i_data_bus[703]), .A2(n6943), .B1(
        i_data_bus[671]), .B2(n6942), .ZN(n6928) );
  ND2D1BWP30P140LVT U10179 ( .A1(n6929), .A2(n6928), .ZN(N2788) );
  AOI22D1BWP30P140LVT U10180 ( .A1(i_data_bus[733]), .A2(n6941), .B1(
        i_data_bus[701]), .B2(n6943), .ZN(n6931) );
  AOI22D1BWP30P140LVT U10181 ( .A1(i_data_bus[765]), .A2(n6940), .B1(
        i_data_bus[669]), .B2(n6942), .ZN(n6930) );
  ND2D1BWP30P140LVT U10182 ( .A1(n6931), .A2(n6930), .ZN(N2786) );
  AOI22D1BWP30P140LVT U10183 ( .A1(i_data_bus[761]), .A2(n6940), .B1(
        i_data_bus[729]), .B2(n6941), .ZN(n6933) );
  AOI22D1BWP30P140LVT U10184 ( .A1(i_data_bus[697]), .A2(n6943), .B1(
        i_data_bus[665]), .B2(n6942), .ZN(n6932) );
  ND2D1BWP30P140LVT U10185 ( .A1(n6933), .A2(n6932), .ZN(N2782) );
  AOI22D1BWP30P140LVT U10186 ( .A1(i_data_bus[753]), .A2(n6940), .B1(
        i_data_bus[721]), .B2(n6941), .ZN(n6935) );
  AOI22D1BWP30P140LVT U10187 ( .A1(i_data_bus[689]), .A2(n6943), .B1(
        i_data_bus[657]), .B2(n6942), .ZN(n6934) );
  ND2D1BWP30P140LVT U10188 ( .A1(n6935), .A2(n6934), .ZN(N2774) );
  AOI22D1BWP30P140LVT U10189 ( .A1(i_data_bus[743]), .A2(n6940), .B1(
        i_data_bus[679]), .B2(n6943), .ZN(n6937) );
  AOI22D1BWP30P140LVT U10190 ( .A1(i_data_bus[711]), .A2(n6941), .B1(
        i_data_bus[647]), .B2(n6942), .ZN(n6936) );
  ND2D1BWP30P140LVT U10191 ( .A1(n6937), .A2(n6936), .ZN(N2764) );
  AOI22D1BWP30P140LVT U10192 ( .A1(i_data_bus[678]), .A2(n6943), .B1(
        i_data_bus[710]), .B2(n6941), .ZN(n6939) );
  AOI22D1BWP30P140LVT U10193 ( .A1(i_data_bus[742]), .A2(n6940), .B1(
        i_data_bus[646]), .B2(n6942), .ZN(n6938) );
  ND2D1BWP30P140LVT U10194 ( .A1(n6939), .A2(n6938), .ZN(N2763) );
  AOI22D1BWP30P140LVT U10195 ( .A1(i_data_bus[704]), .A2(n6941), .B1(
        i_data_bus[736]), .B2(n6940), .ZN(n6945) );
  AOI22D1BWP30P140LVT U10196 ( .A1(i_data_bus[672]), .A2(n6943), .B1(
        i_data_bus[640]), .B2(n6942), .ZN(n6944) );
  ND2D1BWP30P140LVT U10197 ( .A1(n6945), .A2(n6944), .ZN(N2757) );
  AOI22D1BWP30P140LVT U10198 ( .A1(n6987), .A2(i_data_bus[702]), .B1(n6986), 
        .B2(i_data_bus[670]), .ZN(n6947) );
  AOI22D1BWP30P140LVT U10199 ( .A1(n6985), .A2(i_data_bus[734]), .B1(n6984), 
        .B2(i_data_bus[766]), .ZN(n6946) );
  ND2D1BWP30P140LVT U10200 ( .A1(n6947), .A2(n6946), .ZN(N1673) );
  AOI22D1BWP30P140LVT U10201 ( .A1(n6987), .A2(i_data_bus[701]), .B1(n6986), 
        .B2(i_data_bus[669]), .ZN(n6949) );
  AOI22D1BWP30P140LVT U10202 ( .A1(n6985), .A2(i_data_bus[733]), .B1(n6984), 
        .B2(i_data_bus[765]), .ZN(n6948) );
  ND2D1BWP30P140LVT U10203 ( .A1(n6949), .A2(n6948), .ZN(N1672) );
  AOI22D1BWP30P140LVT U10204 ( .A1(n6987), .A2(i_data_bus[698]), .B1(n6986), 
        .B2(i_data_bus[666]), .ZN(n6951) );
  AOI22D1BWP30P140LVT U10205 ( .A1(n6985), .A2(i_data_bus[730]), .B1(n6984), 
        .B2(i_data_bus[762]), .ZN(n6950) );
  ND2D1BWP30P140LVT U10206 ( .A1(n6951), .A2(n6950), .ZN(N1669) );
  AOI22D1BWP30P140LVT U10207 ( .A1(n6985), .A2(i_data_bus[729]), .B1(n6986), 
        .B2(i_data_bus[665]), .ZN(n6953) );
  AOI22D1BWP30P140LVT U10208 ( .A1(n6987), .A2(i_data_bus[697]), .B1(n6984), 
        .B2(i_data_bus[761]), .ZN(n6952) );
  ND2D1BWP30P140LVT U10209 ( .A1(n6953), .A2(n6952), .ZN(N1668) );
  AOI22D1BWP30P140LVT U10210 ( .A1(n6987), .A2(i_data_bus[689]), .B1(n6986), 
        .B2(i_data_bus[657]), .ZN(n6955) );
  AOI22D1BWP30P140LVT U10211 ( .A1(n6985), .A2(i_data_bus[721]), .B1(n6984), 
        .B2(i_data_bus[753]), .ZN(n6954) );
  ND2D1BWP30P140LVT U10212 ( .A1(n6955), .A2(n6954), .ZN(N1660) );
  AOI22D1BWP30P140LVT U10213 ( .A1(n6987), .A2(i_data_bus[683]), .B1(n6986), 
        .B2(i_data_bus[651]), .ZN(n6957) );
  AOI22D1BWP30P140LVT U10214 ( .A1(n6985), .A2(i_data_bus[715]), .B1(n6984), 
        .B2(i_data_bus[747]), .ZN(n6956) );
  ND2D1BWP30P140LVT U10215 ( .A1(n6957), .A2(n6956), .ZN(N1654) );
  AOI22D1BWP30P140LVT U10216 ( .A1(n6987), .A2(i_data_bus[680]), .B1(n6986), 
        .B2(i_data_bus[648]), .ZN(n6959) );
  AOI22D1BWP30P140LVT U10217 ( .A1(n6985), .A2(i_data_bus[712]), .B1(n6984), 
        .B2(i_data_bus[744]), .ZN(n6958) );
  ND2D1BWP30P140LVT U10218 ( .A1(n6959), .A2(n6958), .ZN(N1651) );
  AOI22D1BWP30P140LVT U10219 ( .A1(n6987), .A2(i_data_bus[679]), .B1(n6986), 
        .B2(i_data_bus[647]), .ZN(n6961) );
  AOI22D1BWP30P140LVT U10220 ( .A1(n6985), .A2(i_data_bus[711]), .B1(n6984), 
        .B2(i_data_bus[743]), .ZN(n6960) );
  ND2D1BWP30P140LVT U10221 ( .A1(n6961), .A2(n6960), .ZN(N1650) );
  AOI22D1BWP30P140LVT U10222 ( .A1(n6987), .A2(i_data_bus[676]), .B1(n6986), 
        .B2(i_data_bus[644]), .ZN(n6963) );
  AOI22D1BWP30P140LVT U10223 ( .A1(n6985), .A2(i_data_bus[708]), .B1(n6984), 
        .B2(i_data_bus[740]), .ZN(n6962) );
  ND2D1BWP30P140LVT U10224 ( .A1(n6963), .A2(n6962), .ZN(N1647) );
  AOI22D1BWP30P140LVT U10225 ( .A1(n6985), .A2(i_data_bus[706]), .B1(n6986), 
        .B2(i_data_bus[642]), .ZN(n6965) );
  AOI22D1BWP30P140LVT U10226 ( .A1(n6987), .A2(i_data_bus[674]), .B1(n6984), 
        .B2(i_data_bus[738]), .ZN(n6964) );
  ND2D1BWP30P140LVT U10227 ( .A1(n6965), .A2(n6964), .ZN(N1645) );
  AOI22D1BWP30P140LVT U10228 ( .A1(n6985), .A2(i_data_bus[705]), .B1(n6986), 
        .B2(i_data_bus[641]), .ZN(n6967) );
  AOI22D1BWP30P140LVT U10229 ( .A1(n6987), .A2(i_data_bus[673]), .B1(n6984), 
        .B2(i_data_bus[737]), .ZN(n6966) );
  ND2D1BWP30P140LVT U10230 ( .A1(n6967), .A2(n6966), .ZN(N1644) );
  AOI22D1BWP30P140LVT U10231 ( .A1(n6987), .A2(i_data_bus[699]), .B1(n6984), 
        .B2(i_data_bus[763]), .ZN(n6969) );
  AOI22D1BWP30P140LVT U10232 ( .A1(n6985), .A2(i_data_bus[731]), .B1(n6986), 
        .B2(i_data_bus[667]), .ZN(n6968) );
  ND2D1BWP30P140LVT U10233 ( .A1(n6969), .A2(n6968), .ZN(N1670) );
  AOI22D1BWP30P140LVT U10234 ( .A1(n6987), .A2(i_data_bus[696]), .B1(n6984), 
        .B2(i_data_bus[760]), .ZN(n6971) );
  AOI22D1BWP30P140LVT U10235 ( .A1(n6985), .A2(i_data_bus[728]), .B1(n6986), 
        .B2(i_data_bus[664]), .ZN(n6970) );
  ND2D1BWP30P140LVT U10236 ( .A1(n6971), .A2(n6970), .ZN(N1667) );
  AOI22D1BWP30P140LVT U10237 ( .A1(n6985), .A2(i_data_bus[726]), .B1(n6984), 
        .B2(i_data_bus[758]), .ZN(n6973) );
  AOI22D1BWP30P140LVT U10238 ( .A1(n6987), .A2(i_data_bus[694]), .B1(n6986), 
        .B2(i_data_bus[662]), .ZN(n6972) );
  ND2D1BWP30P140LVT U10239 ( .A1(n6973), .A2(n6972), .ZN(N1665) );
  AOI22D1BWP30P140LVT U10240 ( .A1(n6985), .A2(i_data_bus[719]), .B1(n6984), 
        .B2(i_data_bus[751]), .ZN(n6975) );
  AOI22D1BWP30P140LVT U10241 ( .A1(n6987), .A2(i_data_bus[687]), .B1(n6986), 
        .B2(i_data_bus[655]), .ZN(n6974) );
  ND2D1BWP30P140LVT U10242 ( .A1(n6975), .A2(n6974), .ZN(N1658) );
  AOI22D1BWP30P140LVT U10243 ( .A1(n6985), .A2(i_data_bus[718]), .B1(n6984), 
        .B2(i_data_bus[750]), .ZN(n6977) );
  AOI22D1BWP30P140LVT U10244 ( .A1(n6987), .A2(i_data_bus[686]), .B1(n6986), 
        .B2(i_data_bus[654]), .ZN(n6976) );
  ND2D1BWP30P140LVT U10245 ( .A1(n6977), .A2(n6976), .ZN(N1657) );
  AOI22D1BWP30P140LVT U10246 ( .A1(n6985), .A2(i_data_bus[717]), .B1(n6984), 
        .B2(i_data_bus[749]), .ZN(n6979) );
  AOI22D1BWP30P140LVT U10247 ( .A1(n6987), .A2(i_data_bus[685]), .B1(n6986), 
        .B2(i_data_bus[653]), .ZN(n6978) );
  ND2D1BWP30P140LVT U10248 ( .A1(n6979), .A2(n6978), .ZN(N1656) );
  AOI22D1BWP30P140LVT U10249 ( .A1(n6987), .A2(i_data_bus[684]), .B1(n6984), 
        .B2(i_data_bus[748]), .ZN(n6981) );
  AOI22D1BWP30P140LVT U10250 ( .A1(n6985), .A2(i_data_bus[716]), .B1(n6986), 
        .B2(i_data_bus[652]), .ZN(n6980) );
  ND2D1BWP30P140LVT U10251 ( .A1(n6981), .A2(n6980), .ZN(N1655) );
  AOI22D1BWP30P140LVT U10252 ( .A1(n6985), .A2(i_data_bus[713]), .B1(n6984), 
        .B2(i_data_bus[745]), .ZN(n6983) );
  AOI22D1BWP30P140LVT U10253 ( .A1(n6987), .A2(i_data_bus[681]), .B1(n6986), 
        .B2(i_data_bus[649]), .ZN(n6982) );
  ND2D1BWP30P140LVT U10254 ( .A1(n6983), .A2(n6982), .ZN(N1652) );
  AOI22D1BWP30P140LVT U10255 ( .A1(n6985), .A2(i_data_bus[707]), .B1(n6984), 
        .B2(i_data_bus[739]), .ZN(n6989) );
  AOI22D1BWP30P140LVT U10256 ( .A1(n6987), .A2(i_data_bus[675]), .B1(n6986), 
        .B2(i_data_bus[643]), .ZN(n6988) );
  ND2D1BWP30P140LVT U10257 ( .A1(n6989), .A2(n6988), .ZN(N1646) );
  NR3D0P7BWP30P140LVT U10258 ( .A1(i_cmd[207]), .A2(i_cmd[223]), .A3(
        i_cmd[215]), .ZN(n10915) );
  NR4D1BWP30P140LVT U10259 ( .A1(i_cmd[207]), .A2(n7179), .A3(n10918), .A4(
        n6990), .ZN(n7333) );
  AOI22D1BWP30P140LVT U10260 ( .A1(i_data_bus[781]), .A2(n7335), .B1(
        i_data_bus[877]), .B2(n7333), .ZN(n6992) );
  INR4D1BWP30P140LVT U10261 ( .A1(i_cmd[215]), .B1(i_cmd[199]), .B2(n7181), 
        .B3(n10916), .ZN(n7334) );
  AOI22D1BWP30P140LVT U10262 ( .A1(i_data_bus[845]), .A2(n7334), .B1(
        i_data_bus[813]), .B2(n7336), .ZN(n6991) );
  ND2D1BWP30P140LVT U10263 ( .A1(n6992), .A2(n6991), .ZN(N11030) );
  AOI22D1BWP30P140LVT U10264 ( .A1(i_data_bus[772]), .A2(n7335), .B1(
        i_data_bus[836]), .B2(n7334), .ZN(n6994) );
  AOI22D1BWP30P140LVT U10265 ( .A1(i_data_bus[868]), .A2(n7333), .B1(
        i_data_bus[804]), .B2(n7336), .ZN(n6993) );
  ND2D1BWP30P140LVT U10266 ( .A1(n6994), .A2(n6993), .ZN(N11021) );
  NR3D0P7BWP30P140LVT U10267 ( .A1(i_cmd[213]), .A2(i_cmd[221]), .A3(
        i_cmd[205]), .ZN(n10973) );
  INVD1BWP30P140LVT U10268 ( .I(i_cmd[205]), .ZN(n6995) );
  AOI22D1BWP30P140LVT U10269 ( .A1(i_data_bus[794]), .A2(n7325), .B1(
        i_data_bus[826]), .B2(n7326), .ZN(n6999) );
  INVD1BWP30P140LVT U10270 ( .I(i_cmd[221]), .ZN(n6997) );
  INR4D1BWP30P140LVT U10271 ( .A1(i_cmd[213]), .B1(i_cmd[197]), .B2(n7181), 
        .B3(n10977), .ZN(n7324) );
  NR4D1BWP30P140LVT U10272 ( .A1(i_cmd[205]), .A2(n6997), .A3(n7179), .A4(
        n6996), .ZN(n7323) );
  AOI22D1BWP30P140LVT U10273 ( .A1(i_data_bus[858]), .A2(n7324), .B1(
        i_data_bus[890]), .B2(n7323), .ZN(n6998) );
  ND2D1BWP30P140LVT U10274 ( .A1(n6999), .A2(n6998), .ZN(N8319) );
  AOI22D1BWP30P140LVT U10275 ( .A1(i_data_bus[784]), .A2(n7325), .B1(
        i_data_bus[848]), .B2(n7324), .ZN(n7001) );
  AOI22D1BWP30P140LVT U10276 ( .A1(i_data_bus[816]), .A2(n7326), .B1(
        i_data_bus[880]), .B2(n7323), .ZN(n7000) );
  ND2D1BWP30P140LVT U10277 ( .A1(n7001), .A2(n7000), .ZN(N8309) );
  AOI22D1BWP30P140LVT U10278 ( .A1(i_data_bus[776]), .A2(n7325), .B1(
        i_data_bus[808]), .B2(n7326), .ZN(n7003) );
  AOI22D1BWP30P140LVT U10279 ( .A1(i_data_bus[840]), .A2(n7324), .B1(
        i_data_bus[872]), .B2(n7323), .ZN(n7002) );
  ND2D1BWP30P140LVT U10280 ( .A1(n7003), .A2(n7002), .ZN(N8301) );
  AOI22D1BWP30P140LVT U10281 ( .A1(i_data_bus[795]), .A2(n7335), .B1(
        i_data_bus[859]), .B2(n7334), .ZN(n7005) );
  AOI22D1BWP30P140LVT U10282 ( .A1(i_data_bus[827]), .A2(n7336), .B1(
        i_data_bus[891]), .B2(n7333), .ZN(n7004) );
  ND2D1BWP30P140LVT U10283 ( .A1(n7005), .A2(n7004), .ZN(N11044) );
  AOI22D1BWP30P140LVT U10284 ( .A1(i_data_bus[789]), .A2(n7335), .B1(
        i_data_bus[853]), .B2(n7334), .ZN(n7007) );
  AOI22D1BWP30P140LVT U10285 ( .A1(i_data_bus[821]), .A2(n7336), .B1(
        i_data_bus[885]), .B2(n7333), .ZN(n7006) );
  ND2D1BWP30P140LVT U10286 ( .A1(n7007), .A2(n7006), .ZN(N11038) );
  AOI22D1BWP30P140LVT U10287 ( .A1(i_data_bus[799]), .A2(n7325), .B1(
        i_data_bus[863]), .B2(n7324), .ZN(n7009) );
  AOI22D1BWP30P140LVT U10288 ( .A1(i_data_bus[895]), .A2(n7323), .B1(
        i_data_bus[831]), .B2(n7326), .ZN(n7008) );
  ND2D1BWP30P140LVT U10289 ( .A1(n7009), .A2(n7008), .ZN(N8324) );
  AOI22D1BWP30P140LVT U10290 ( .A1(i_data_bus[797]), .A2(n7325), .B1(
        i_data_bus[861]), .B2(n7324), .ZN(n7011) );
  AOI22D1BWP30P140LVT U10291 ( .A1(i_data_bus[893]), .A2(n7323), .B1(
        i_data_bus[829]), .B2(n7326), .ZN(n7010) );
  ND2D1BWP30P140LVT U10292 ( .A1(n7011), .A2(n7010), .ZN(N8322) );
  AOI22D1BWP30P140LVT U10293 ( .A1(i_data_bus[785]), .A2(n7325), .B1(
        i_data_bus[849]), .B2(n7324), .ZN(n7013) );
  AOI22D1BWP30P140LVT U10294 ( .A1(i_data_bus[881]), .A2(n7323), .B1(
        i_data_bus[817]), .B2(n7326), .ZN(n7012) );
  ND2D1BWP30P140LVT U10295 ( .A1(n7013), .A2(n7012), .ZN(N8310) );
  AOI22D1BWP30P140LVT U10296 ( .A1(i_data_bus[779]), .A2(n7325), .B1(
        i_data_bus[875]), .B2(n7323), .ZN(n7015) );
  AOI22D1BWP30P140LVT U10297 ( .A1(i_data_bus[843]), .A2(n7324), .B1(
        i_data_bus[811]), .B2(n7326), .ZN(n7014) );
  ND2D1BWP30P140LVT U10298 ( .A1(n7015), .A2(n7014), .ZN(N8304) );
  AOI22D1BWP30P140LVT U10299 ( .A1(i_data_bus[778]), .A2(n7325), .B1(
        i_data_bus[842]), .B2(n7324), .ZN(n7017) );
  AOI22D1BWP30P140LVT U10300 ( .A1(i_data_bus[874]), .A2(n7323), .B1(
        i_data_bus[810]), .B2(n7326), .ZN(n7016) );
  ND2D1BWP30P140LVT U10301 ( .A1(n7017), .A2(n7016), .ZN(N8303) );
  AOI22D1BWP30P140LVT U10302 ( .A1(i_data_bus[772]), .A2(n7325), .B1(
        i_data_bus[836]), .B2(n7324), .ZN(n7019) );
  AOI22D1BWP30P140LVT U10303 ( .A1(i_data_bus[868]), .A2(n7323), .B1(
        i_data_bus[804]), .B2(n7326), .ZN(n7018) );
  ND2D1BWP30P140LVT U10304 ( .A1(n7019), .A2(n7018), .ZN(N8297) );
  NR3D0P7BWP30P140LVT U10305 ( .A1(i_cmd[210]), .A2(i_cmd[202]), .A3(
        i_cmd[218]), .ZN(n11096) );
  ND2D1BWP30P140LVT U10306 ( .A1(n11096), .A2(i_cmd[194]), .ZN(n11098) );
  OR2D1BWP30P140LVT U10307 ( .A1(i_cmd[202]), .A2(i_cmd[218]), .Z(n11100) );
  INR4D1BWP30P140LVT U10308 ( .A1(i_cmd[210]), .B1(i_cmd[194]), .B2(n7181), 
        .B3(n11100), .ZN(n7302) );
  AOI22D1BWP30P140LVT U10309 ( .A1(i_data_bus[787]), .A2(n7303), .B1(
        i_data_bus[851]), .B2(n7302), .ZN(n7022) );
  INR4D1BWP30P140LVT U10310 ( .A1(i_cmd[218]), .B1(i_cmd[202]), .B2(n7179), 
        .B3(n7020), .ZN(n7301) );
  INR4D1BWP30P140LVT U10311 ( .A1(i_cmd[202]), .B1(i_cmd[218]), .B2(n7183), 
        .B3(n7020), .ZN(n7304) );
  AOI22D1BWP30P140LVT U10312 ( .A1(i_data_bus[883]), .A2(n7301), .B1(
        i_data_bus[819]), .B2(n7304), .ZN(n7021) );
  ND2D1BWP30P140LVT U10313 ( .A1(n7022), .A2(n7021), .ZN(N4610) );
  AOI22D1BWP30P140LVT U10314 ( .A1(i_data_bus[781]), .A2(n7303), .B1(
        i_data_bus[877]), .B2(n7301), .ZN(n7024) );
  AOI22D1BWP30P140LVT U10315 ( .A1(i_data_bus[845]), .A2(n7302), .B1(
        i_data_bus[813]), .B2(n7304), .ZN(n7023) );
  ND2D1BWP30P140LVT U10316 ( .A1(n7024), .A2(n7023), .ZN(N4604) );
  NR3D0P7BWP30P140LVT U10317 ( .A1(i_cmd[201]), .A2(i_cmd[217]), .A3(
        i_cmd[209]), .ZN(n11120) );
  OR2D1BWP30P140LVT U10318 ( .A1(i_cmd[201]), .A2(i_cmd[217]), .Z(n11124) );
  INR4D1BWP30P140LVT U10319 ( .A1(i_cmd[209]), .B1(i_cmd[193]), .B2(n7181), 
        .B3(n11124), .ZN(n7351) );
  AOI22D1BWP30P140LVT U10320 ( .A1(i_data_bus[789]), .A2(n7353), .B1(
        i_data_bus[853]), .B2(n7351), .ZN(n7027) );
  INR4D1BWP30P140LVT U10321 ( .A1(i_cmd[201]), .B1(i_cmd[217]), .B2(n7183), 
        .B3(n7025), .ZN(n7352) );
  INR4D1BWP30P140LVT U10322 ( .A1(i_cmd[217]), .B1(i_cmd[201]), .B2(n7179), 
        .B3(n7025), .ZN(n7354) );
  AOI22D1BWP30P140LVT U10323 ( .A1(i_data_bus[821]), .A2(n7352), .B1(
        i_data_bus[885]), .B2(n7354), .ZN(n7026) );
  ND2D1BWP30P140LVT U10324 ( .A1(n7027), .A2(n7026), .ZN(N2866) );
  AOI22D1BWP30P140LVT U10325 ( .A1(i_data_bus[786]), .A2(n7353), .B1(
        i_data_bus[850]), .B2(n7351), .ZN(n7029) );
  AOI22D1BWP30P140LVT U10326 ( .A1(i_data_bus[818]), .A2(n7352), .B1(
        i_data_bus[882]), .B2(n7354), .ZN(n7028) );
  ND2D1BWP30P140LVT U10327 ( .A1(n7029), .A2(n7028), .ZN(N2863) );
  AOI22D1BWP30P140LVT U10328 ( .A1(i_data_bus[776]), .A2(n7353), .B1(
        i_data_bus[808]), .B2(n7352), .ZN(n7031) );
  AOI22D1BWP30P140LVT U10329 ( .A1(i_data_bus[840]), .A2(n7351), .B1(
        i_data_bus[872]), .B2(n7354), .ZN(n7030) );
  ND2D1BWP30P140LVT U10330 ( .A1(n7031), .A2(n7030), .ZN(N2853) );
  AOI22D1BWP30P140LVT U10331 ( .A1(i_data_bus[770]), .A2(n7353), .B1(
        i_data_bus[802]), .B2(n7352), .ZN(n7033) );
  AOI22D1BWP30P140LVT U10332 ( .A1(i_data_bus[834]), .A2(n7351), .B1(
        i_data_bus[866]), .B2(n7354), .ZN(n7032) );
  ND2D1BWP30P140LVT U10333 ( .A1(n7033), .A2(n7032), .ZN(N2847) );
  AOI22D1BWP30P140LVT U10334 ( .A1(i_data_bus[797]), .A2(n7353), .B1(
        i_data_bus[861]), .B2(n7351), .ZN(n7035) );
  AOI22D1BWP30P140LVT U10335 ( .A1(i_data_bus[893]), .A2(n7354), .B1(
        i_data_bus[829]), .B2(n7352), .ZN(n7034) );
  ND2D1BWP30P140LVT U10336 ( .A1(n7035), .A2(n7034), .ZN(N2874) );
  AOI22D1BWP30P140LVT U10337 ( .A1(i_data_bus[781]), .A2(n7353), .B1(
        i_data_bus[877]), .B2(n7354), .ZN(n7037) );
  AOI22D1BWP30P140LVT U10338 ( .A1(i_data_bus[845]), .A2(n7351), .B1(
        i_data_bus[813]), .B2(n7352), .ZN(n7036) );
  ND2D1BWP30P140LVT U10339 ( .A1(n7037), .A2(n7036), .ZN(N2858) );
  AOI22D1BWP30P140LVT U10340 ( .A1(i_data_bus[772]), .A2(n7353), .B1(
        i_data_bus[836]), .B2(n7351), .ZN(n7039) );
  AOI22D1BWP30P140LVT U10341 ( .A1(i_data_bus[868]), .A2(n7354), .B1(
        i_data_bus[804]), .B2(n7352), .ZN(n7038) );
  ND2D1BWP30P140LVT U10342 ( .A1(n7039), .A2(n7038), .ZN(N2849) );
  AOI22D1BWP30P140LVT U10343 ( .A1(i_data_bus[793]), .A2(n7325), .B1(
        i_data_bus[825]), .B2(n7326), .ZN(n7041) );
  AOI22D1BWP30P140LVT U10344 ( .A1(i_data_bus[889]), .A2(n7323), .B1(
        i_data_bus[857]), .B2(n7324), .ZN(n7040) );
  ND2D1BWP30P140LVT U10345 ( .A1(n7041), .A2(n7040), .ZN(N8318) );
  AOI22D1BWP30P140LVT U10346 ( .A1(i_data_bus[786]), .A2(n7325), .B1(
        i_data_bus[882]), .B2(n7323), .ZN(n7043) );
  AOI22D1BWP30P140LVT U10347 ( .A1(i_data_bus[818]), .A2(n7326), .B1(
        i_data_bus[850]), .B2(n7324), .ZN(n7042) );
  ND2D1BWP30P140LVT U10348 ( .A1(n7043), .A2(n7042), .ZN(N8311) );
  AOI22D1BWP30P140LVT U10349 ( .A1(i_data_bus[775]), .A2(n7325), .B1(
        i_data_bus[807]), .B2(n7326), .ZN(n7045) );
  AOI22D1BWP30P140LVT U10350 ( .A1(i_data_bus[871]), .A2(n7323), .B1(
        i_data_bus[839]), .B2(n7324), .ZN(n7044) );
  ND2D1BWP30P140LVT U10351 ( .A1(n7045), .A2(n7044), .ZN(N8300) );
  AOI22D1BWP30P140LVT U10352 ( .A1(i_data_bus[771]), .A2(n7325), .B1(
        i_data_bus[803]), .B2(n7326), .ZN(n7047) );
  AOI22D1BWP30P140LVT U10353 ( .A1(i_data_bus[867]), .A2(n7323), .B1(
        i_data_bus[835]), .B2(n7324), .ZN(n7046) );
  ND2D1BWP30P140LVT U10354 ( .A1(n7047), .A2(n7046), .ZN(N8296) );
  AOI22D1BWP30P140LVT U10355 ( .A1(i_data_bus[796]), .A2(n7335), .B1(
        i_data_bus[828]), .B2(n7336), .ZN(n7049) );
  AOI22D1BWP30P140LVT U10356 ( .A1(i_data_bus[892]), .A2(n7333), .B1(
        i_data_bus[860]), .B2(n7334), .ZN(n7048) );
  ND2D1BWP30P140LVT U10357 ( .A1(n7049), .A2(n7048), .ZN(N11045) );
  AOI22D1BWP30P140LVT U10358 ( .A1(i_data_bus[793]), .A2(n7335), .B1(
        i_data_bus[889]), .B2(n7333), .ZN(n7051) );
  AOI22D1BWP30P140LVT U10359 ( .A1(i_data_bus[825]), .A2(n7336), .B1(
        i_data_bus[857]), .B2(n7334), .ZN(n7050) );
  ND2D1BWP30P140LVT U10360 ( .A1(n7051), .A2(n7050), .ZN(N11042) );
  AOI22D1BWP30P140LVT U10361 ( .A1(i_data_bus[792]), .A2(n7335), .B1(
        i_data_bus[824]), .B2(n7336), .ZN(n7053) );
  AOI22D1BWP30P140LVT U10362 ( .A1(i_data_bus[888]), .A2(n7333), .B1(
        i_data_bus[856]), .B2(n7334), .ZN(n7052) );
  ND2D1BWP30P140LVT U10363 ( .A1(n7053), .A2(n7052), .ZN(N11041) );
  AOI22D1BWP30P140LVT U10364 ( .A1(i_data_bus[786]), .A2(n7335), .B1(
        i_data_bus[818]), .B2(n7336), .ZN(n7055) );
  AOI22D1BWP30P140LVT U10365 ( .A1(i_data_bus[882]), .A2(n7333), .B1(
        i_data_bus[850]), .B2(n7334), .ZN(n7054) );
  ND2D1BWP30P140LVT U10366 ( .A1(n7055), .A2(n7054), .ZN(N11035) );
  AOI22D1BWP30P140LVT U10367 ( .A1(i_data_bus[771]), .A2(n7335), .B1(
        i_data_bus[803]), .B2(n7336), .ZN(n7057) );
  AOI22D1BWP30P140LVT U10368 ( .A1(i_data_bus[867]), .A2(n7333), .B1(
        i_data_bus[835]), .B2(n7334), .ZN(n7056) );
  ND2D1BWP30P140LVT U10369 ( .A1(n7057), .A2(n7056), .ZN(N11020) );
  AOI22D1BWP30P140LVT U10370 ( .A1(i_data_bus[796]), .A2(n7303), .B1(
        i_data_bus[828]), .B2(n7304), .ZN(n7059) );
  AOI22D1BWP30P140LVT U10371 ( .A1(i_data_bus[892]), .A2(n7301), .B1(
        i_data_bus[860]), .B2(n7302), .ZN(n7058) );
  ND2D1BWP30P140LVT U10372 ( .A1(n7059), .A2(n7058), .ZN(N4619) );
  AOI22D1BWP30P140LVT U10373 ( .A1(i_data_bus[795]), .A2(n7303), .B1(
        i_data_bus[827]), .B2(n7304), .ZN(n7061) );
  AOI22D1BWP30P140LVT U10374 ( .A1(i_data_bus[891]), .A2(n7301), .B1(
        i_data_bus[859]), .B2(n7302), .ZN(n7060) );
  ND2D1BWP30P140LVT U10375 ( .A1(n7061), .A2(n7060), .ZN(N4618) );
  AOI22D1BWP30P140LVT U10376 ( .A1(i_data_bus[792]), .A2(n7303), .B1(
        i_data_bus[824]), .B2(n7304), .ZN(n7063) );
  AOI22D1BWP30P140LVT U10377 ( .A1(i_data_bus[888]), .A2(n7301), .B1(
        i_data_bus[856]), .B2(n7302), .ZN(n7062) );
  ND2D1BWP30P140LVT U10378 ( .A1(n7063), .A2(n7062), .ZN(N4615) );
  AOI22D1BWP30P140LVT U10379 ( .A1(i_data_bus[788]), .A2(n7303), .B1(
        i_data_bus[884]), .B2(n7301), .ZN(n7065) );
  AOI22D1BWP30P140LVT U10380 ( .A1(i_data_bus[820]), .A2(n7304), .B1(
        i_data_bus[852]), .B2(n7302), .ZN(n7064) );
  ND2D1BWP30P140LVT U10381 ( .A1(n7065), .A2(n7064), .ZN(N4611) );
  AOI22D1BWP30P140LVT U10382 ( .A1(i_data_bus[778]), .A2(n7303), .B1(
        i_data_bus[874]), .B2(n7301), .ZN(n7067) );
  AOI22D1BWP30P140LVT U10383 ( .A1(i_data_bus[810]), .A2(n7304), .B1(
        i_data_bus[842]), .B2(n7302), .ZN(n7066) );
  ND2D1BWP30P140LVT U10384 ( .A1(n7067), .A2(n7066), .ZN(N4601) );
  AOI22D1BWP30P140LVT U10385 ( .A1(i_data_bus[771]), .A2(n7303), .B1(
        i_data_bus[867]), .B2(n7301), .ZN(n7069) );
  AOI22D1BWP30P140LVT U10386 ( .A1(i_data_bus[803]), .A2(n7304), .B1(
        i_data_bus[835]), .B2(n7302), .ZN(n7068) );
  ND2D1BWP30P140LVT U10387 ( .A1(n7069), .A2(n7068), .ZN(N4594) );
  AOI22D1BWP30P140LVT U10388 ( .A1(i_data_bus[799]), .A2(n7353), .B1(
        i_data_bus[895]), .B2(n7354), .ZN(n7071) );
  AOI22D1BWP30P140LVT U10389 ( .A1(i_data_bus[831]), .A2(n7352), .B1(
        i_data_bus[863]), .B2(n7351), .ZN(n7070) );
  ND2D1BWP30P140LVT U10390 ( .A1(n7071), .A2(n7070), .ZN(N2876) );
  AOI22D1BWP30P140LVT U10391 ( .A1(i_data_bus[793]), .A2(n7353), .B1(
        i_data_bus[825]), .B2(n7352), .ZN(n7073) );
  AOI22D1BWP30P140LVT U10392 ( .A1(i_data_bus[889]), .A2(n7354), .B1(
        i_data_bus[857]), .B2(n7351), .ZN(n7072) );
  ND2D1BWP30P140LVT U10393 ( .A1(n7073), .A2(n7072), .ZN(N2870) );
  AOI22D1BWP30P140LVT U10394 ( .A1(i_data_bus[792]), .A2(n7353), .B1(
        i_data_bus[824]), .B2(n7352), .ZN(n7075) );
  AOI22D1BWP30P140LVT U10395 ( .A1(i_data_bus[888]), .A2(n7354), .B1(
        i_data_bus[856]), .B2(n7351), .ZN(n7074) );
  ND2D1BWP30P140LVT U10396 ( .A1(n7075), .A2(n7074), .ZN(N2869) );
  AOI22D1BWP30P140LVT U10397 ( .A1(i_data_bus[776]), .A2(n7365), .B1(
        i_data_bus[808]), .B2(n7366), .ZN(n7081) );
  AOI22D1BWP30P140LVT U10398 ( .A1(i_data_bus[840]), .A2(n7364), .B1(
        i_data_bus[872]), .B2(n7363), .ZN(n7080) );
  ND2D1BWP30P140LVT U10399 ( .A1(n7081), .A2(n7080), .ZN(N10047) );
  AOI22D1BWP30P140LVT U10400 ( .A1(i_data_bus[791]), .A2(n7365), .B1(
        i_data_bus[855]), .B2(n7364), .ZN(n7083) );
  AOI22D1BWP30P140LVT U10401 ( .A1(i_data_bus[887]), .A2(n7363), .B1(
        i_data_bus[823]), .B2(n7366), .ZN(n7082) );
  ND2D1BWP30P140LVT U10402 ( .A1(n7083), .A2(n7082), .ZN(N10062) );
  AOI22D1BWP30P140LVT U10403 ( .A1(i_data_bus[779]), .A2(n7365), .B1(
        i_data_bus[843]), .B2(n7364), .ZN(n7085) );
  AOI22D1BWP30P140LVT U10404 ( .A1(i_data_bus[875]), .A2(n7363), .B1(
        i_data_bus[811]), .B2(n7366), .ZN(n7084) );
  ND2D1BWP30P140LVT U10405 ( .A1(n7085), .A2(n7084), .ZN(N10050) );
  AOI22D1BWP30P140LVT U10406 ( .A1(i_data_bus[789]), .A2(n7365), .B1(
        i_data_bus[885]), .B2(n7363), .ZN(n7087) );
  AOI22D1BWP30P140LVT U10407 ( .A1(i_data_bus[853]), .A2(n7364), .B1(
        i_data_bus[821]), .B2(n7366), .ZN(n7086) );
  ND2D1BWP30P140LVT U10408 ( .A1(n7087), .A2(n7086), .ZN(N10060) );
  AOI22D1BWP30P140LVT U10409 ( .A1(i_data_bus[786]), .A2(n7365), .B1(
        i_data_bus[850]), .B2(n7364), .ZN(n7089) );
  AOI22D1BWP30P140LVT U10410 ( .A1(i_data_bus[818]), .A2(n7366), .B1(
        i_data_bus[882]), .B2(n7363), .ZN(n7088) );
  ND2D1BWP30P140LVT U10411 ( .A1(n7089), .A2(n7088), .ZN(N10057) );
  AOI22D1BWP30P140LVT U10412 ( .A1(i_data_bus[772]), .A2(n7365), .B1(
        i_data_bus[868]), .B2(n7363), .ZN(n7091) );
  AOI22D1BWP30P140LVT U10413 ( .A1(i_data_bus[836]), .A2(n7364), .B1(
        i_data_bus[804]), .B2(n7366), .ZN(n7090) );
  ND2D1BWP30P140LVT U10414 ( .A1(n7091), .A2(n7090), .ZN(N10043) );
  AOI22D1BWP30P140LVT U10415 ( .A1(i_data_bus[778]), .A2(n7365), .B1(
        i_data_bus[874]), .B2(n7363), .ZN(n7093) );
  AOI22D1BWP30P140LVT U10416 ( .A1(i_data_bus[810]), .A2(n7366), .B1(
        i_data_bus[842]), .B2(n7364), .ZN(n7092) );
  ND2D1BWP30P140LVT U10417 ( .A1(n7093), .A2(n7092), .ZN(N10049) );
  AOI22D1BWP30P140LVT U10418 ( .A1(i_data_bus[775]), .A2(n7365), .B1(
        i_data_bus[871]), .B2(n7363), .ZN(n7095) );
  AOI22D1BWP30P140LVT U10419 ( .A1(i_data_bus[807]), .A2(n7366), .B1(
        i_data_bus[839]), .B2(n7364), .ZN(n7094) );
  ND2D1BWP30P140LVT U10420 ( .A1(n7095), .A2(n7094), .ZN(N10046) );
  AOI22D1BWP30P140LVT U10421 ( .A1(i_data_bus[895]), .A2(n7333), .B1(
        i_data_bus[863]), .B2(n7334), .ZN(n7097) );
  AOI22D1BWP30P140LVT U10422 ( .A1(i_data_bus[799]), .A2(n7335), .B1(
        i_data_bus[831]), .B2(n7336), .ZN(n7096) );
  ND2D1BWP30P140LVT U10423 ( .A1(n7097), .A2(n7096), .ZN(N11048) );
  AOI22D1BWP30P140LVT U10424 ( .A1(i_data_bus[820]), .A2(n7336), .B1(
        i_data_bus[852]), .B2(n7334), .ZN(n7099) );
  AOI22D1BWP30P140LVT U10425 ( .A1(i_data_bus[788]), .A2(n7335), .B1(
        i_data_bus[884]), .B2(n7333), .ZN(n7098) );
  ND2D1BWP30P140LVT U10426 ( .A1(n7099), .A2(n7098), .ZN(N11037) );
  AOI22D1BWP30P140LVT U10427 ( .A1(i_data_bus[883]), .A2(n7333), .B1(
        i_data_bus[819]), .B2(n7336), .ZN(n7101) );
  AOI22D1BWP30P140LVT U10428 ( .A1(i_data_bus[787]), .A2(n7335), .B1(
        i_data_bus[851]), .B2(n7334), .ZN(n7100) );
  ND2D1BWP30P140LVT U10429 ( .A1(n7101), .A2(n7100), .ZN(N11036) );
  AOI22D1BWP30P140LVT U10430 ( .A1(i_data_bus[843]), .A2(n7334), .B1(
        i_data_bus[811]), .B2(n7336), .ZN(n7103) );
  AOI22D1BWP30P140LVT U10431 ( .A1(i_data_bus[779]), .A2(n7335), .B1(
        i_data_bus[875]), .B2(n7333), .ZN(n7102) );
  ND2D1BWP30P140LVT U10432 ( .A1(n7103), .A2(n7102), .ZN(N11028) );
  AOI22D1BWP30P140LVT U10433 ( .A1(i_data_bus[810]), .A2(n7336), .B1(
        i_data_bus[842]), .B2(n7334), .ZN(n7105) );
  AOI22D1BWP30P140LVT U10434 ( .A1(i_data_bus[778]), .A2(n7335), .B1(
        i_data_bus[874]), .B2(n7333), .ZN(n7104) );
  ND2D1BWP30P140LVT U10435 ( .A1(n7105), .A2(n7104), .ZN(N11027) );
  AOI22D1BWP30P140LVT U10436 ( .A1(i_data_bus[840]), .A2(n7334), .B1(
        i_data_bus[808]), .B2(n7336), .ZN(n7107) );
  AOI22D1BWP30P140LVT U10437 ( .A1(i_data_bus[776]), .A2(n7335), .B1(
        i_data_bus[872]), .B2(n7333), .ZN(n7106) );
  ND2D1BWP30P140LVT U10438 ( .A1(n7107), .A2(n7106), .ZN(N11025) );
  AOI22D1BWP30P140LVT U10439 ( .A1(i_data_bus[871]), .A2(n7333), .B1(
        i_data_bus[807]), .B2(n7336), .ZN(n7109) );
  AOI22D1BWP30P140LVT U10440 ( .A1(i_data_bus[775]), .A2(n7335), .B1(
        i_data_bus[839]), .B2(n7334), .ZN(n7108) );
  ND2D1BWP30P140LVT U10441 ( .A1(n7109), .A2(n7108), .ZN(N11024) );
  AOI22D1BWP30P140LVT U10442 ( .A1(i_data_bus[870]), .A2(n7333), .B1(
        i_data_bus[806]), .B2(n7336), .ZN(n7111) );
  AOI22D1BWP30P140LVT U10443 ( .A1(i_data_bus[774]), .A2(n7335), .B1(
        i_data_bus[838]), .B2(n7334), .ZN(n7110) );
  ND2D1BWP30P140LVT U10444 ( .A1(n7111), .A2(n7110), .ZN(N11023) );
  AOI22D1BWP30P140LVT U10445 ( .A1(i_data_bus[802]), .A2(n7336), .B1(
        i_data_bus[866]), .B2(n7333), .ZN(n7113) );
  AOI22D1BWP30P140LVT U10446 ( .A1(i_data_bus[770]), .A2(n7335), .B1(
        i_data_bus[834]), .B2(n7334), .ZN(n7112) );
  ND2D1BWP30P140LVT U10447 ( .A1(n7113), .A2(n7112), .ZN(N11019) );
  AOI22D1BWP30P140LVT U10448 ( .A1(i_data_bus[895]), .A2(n7301), .B1(
        i_data_bus[831]), .B2(n7304), .ZN(n7115) );
  AOI22D1BWP30P140LVT U10449 ( .A1(i_data_bus[799]), .A2(n7303), .B1(
        i_data_bus[863]), .B2(n7302), .ZN(n7114) );
  ND2D1BWP30P140LVT U10450 ( .A1(n7115), .A2(n7114), .ZN(N4622) );
  AOI22D1BWP30P140LVT U10451 ( .A1(i_data_bus[893]), .A2(n7301), .B1(
        i_data_bus[829]), .B2(n7304), .ZN(n7117) );
  AOI22D1BWP30P140LVT U10452 ( .A1(i_data_bus[797]), .A2(n7303), .B1(
        i_data_bus[861]), .B2(n7302), .ZN(n7116) );
  ND2D1BWP30P140LVT U10453 ( .A1(n7117), .A2(n7116), .ZN(N4620) );
  AOI22D1BWP30P140LVT U10454 ( .A1(i_data_bus[825]), .A2(n7304), .B1(
        i_data_bus[857]), .B2(n7302), .ZN(n7119) );
  AOI22D1BWP30P140LVT U10455 ( .A1(i_data_bus[793]), .A2(n7303), .B1(
        i_data_bus[889]), .B2(n7301), .ZN(n7118) );
  ND2D1BWP30P140LVT U10456 ( .A1(n7119), .A2(n7118), .ZN(N4616) );
  AOI22D1BWP30P140LVT U10457 ( .A1(i_data_bus[821]), .A2(n7304), .B1(
        i_data_bus[885]), .B2(n7301), .ZN(n7121) );
  AOI22D1BWP30P140LVT U10458 ( .A1(i_data_bus[789]), .A2(n7303), .B1(
        i_data_bus[853]), .B2(n7302), .ZN(n7120) );
  ND2D1BWP30P140LVT U10459 ( .A1(n7121), .A2(n7120), .ZN(N4612) );
  AOI22D1BWP30P140LVT U10460 ( .A1(i_data_bus[818]), .A2(n7304), .B1(
        i_data_bus[882]), .B2(n7301), .ZN(n7123) );
  AOI22D1BWP30P140LVT U10461 ( .A1(i_data_bus[786]), .A2(n7303), .B1(
        i_data_bus[850]), .B2(n7302), .ZN(n7122) );
  ND2D1BWP30P140LVT U10462 ( .A1(n7123), .A2(n7122), .ZN(N4609) );
  AOI22D1BWP30P140LVT U10463 ( .A1(i_data_bus[843]), .A2(n7302), .B1(
        i_data_bus[811]), .B2(n7304), .ZN(n7125) );
  AOI22D1BWP30P140LVT U10464 ( .A1(i_data_bus[779]), .A2(n7303), .B1(
        i_data_bus[875]), .B2(n7301), .ZN(n7124) );
  ND2D1BWP30P140LVT U10465 ( .A1(n7125), .A2(n7124), .ZN(N4602) );
  AOI22D1BWP30P140LVT U10466 ( .A1(i_data_bus[808]), .A2(n7304), .B1(
        i_data_bus[872]), .B2(n7301), .ZN(n7127) );
  AOI22D1BWP30P140LVT U10467 ( .A1(i_data_bus[776]), .A2(n7303), .B1(
        i_data_bus[840]), .B2(n7302), .ZN(n7126) );
  ND2D1BWP30P140LVT U10468 ( .A1(n7127), .A2(n7126), .ZN(N4599) );
  AOI22D1BWP30P140LVT U10469 ( .A1(i_data_bus[871]), .A2(n7301), .B1(
        i_data_bus[807]), .B2(n7304), .ZN(n7129) );
  AOI22D1BWP30P140LVT U10470 ( .A1(i_data_bus[775]), .A2(n7303), .B1(
        i_data_bus[839]), .B2(n7302), .ZN(n7128) );
  ND2D1BWP30P140LVT U10471 ( .A1(n7129), .A2(n7128), .ZN(N4598) );
  AOI22D1BWP30P140LVT U10472 ( .A1(i_data_bus[868]), .A2(n7301), .B1(
        i_data_bus[804]), .B2(n7304), .ZN(n7131) );
  AOI22D1BWP30P140LVT U10473 ( .A1(i_data_bus[772]), .A2(n7303), .B1(
        i_data_bus[836]), .B2(n7302), .ZN(n7130) );
  ND2D1BWP30P140LVT U10474 ( .A1(n7131), .A2(n7130), .ZN(N4595) );
  AOI22D1BWP30P140LVT U10475 ( .A1(i_data_bus[802]), .A2(n7304), .B1(
        i_data_bus[866]), .B2(n7301), .ZN(n7133) );
  AOI22D1BWP30P140LVT U10476 ( .A1(i_data_bus[770]), .A2(n7303), .B1(
        i_data_bus[834]), .B2(n7302), .ZN(n7132) );
  ND2D1BWP30P140LVT U10477 ( .A1(n7133), .A2(n7132), .ZN(N4593) );
  AOI22D1BWP30P140LVT U10478 ( .A1(i_data_bus[891]), .A2(n7323), .B1(
        i_data_bus[859]), .B2(n7324), .ZN(n7135) );
  AOI22D1BWP30P140LVT U10479 ( .A1(i_data_bus[795]), .A2(n7325), .B1(
        i_data_bus[827]), .B2(n7326), .ZN(n7134) );
  ND2D1BWP30P140LVT U10480 ( .A1(n7135), .A2(n7134), .ZN(N8320) );
  AOI22D1BWP30P140LVT U10481 ( .A1(i_data_bus[888]), .A2(n7323), .B1(
        i_data_bus[856]), .B2(n7324), .ZN(n7137) );
  AOI22D1BWP30P140LVT U10482 ( .A1(i_data_bus[792]), .A2(n7325), .B1(
        i_data_bus[824]), .B2(n7326), .ZN(n7136) );
  ND2D1BWP30P140LVT U10483 ( .A1(n7137), .A2(n7136), .ZN(N8317) );
  AOI22D1BWP30P140LVT U10484 ( .A1(i_data_bus[853]), .A2(n7324), .B1(
        i_data_bus[821]), .B2(n7326), .ZN(n7139) );
  AOI22D1BWP30P140LVT U10485 ( .A1(i_data_bus[789]), .A2(n7325), .B1(
        i_data_bus[885]), .B2(n7323), .ZN(n7138) );
  ND2D1BWP30P140LVT U10486 ( .A1(n7139), .A2(n7138), .ZN(N8314) );
  AOI22D1BWP30P140LVT U10487 ( .A1(i_data_bus[870]), .A2(n7323), .B1(
        i_data_bus[806]), .B2(n7326), .ZN(n7141) );
  AOI22D1BWP30P140LVT U10488 ( .A1(i_data_bus[774]), .A2(n7325), .B1(
        i_data_bus[838]), .B2(n7324), .ZN(n7140) );
  ND2D1BWP30P140LVT U10489 ( .A1(n7141), .A2(n7140), .ZN(N8299) );
  AOI22D1BWP30P140LVT U10490 ( .A1(i_data_bus[802]), .A2(n7326), .B1(
        i_data_bus[866]), .B2(n7323), .ZN(n7143) );
  AOI22D1BWP30P140LVT U10491 ( .A1(i_data_bus[770]), .A2(n7325), .B1(
        i_data_bus[834]), .B2(n7324), .ZN(n7142) );
  ND2D1BWP30P140LVT U10492 ( .A1(n7143), .A2(n7142), .ZN(N8295) );
  AOI22D1BWP30P140LVT U10493 ( .A1(i_data_bus[827]), .A2(n7352), .B1(
        i_data_bus[891]), .B2(n7354), .ZN(n7145) );
  AOI22D1BWP30P140LVT U10494 ( .A1(i_data_bus[795]), .A2(n7353), .B1(
        i_data_bus[859]), .B2(n7351), .ZN(n7144) );
  ND2D1BWP30P140LVT U10495 ( .A1(n7145), .A2(n7144), .ZN(N2872) );
  AOI22D1BWP30P140LVT U10496 ( .A1(i_data_bus[883]), .A2(n7354), .B1(
        i_data_bus[819]), .B2(n7352), .ZN(n7147) );
  AOI22D1BWP30P140LVT U10497 ( .A1(i_data_bus[787]), .A2(n7353), .B1(
        i_data_bus[851]), .B2(n7351), .ZN(n7146) );
  ND2D1BWP30P140LVT U10498 ( .A1(n7147), .A2(n7146), .ZN(N2864) );
  AOI22D1BWP30P140LVT U10499 ( .A1(i_data_bus[844]), .A2(n7351), .B1(
        i_data_bus[812]), .B2(n7352), .ZN(n7149) );
  AOI22D1BWP30P140LVT U10500 ( .A1(i_data_bus[780]), .A2(n7353), .B1(
        i_data_bus[876]), .B2(n7354), .ZN(n7148) );
  ND2D1BWP30P140LVT U10501 ( .A1(n7149), .A2(n7148), .ZN(N2857) );
  AOI22D1BWP30P140LVT U10502 ( .A1(i_data_bus[875]), .A2(n7354), .B1(
        i_data_bus[811]), .B2(n7352), .ZN(n7151) );
  AOI22D1BWP30P140LVT U10503 ( .A1(i_data_bus[779]), .A2(n7353), .B1(
        i_data_bus[843]), .B2(n7351), .ZN(n7150) );
  ND2D1BWP30P140LVT U10504 ( .A1(n7151), .A2(n7150), .ZN(N2856) );
  AOI22D1BWP30P140LVT U10505 ( .A1(i_data_bus[810]), .A2(n7352), .B1(
        i_data_bus[842]), .B2(n7351), .ZN(n7153) );
  AOI22D1BWP30P140LVT U10506 ( .A1(i_data_bus[778]), .A2(n7353), .B1(
        i_data_bus[874]), .B2(n7354), .ZN(n7152) );
  ND2D1BWP30P140LVT U10507 ( .A1(n7153), .A2(n7152), .ZN(N2855) );
  AOI22D1BWP30P140LVT U10508 ( .A1(i_data_bus[871]), .A2(n7354), .B1(
        i_data_bus[839]), .B2(n7351), .ZN(n7155) );
  AOI22D1BWP30P140LVT U10509 ( .A1(i_data_bus[775]), .A2(n7353), .B1(
        i_data_bus[807]), .B2(n7352), .ZN(n7154) );
  ND2D1BWP30P140LVT U10510 ( .A1(n7155), .A2(n7154), .ZN(N2852) );
  AOI22D1BWP30P140LVT U10511 ( .A1(i_data_bus[867]), .A2(n7354), .B1(
        i_data_bus[835]), .B2(n7351), .ZN(n7157) );
  AOI22D1BWP30P140LVT U10512 ( .A1(i_data_bus[771]), .A2(n7353), .B1(
        i_data_bus[803]), .B2(n7352), .ZN(n7156) );
  ND2D1BWP30P140LVT U10513 ( .A1(n7157), .A2(n7156), .ZN(N2848) );
  AOI22D1BWP30P140LVT U10514 ( .A1(i_data_bus[832]), .A2(n7351), .B1(
        i_data_bus[800]), .B2(n7352), .ZN(n7159) );
  AOI22D1BWP30P140LVT U10515 ( .A1(i_data_bus[768]), .A2(n7353), .B1(
        i_data_bus[864]), .B2(n7354), .ZN(n7158) );
  ND2D1BWP30P140LVT U10516 ( .A1(n7159), .A2(n7158), .ZN(N2845) );
  AOI22D1BWP30P140LVT U10517 ( .A1(i_data_bus[827]), .A2(n7366), .B1(
        i_data_bus[891]), .B2(n7363), .ZN(n7161) );
  AOI22D1BWP30P140LVT U10518 ( .A1(i_data_bus[795]), .A2(n7365), .B1(
        i_data_bus[859]), .B2(n7364), .ZN(n7160) );
  ND2D1BWP30P140LVT U10519 ( .A1(n7161), .A2(n7160), .ZN(N10066) );
  AOI22D1BWP30P140LVT U10520 ( .A1(i_data_bus[825]), .A2(n7366), .B1(
        i_data_bus[889]), .B2(n7363), .ZN(n7163) );
  AOI22D1BWP30P140LVT U10521 ( .A1(i_data_bus[793]), .A2(n7365), .B1(
        i_data_bus[857]), .B2(n7364), .ZN(n7162) );
  ND2D1BWP30P140LVT U10522 ( .A1(n7163), .A2(n7162), .ZN(N10064) );
  AOI22D1BWP30P140LVT U10523 ( .A1(i_data_bus[870]), .A2(n7363), .B1(
        i_data_bus[806]), .B2(n7366), .ZN(n7165) );
  AOI22D1BWP30P140LVT U10524 ( .A1(i_data_bus[774]), .A2(n7365), .B1(
        i_data_bus[838]), .B2(n7364), .ZN(n7164) );
  ND2D1BWP30P140LVT U10525 ( .A1(n7165), .A2(n7164), .ZN(N10045) );
  AOI22D1BWP30P140LVT U10526 ( .A1(i_data_bus[803]), .A2(n7366), .B1(
        i_data_bus[867]), .B2(n7363), .ZN(n7167) );
  AOI22D1BWP30P140LVT U10527 ( .A1(i_data_bus[771]), .A2(n7365), .B1(
        i_data_bus[835]), .B2(n7364), .ZN(n7166) );
  ND2D1BWP30P140LVT U10528 ( .A1(n7167), .A2(n7166), .ZN(N10042) );
  AOI22D1BWP30P140LVT U10529 ( .A1(i_data_bus[831]), .A2(n7366), .B1(
        i_data_bus[863]), .B2(n7364), .ZN(n7169) );
  AOI22D1BWP30P140LVT U10530 ( .A1(i_data_bus[799]), .A2(n7365), .B1(
        i_data_bus[895]), .B2(n7363), .ZN(n7168) );
  ND2D1BWP30P140LVT U10531 ( .A1(n7169), .A2(n7168), .ZN(N10070) );
  AOI22D1BWP30P140LVT U10532 ( .A1(i_data_bus[856]), .A2(n7364), .B1(
        i_data_bus[824]), .B2(n7366), .ZN(n7171) );
  AOI22D1BWP30P140LVT U10533 ( .A1(i_data_bus[792]), .A2(n7365), .B1(
        i_data_bus[888]), .B2(n7363), .ZN(n7170) );
  ND2D1BWP30P140LVT U10534 ( .A1(n7171), .A2(n7170), .ZN(N10063) );
  AOI22D1BWP30P140LVT U10535 ( .A1(i_data_bus[820]), .A2(n7366), .B1(
        i_data_bus[852]), .B2(n7364), .ZN(n7173) );
  AOI22D1BWP30P140LVT U10536 ( .A1(i_data_bus[788]), .A2(n7365), .B1(
        i_data_bus[884]), .B2(n7363), .ZN(n7172) );
  ND2D1BWP30P140LVT U10537 ( .A1(n7173), .A2(n7172), .ZN(N10059) );
  AOI22D1BWP30P140LVT U10538 ( .A1(i_data_bus[844]), .A2(n7364), .B1(
        i_data_bus[812]), .B2(n7366), .ZN(n7175) );
  AOI22D1BWP30P140LVT U10539 ( .A1(i_data_bus[780]), .A2(n7365), .B1(
        i_data_bus[876]), .B2(n7363), .ZN(n7174) );
  ND2D1BWP30P140LVT U10540 ( .A1(n7175), .A2(n7174), .ZN(N10051) );
  AOI22D1BWP30P140LVT U10541 ( .A1(i_data_bus[834]), .A2(n7364), .B1(
        i_data_bus[802]), .B2(n7366), .ZN(n7177) );
  AOI22D1BWP30P140LVT U10542 ( .A1(i_data_bus[770]), .A2(n7365), .B1(
        i_data_bus[866]), .B2(n7363), .ZN(n7176) );
  ND2D1BWP30P140LVT U10543 ( .A1(n7177), .A2(n7176), .ZN(N10041) );
  NR3D0P7BWP30P140LVT U10544 ( .A1(i_cmd[208]), .A2(i_cmd[200]), .A3(
        i_cmd[216]), .ZN(n11151) );
  INVD1BWP30P140LVT U10545 ( .I(i_cmd[216]), .ZN(n7180) );
  NR4D1BWP30P140LVT U10546 ( .A1(i_cmd[200]), .A2(n7180), .A3(n7182), .A4(
        n7179), .ZN(n7422) );
  AOI22D1BWP30P140LVT U10547 ( .A1(i_data_bus[768]), .A2(n7424), .B1(
        i_data_bus[864]), .B2(n7422), .ZN(n7186) );
  INVD1BWP30P140LVT U10548 ( .I(i_cmd[200]), .ZN(n7184) );
  INR4D1BWP30P140LVT U10549 ( .A1(i_cmd[208]), .B1(i_cmd[192]), .B2(n7181), 
        .B3(n11155), .ZN(n7425) );
  AOI22D1BWP30P140LVT U10550 ( .A1(i_data_bus[832]), .A2(n7425), .B1(
        i_data_bus[800]), .B2(n7423), .ZN(n7185) );
  ND2D1BWP30P140LVT U10551 ( .A1(n7186), .A2(n7185), .ZN(N1863) );
  AOI22D1BWP30P140LVT U10552 ( .A1(n7424), .A2(i_data_bus[788]), .B1(n7422), 
        .B2(i_data_bus[884]), .ZN(n7188) );
  AOI22D1BWP30P140LVT U10553 ( .A1(n7425), .A2(i_data_bus[852]), .B1(n7423), 
        .B2(i_data_bus[820]), .ZN(n7187) );
  ND2D1BWP30P140LVT U10554 ( .A1(n7188), .A2(n7187), .ZN(N1883) );
  AOI22D1BWP30P140LVT U10555 ( .A1(n7424), .A2(i_data_bus[782]), .B1(n7422), 
        .B2(i_data_bus[878]), .ZN(n7190) );
  AOI22D1BWP30P140LVT U10556 ( .A1(n7425), .A2(i_data_bus[846]), .B1(n7423), 
        .B2(i_data_bus[814]), .ZN(n7189) );
  ND2D1BWP30P140LVT U10557 ( .A1(n7190), .A2(n7189), .ZN(N1877) );
  AOI22D1BWP30P140LVT U10558 ( .A1(n7424), .A2(i_data_bus[781]), .B1(n7422), 
        .B2(i_data_bus[877]), .ZN(n7192) );
  AOI22D1BWP30P140LVT U10559 ( .A1(n7425), .A2(i_data_bus[845]), .B1(n7423), 
        .B2(i_data_bus[813]), .ZN(n7191) );
  ND2D1BWP30P140LVT U10560 ( .A1(n7192), .A2(n7191), .ZN(N1876) );
  AOI22D1BWP30P140LVT U10561 ( .A1(n7424), .A2(i_data_bus[780]), .B1(n7422), 
        .B2(i_data_bus[876]), .ZN(n7194) );
  AOI22D1BWP30P140LVT U10562 ( .A1(n7425), .A2(i_data_bus[844]), .B1(n7423), 
        .B2(i_data_bus[812]), .ZN(n7193) );
  ND2D1BWP30P140LVT U10563 ( .A1(n7194), .A2(n7193), .ZN(N1875) );
  AOI22D1BWP30P140LVT U10564 ( .A1(n7424), .A2(i_data_bus[777]), .B1(n7422), 
        .B2(i_data_bus[873]), .ZN(n7196) );
  AOI22D1BWP30P140LVT U10565 ( .A1(n7425), .A2(i_data_bus[841]), .B1(n7423), 
        .B2(i_data_bus[809]), .ZN(n7195) );
  ND2D1BWP30P140LVT U10566 ( .A1(n7196), .A2(n7195), .ZN(N1872) );
  AOI22D1BWP30P140LVT U10567 ( .A1(i_data_bus[873]), .A2(n7333), .B1(
        i_data_bus[777]), .B2(n7335), .ZN(n7198) );
  AOI22D1BWP30P140LVT U10568 ( .A1(i_data_bus[841]), .A2(n7334), .B1(
        i_data_bus[809]), .B2(n7336), .ZN(n7197) );
  ND2D1BWP30P140LVT U10569 ( .A1(n7198), .A2(n7197), .ZN(N11026) );
  AOI22D1BWP30P140LVT U10570 ( .A1(i_data_bus[822]), .A2(n7326), .B1(
        i_data_bus[790]), .B2(n7325), .ZN(n7200) );
  AOI22D1BWP30P140LVT U10571 ( .A1(i_data_bus[854]), .A2(n7324), .B1(
        i_data_bus[886]), .B2(n7323), .ZN(n7199) );
  ND2D1BWP30P140LVT U10572 ( .A1(n7200), .A2(n7199), .ZN(N8315) );
  AOI22D1BWP30P140LVT U10573 ( .A1(i_data_bus[846]), .A2(n7324), .B1(
        i_data_bus[782]), .B2(n7325), .ZN(n7202) );
  AOI22D1BWP30P140LVT U10574 ( .A1(i_data_bus[814]), .A2(n7326), .B1(
        i_data_bus[878]), .B2(n7323), .ZN(n7201) );
  ND2D1BWP30P140LVT U10575 ( .A1(n7202), .A2(n7201), .ZN(N8307) );
  AOI22D1BWP30P140LVT U10576 ( .A1(i_data_bus[845]), .A2(n7324), .B1(
        i_data_bus[781]), .B2(n7325), .ZN(n7204) );
  AOI22D1BWP30P140LVT U10577 ( .A1(i_data_bus[813]), .A2(n7326), .B1(
        i_data_bus[877]), .B2(n7323), .ZN(n7203) );
  ND2D1BWP30P140LVT U10578 ( .A1(n7204), .A2(n7203), .ZN(N8306) );
  AOI22D1BWP30P140LVT U10579 ( .A1(i_data_bus[809]), .A2(n7326), .B1(
        i_data_bus[777]), .B2(n7325), .ZN(n7206) );
  AOI22D1BWP30P140LVT U10580 ( .A1(i_data_bus[841]), .A2(n7324), .B1(
        i_data_bus[873]), .B2(n7323), .ZN(n7205) );
  ND2D1BWP30P140LVT U10581 ( .A1(n7206), .A2(n7205), .ZN(N8302) );
  AOI22D1BWP30P140LVT U10582 ( .A1(i_data_bus[844]), .A2(n7334), .B1(
        i_data_bus[780]), .B2(n7335), .ZN(n7208) );
  AOI22D1BWP30P140LVT U10583 ( .A1(i_data_bus[812]), .A2(n7336), .B1(
        i_data_bus[876]), .B2(n7333), .ZN(n7207) );
  ND2D1BWP30P140LVT U10584 ( .A1(n7208), .A2(n7207), .ZN(N11029) );
  AOI22D1BWP30P140LVT U10585 ( .A1(i_data_bus[832]), .A2(n7334), .B1(
        i_data_bus[768]), .B2(n7335), .ZN(n7210) );
  AOI22D1BWP30P140LVT U10586 ( .A1(i_data_bus[800]), .A2(n7336), .B1(
        i_data_bus[864]), .B2(n7333), .ZN(n7209) );
  ND2D1BWP30P140LVT U10587 ( .A1(n7210), .A2(n7209), .ZN(N11017) );
  AOI22D1BWP30P140LVT U10588 ( .A1(i_data_bus[860]), .A2(n7324), .B1(
        i_data_bus[796]), .B2(n7325), .ZN(n7212) );
  AOI22D1BWP30P140LVT U10589 ( .A1(i_data_bus[892]), .A2(n7323), .B1(
        i_data_bus[828]), .B2(n7326), .ZN(n7211) );
  ND2D1BWP30P140LVT U10590 ( .A1(n7212), .A2(n7211), .ZN(N8321) );
  AOI22D1BWP30P140LVT U10591 ( .A1(i_data_bus[890]), .A2(n7301), .B1(
        i_data_bus[794]), .B2(n7303), .ZN(n7214) );
  AOI22D1BWP30P140LVT U10592 ( .A1(i_data_bus[858]), .A2(n7302), .B1(
        i_data_bus[826]), .B2(n7304), .ZN(n7213) );
  ND2D1BWP30P140LVT U10593 ( .A1(n7214), .A2(n7213), .ZN(N4617) );
  AOI22D1BWP30P140LVT U10594 ( .A1(i_data_bus[820]), .A2(n7352), .B1(
        i_data_bus[788]), .B2(n7353), .ZN(n7216) );
  AOI22D1BWP30P140LVT U10595 ( .A1(i_data_bus[852]), .A2(n7351), .B1(
        i_data_bus[884]), .B2(n7354), .ZN(n7215) );
  ND2D1BWP30P140LVT U10596 ( .A1(n7216), .A2(n7215), .ZN(N2865) );
  AOI22D1BWP30P140LVT U10597 ( .A1(i_data_bus[809]), .A2(n7352), .B1(
        i_data_bus[777]), .B2(n7353), .ZN(n7218) );
  AOI22D1BWP30P140LVT U10598 ( .A1(i_data_bus[841]), .A2(n7351), .B1(
        i_data_bus[873]), .B2(n7354), .ZN(n7217) );
  ND2D1BWP30P140LVT U10599 ( .A1(n7218), .A2(n7217), .ZN(N2854) );
  AOI22D1BWP30P140LVT U10600 ( .A1(i_data_bus[833]), .A2(n7302), .B1(
        i_data_bus[769]), .B2(n7303), .ZN(n7220) );
  AOI22D1BWP30P140LVT U10601 ( .A1(i_data_bus[801]), .A2(n7304), .B1(
        i_data_bus[865]), .B2(n7301), .ZN(n7219) );
  ND2D1BWP30P140LVT U10602 ( .A1(n7220), .A2(n7219), .ZN(N4592) );
  AOI22D1BWP30P140LVT U10603 ( .A1(i_data_bus[854]), .A2(n7351), .B1(
        i_data_bus[790]), .B2(n7353), .ZN(n7222) );
  AOI22D1BWP30P140LVT U10604 ( .A1(i_data_bus[886]), .A2(n7354), .B1(
        i_data_bus[822]), .B2(n7352), .ZN(n7221) );
  ND2D1BWP30P140LVT U10605 ( .A1(n7222), .A2(n7221), .ZN(N2867) );
  AOI22D1BWP30P140LVT U10606 ( .A1(i_data_bus[829]), .A2(n7336), .B1(
        i_data_bus[797]), .B2(n7335), .ZN(n7224) );
  AOI22D1BWP30P140LVT U10607 ( .A1(i_data_bus[893]), .A2(n7333), .B1(
        i_data_bus[861]), .B2(n7334), .ZN(n7223) );
  ND2D1BWP30P140LVT U10608 ( .A1(n7224), .A2(n7223), .ZN(N11046) );
  AOI22D1BWP30P140LVT U10609 ( .A1(i_data_bus[823]), .A2(n7336), .B1(
        i_data_bus[791]), .B2(n7335), .ZN(n7226) );
  AOI22D1BWP30P140LVT U10610 ( .A1(i_data_bus[887]), .A2(n7333), .B1(
        i_data_bus[855]), .B2(n7334), .ZN(n7225) );
  ND2D1BWP30P140LVT U10611 ( .A1(n7226), .A2(n7225), .ZN(N11040) );
  AOI22D1BWP30P140LVT U10612 ( .A1(i_data_bus[817]), .A2(n7336), .B1(
        i_data_bus[785]), .B2(n7335), .ZN(n7228) );
  AOI22D1BWP30P140LVT U10613 ( .A1(i_data_bus[881]), .A2(n7333), .B1(
        i_data_bus[849]), .B2(n7334), .ZN(n7227) );
  ND2D1BWP30P140LVT U10614 ( .A1(n7228), .A2(n7227), .ZN(N11034) );
  AOI22D1BWP30P140LVT U10615 ( .A1(i_data_bus[869]), .A2(n7333), .B1(
        i_data_bus[773]), .B2(n7335), .ZN(n7230) );
  AOI22D1BWP30P140LVT U10616 ( .A1(i_data_bus[805]), .A2(n7336), .B1(
        i_data_bus[837]), .B2(n7334), .ZN(n7229) );
  ND2D1BWP30P140LVT U10617 ( .A1(n7230), .A2(n7229), .ZN(N11022) );
  AOI22D1BWP30P140LVT U10618 ( .A1(i_data_bus[830]), .A2(n7352), .B1(
        i_data_bus[798]), .B2(n7353), .ZN(n7232) );
  AOI22D1BWP30P140LVT U10619 ( .A1(i_data_bus[894]), .A2(n7354), .B1(
        i_data_bus[862]), .B2(n7351), .ZN(n7231) );
  ND2D1BWP30P140LVT U10620 ( .A1(n7232), .A2(n7231), .ZN(N2875) );
  AOI22D1BWP30P140LVT U10621 ( .A1(i_data_bus[887]), .A2(n7354), .B1(
        i_data_bus[791]), .B2(n7353), .ZN(n7234) );
  AOI22D1BWP30P140LVT U10622 ( .A1(i_data_bus[823]), .A2(n7352), .B1(
        i_data_bus[855]), .B2(n7351), .ZN(n7233) );
  ND2D1BWP30P140LVT U10623 ( .A1(n7234), .A2(n7233), .ZN(N2868) );
  AOI22D1BWP30P140LVT U10624 ( .A1(i_data_bus[817]), .A2(n7352), .B1(
        i_data_bus[785]), .B2(n7353), .ZN(n7236) );
  AOI22D1BWP30P140LVT U10625 ( .A1(i_data_bus[881]), .A2(n7354), .B1(
        i_data_bus[849]), .B2(n7351), .ZN(n7235) );
  ND2D1BWP30P140LVT U10626 ( .A1(n7236), .A2(n7235), .ZN(N2862) );
  AOI22D1BWP30P140LVT U10627 ( .A1(i_data_bus[878]), .A2(n7354), .B1(
        i_data_bus[782]), .B2(n7353), .ZN(n7238) );
  AOI22D1BWP30P140LVT U10628 ( .A1(i_data_bus[814]), .A2(n7352), .B1(
        i_data_bus[846]), .B2(n7351), .ZN(n7237) );
  ND2D1BWP30P140LVT U10629 ( .A1(n7238), .A2(n7237), .ZN(N2859) );
  AOI22D1BWP30P140LVT U10630 ( .A1(i_data_bus[823]), .A2(n7304), .B1(
        i_data_bus[791]), .B2(n7303), .ZN(n7240) );
  AOI22D1BWP30P140LVT U10631 ( .A1(i_data_bus[887]), .A2(n7301), .B1(
        i_data_bus[855]), .B2(n7302), .ZN(n7239) );
  ND2D1BWP30P140LVT U10632 ( .A1(n7240), .A2(n7239), .ZN(N4614) );
  AOI22D1BWP30P140LVT U10633 ( .A1(i_data_bus[879]), .A2(n7301), .B1(
        i_data_bus[783]), .B2(n7303), .ZN(n7242) );
  AOI22D1BWP30P140LVT U10634 ( .A1(i_data_bus[815]), .A2(n7304), .B1(
        i_data_bus[847]), .B2(n7302), .ZN(n7241) );
  ND2D1BWP30P140LVT U10635 ( .A1(n7242), .A2(n7241), .ZN(N4606) );
  AOI22D1BWP30P140LVT U10636 ( .A1(i_data_bus[806]), .A2(n7304), .B1(
        i_data_bus[774]), .B2(n7303), .ZN(n7244) );
  AOI22D1BWP30P140LVT U10637 ( .A1(i_data_bus[870]), .A2(n7301), .B1(
        i_data_bus[838]), .B2(n7302), .ZN(n7243) );
  ND2D1BWP30P140LVT U10638 ( .A1(n7244), .A2(n7243), .ZN(N4597) );
  AOI22D1BWP30P140LVT U10639 ( .A1(i_data_bus[860]), .A2(n7364), .B1(
        i_data_bus[796]), .B2(n7365), .ZN(n7246) );
  AOI22D1BWP30P140LVT U10640 ( .A1(i_data_bus[892]), .A2(n7363), .B1(
        i_data_bus[828]), .B2(n7366), .ZN(n7245) );
  ND2D1BWP30P140LVT U10641 ( .A1(n7246), .A2(n7245), .ZN(N10067) );
  AOI22D1BWP30P140LVT U10642 ( .A1(i_data_bus[830]), .A2(n7366), .B1(
        i_data_bus[798]), .B2(n7365), .ZN(n7248) );
  AOI22D1BWP30P140LVT U10643 ( .A1(i_data_bus[894]), .A2(n7363), .B1(
        i_data_bus[862]), .B2(n7364), .ZN(n7247) );
  ND2D1BWP30P140LVT U10644 ( .A1(n7248), .A2(n7247), .ZN(N10069) );
  AOI22D1BWP30P140LVT U10645 ( .A1(i_data_bus[829]), .A2(n7366), .B1(
        i_data_bus[797]), .B2(n7365), .ZN(n7250) );
  AOI22D1BWP30P140LVT U10646 ( .A1(i_data_bus[893]), .A2(n7363), .B1(
        i_data_bus[861]), .B2(n7364), .ZN(n7249) );
  ND2D1BWP30P140LVT U10647 ( .A1(n7250), .A2(n7249), .ZN(N10068) );
  AOI22D1BWP30P140LVT U10648 ( .A1(i_data_bus[880]), .A2(n7363), .B1(
        i_data_bus[784]), .B2(n7365), .ZN(n7252) );
  AOI22D1BWP30P140LVT U10649 ( .A1(i_data_bus[816]), .A2(n7366), .B1(
        i_data_bus[848]), .B2(n7364), .ZN(n7251) );
  ND2D1BWP30P140LVT U10650 ( .A1(n7252), .A2(n7251), .ZN(N10055) );
  AOI22D1BWP30P140LVT U10651 ( .A1(i_data_bus[878]), .A2(n7363), .B1(
        i_data_bus[782]), .B2(n7365), .ZN(n7254) );
  AOI22D1BWP30P140LVT U10652 ( .A1(i_data_bus[814]), .A2(n7366), .B1(
        i_data_bus[846]), .B2(n7364), .ZN(n7253) );
  ND2D1BWP30P140LVT U10653 ( .A1(n7254), .A2(n7253), .ZN(N10053) );
  AOI22D1BWP30P140LVT U10654 ( .A1(i_data_bus[869]), .A2(n7363), .B1(
        i_data_bus[773]), .B2(n7365), .ZN(n7256) );
  AOI22D1BWP30P140LVT U10655 ( .A1(i_data_bus[805]), .A2(n7366), .B1(
        i_data_bus[837]), .B2(n7364), .ZN(n7255) );
  ND2D1BWP30P140LVT U10656 ( .A1(n7256), .A2(n7255), .ZN(N10044) );
  AOI22D1BWP30P140LVT U10657 ( .A1(i_data_bus[822]), .A2(n7366), .B1(
        i_data_bus[790]), .B2(n7365), .ZN(n7258) );
  AOI22D1BWP30P140LVT U10658 ( .A1(i_data_bus[854]), .A2(n7364), .B1(
        i_data_bus[886]), .B2(n7363), .ZN(n7257) );
  ND2D1BWP30P140LVT U10659 ( .A1(n7258), .A2(n7257), .ZN(N10061) );
  AOI22D1BWP30P140LVT U10660 ( .A1(i_data_bus[847]), .A2(n7364), .B1(
        i_data_bus[783]), .B2(n7365), .ZN(n7260) );
  AOI22D1BWP30P140LVT U10661 ( .A1(i_data_bus[815]), .A2(n7366), .B1(
        i_data_bus[879]), .B2(n7363), .ZN(n7259) );
  ND2D1BWP30P140LVT U10662 ( .A1(n7260), .A2(n7259), .ZN(N10054) );
  AOI22D1BWP30P140LVT U10663 ( .A1(i_data_bus[813]), .A2(n7366), .B1(
        i_data_bus[781]), .B2(n7365), .ZN(n7262) );
  AOI22D1BWP30P140LVT U10664 ( .A1(i_data_bus[845]), .A2(n7364), .B1(
        i_data_bus[877]), .B2(n7363), .ZN(n7261) );
  ND2D1BWP30P140LVT U10665 ( .A1(n7262), .A2(n7261), .ZN(N10052) );
  AOI22D1BWP30P140LVT U10666 ( .A1(i_data_bus[833]), .A2(n7364), .B1(
        i_data_bus[769]), .B2(n7365), .ZN(n7264) );
  AOI22D1BWP30P140LVT U10667 ( .A1(i_data_bus[801]), .A2(n7366), .B1(
        i_data_bus[865]), .B2(n7363), .ZN(n7263) );
  ND2D1BWP30P140LVT U10668 ( .A1(n7264), .A2(n7263), .ZN(N10040) );
  AOI22D1BWP30P140LVT U10669 ( .A1(i_data_bus[800]), .A2(n7366), .B1(
        i_data_bus[768]), .B2(n7365), .ZN(n7266) );
  AOI22D1BWP30P140LVT U10670 ( .A1(i_data_bus[832]), .A2(n7364), .B1(
        i_data_bus[864]), .B2(n7363), .ZN(n7265) );
  ND2D1BWP30P140LVT U10671 ( .A1(n7266), .A2(n7265), .ZN(N10039) );
  AOI22D1BWP30P140LVT U10672 ( .A1(n7425), .A2(i_data_bus[863]), .B1(n7423), 
        .B2(i_data_bus[831]), .ZN(n7268) );
  AOI22D1BWP30P140LVT U10673 ( .A1(n7424), .A2(i_data_bus[799]), .B1(n7422), 
        .B2(i_data_bus[895]), .ZN(n7267) );
  ND2D1BWP30P140LVT U10674 ( .A1(n7268), .A2(n7267), .ZN(N1894) );
  AOI22D1BWP30P140LVT U10675 ( .A1(n7425), .A2(i_data_bus[856]), .B1(n7423), 
        .B2(i_data_bus[824]), .ZN(n7270) );
  AOI22D1BWP30P140LVT U10676 ( .A1(n7424), .A2(i_data_bus[792]), .B1(n7422), 
        .B2(i_data_bus[888]), .ZN(n7269) );
  ND2D1BWP30P140LVT U10677 ( .A1(n7270), .A2(n7269), .ZN(N1887) );
  AOI22D1BWP30P140LVT U10678 ( .A1(n7425), .A2(i_data_bus[842]), .B1(n7423), 
        .B2(i_data_bus[810]), .ZN(n7272) );
  AOI22D1BWP30P140LVT U10679 ( .A1(n7424), .A2(i_data_bus[778]), .B1(n7422), 
        .B2(i_data_bus[874]), .ZN(n7271) );
  ND2D1BWP30P140LVT U10680 ( .A1(n7272), .A2(n7271), .ZN(N1873) );
  AOI22D1BWP30P140LVT U10681 ( .A1(n7425), .A2(i_data_bus[839]), .B1(n7423), 
        .B2(i_data_bus[807]), .ZN(n7274) );
  AOI22D1BWP30P140LVT U10682 ( .A1(n7424), .A2(i_data_bus[775]), .B1(n7422), 
        .B2(i_data_bus[871]), .ZN(n7273) );
  ND2D1BWP30P140LVT U10683 ( .A1(n7274), .A2(n7273), .ZN(N1870) );
  AOI22D1BWP30P140LVT U10684 ( .A1(n7425), .A2(i_data_bus[836]), .B1(n7423), 
        .B2(i_data_bus[804]), .ZN(n7276) );
  AOI22D1BWP30P140LVT U10685 ( .A1(n7424), .A2(i_data_bus[772]), .B1(n7422), 
        .B2(i_data_bus[868]), .ZN(n7275) );
  ND2D1BWP30P140LVT U10686 ( .A1(n7276), .A2(n7275), .ZN(N1867) );
  AOI22D1BWP30P140LVT U10687 ( .A1(i_data_bus[830]), .A2(n7336), .B1(
        i_data_bus[862]), .B2(n7334), .ZN(n7278) );
  AOI22D1BWP30P140LVT U10688 ( .A1(i_data_bus[894]), .A2(n7333), .B1(
        i_data_bus[798]), .B2(n7335), .ZN(n7277) );
  ND2D1BWP30P140LVT U10689 ( .A1(n7278), .A2(n7277), .ZN(N11047) );
  AOI22D1BWP30P140LVT U10690 ( .A1(i_data_bus[858]), .A2(n7334), .B1(
        i_data_bus[826]), .B2(n7336), .ZN(n7280) );
  AOI22D1BWP30P140LVT U10691 ( .A1(i_data_bus[890]), .A2(n7333), .B1(
        i_data_bus[794]), .B2(n7335), .ZN(n7279) );
  ND2D1BWP30P140LVT U10692 ( .A1(n7280), .A2(n7279), .ZN(N11043) );
  AOI22D1BWP30P140LVT U10693 ( .A1(i_data_bus[879]), .A2(n7333), .B1(
        i_data_bus[847]), .B2(n7334), .ZN(n7282) );
  AOI22D1BWP30P140LVT U10694 ( .A1(i_data_bus[815]), .A2(n7336), .B1(
        i_data_bus[783]), .B2(n7335), .ZN(n7281) );
  ND2D1BWP30P140LVT U10695 ( .A1(n7282), .A2(n7281), .ZN(N11032) );
  AOI22D1BWP30P140LVT U10696 ( .A1(i_data_bus[894]), .A2(n7301), .B1(
        i_data_bus[862]), .B2(n7302), .ZN(n7284) );
  AOI22D1BWP30P140LVT U10697 ( .A1(i_data_bus[830]), .A2(n7304), .B1(
        i_data_bus[798]), .B2(n7303), .ZN(n7283) );
  ND2D1BWP30P140LVT U10698 ( .A1(n7284), .A2(n7283), .ZN(N4621) );
  AOI22D1BWP30P140LVT U10699 ( .A1(i_data_bus[854]), .A2(n7302), .B1(
        i_data_bus[886]), .B2(n7301), .ZN(n7286) );
  AOI22D1BWP30P140LVT U10700 ( .A1(i_data_bus[822]), .A2(n7304), .B1(
        i_data_bus[790]), .B2(n7303), .ZN(n7285) );
  ND2D1BWP30P140LVT U10701 ( .A1(n7286), .A2(n7285), .ZN(N4613) );
  AOI22D1BWP30P140LVT U10702 ( .A1(i_data_bus[817]), .A2(n7304), .B1(
        i_data_bus[849]), .B2(n7302), .ZN(n7288) );
  AOI22D1BWP30P140LVT U10703 ( .A1(i_data_bus[881]), .A2(n7301), .B1(
        i_data_bus[785]), .B2(n7303), .ZN(n7287) );
  ND2D1BWP30P140LVT U10704 ( .A1(n7288), .A2(n7287), .ZN(N4608) );
  AOI22D1BWP30P140LVT U10705 ( .A1(i_data_bus[816]), .A2(n7304), .B1(
        i_data_bus[848]), .B2(n7302), .ZN(n7290) );
  AOI22D1BWP30P140LVT U10706 ( .A1(i_data_bus[880]), .A2(n7301), .B1(
        i_data_bus[784]), .B2(n7303), .ZN(n7289) );
  ND2D1BWP30P140LVT U10707 ( .A1(n7290), .A2(n7289), .ZN(N4607) );
  AOI22D1BWP30P140LVT U10708 ( .A1(i_data_bus[846]), .A2(n7302), .B1(
        i_data_bus[878]), .B2(n7301), .ZN(n7292) );
  AOI22D1BWP30P140LVT U10709 ( .A1(i_data_bus[814]), .A2(n7304), .B1(
        i_data_bus[782]), .B2(n7303), .ZN(n7291) );
  ND2D1BWP30P140LVT U10710 ( .A1(n7292), .A2(n7291), .ZN(N4605) );
  AOI22D1BWP30P140LVT U10711 ( .A1(i_data_bus[812]), .A2(n7304), .B1(
        i_data_bus[876]), .B2(n7301), .ZN(n7294) );
  AOI22D1BWP30P140LVT U10712 ( .A1(i_data_bus[844]), .A2(n7302), .B1(
        i_data_bus[780]), .B2(n7303), .ZN(n7293) );
  ND2D1BWP30P140LVT U10713 ( .A1(n7294), .A2(n7293), .ZN(N4603) );
  AOI22D1BWP30P140LVT U10714 ( .A1(i_data_bus[841]), .A2(n7302), .B1(
        i_data_bus[873]), .B2(n7301), .ZN(n7296) );
  AOI22D1BWP30P140LVT U10715 ( .A1(i_data_bus[809]), .A2(n7304), .B1(
        i_data_bus[777]), .B2(n7303), .ZN(n7295) );
  ND2D1BWP30P140LVT U10716 ( .A1(n7296), .A2(n7295), .ZN(N4600) );
  AOI22D1BWP30P140LVT U10717 ( .A1(i_data_bus[805]), .A2(n7304), .B1(
        i_data_bus[837]), .B2(n7302), .ZN(n7298) );
  AOI22D1BWP30P140LVT U10718 ( .A1(i_data_bus[869]), .A2(n7301), .B1(
        i_data_bus[773]), .B2(n7303), .ZN(n7297) );
  ND2D1BWP30P140LVT U10719 ( .A1(n7298), .A2(n7297), .ZN(N4596) );
  AOI22D1BWP30P140LVT U10720 ( .A1(i_data_bus[801]), .A2(n7336), .B1(
        i_data_bus[865]), .B2(n7333), .ZN(n7300) );
  AOI22D1BWP30P140LVT U10721 ( .A1(i_data_bus[833]), .A2(n7334), .B1(
        i_data_bus[769]), .B2(n7335), .ZN(n7299) );
  ND2D1BWP30P140LVT U10722 ( .A1(n7300), .A2(n7299), .ZN(N11018) );
  AOI22D1BWP30P140LVT U10723 ( .A1(i_data_bus[832]), .A2(n7302), .B1(
        i_data_bus[864]), .B2(n7301), .ZN(n7306) );
  AOI22D1BWP30P140LVT U10724 ( .A1(i_data_bus[800]), .A2(n7304), .B1(
        i_data_bus[768]), .B2(n7303), .ZN(n7305) );
  ND2D1BWP30P140LVT U10725 ( .A1(n7306), .A2(n7305), .ZN(N4591) );
  AOI22D1BWP30P140LVT U10726 ( .A1(i_data_bus[830]), .A2(n7326), .B1(
        i_data_bus[862]), .B2(n7324), .ZN(n7308) );
  AOI22D1BWP30P140LVT U10727 ( .A1(i_data_bus[894]), .A2(n7323), .B1(
        i_data_bus[798]), .B2(n7325), .ZN(n7307) );
  ND2D1BWP30P140LVT U10728 ( .A1(n7308), .A2(n7307), .ZN(N8323) );
  AOI22D1BWP30P140LVT U10729 ( .A1(i_data_bus[887]), .A2(n7323), .B1(
        i_data_bus[855]), .B2(n7324), .ZN(n7310) );
  AOI22D1BWP30P140LVT U10730 ( .A1(i_data_bus[823]), .A2(n7326), .B1(
        i_data_bus[791]), .B2(n7325), .ZN(n7309) );
  ND2D1BWP30P140LVT U10731 ( .A1(n7310), .A2(n7309), .ZN(N8316) );
  AOI22D1BWP30P140LVT U10732 ( .A1(i_data_bus[852]), .A2(n7324), .B1(
        i_data_bus[884]), .B2(n7323), .ZN(n7312) );
  AOI22D1BWP30P140LVT U10733 ( .A1(i_data_bus[820]), .A2(n7326), .B1(
        i_data_bus[788]), .B2(n7325), .ZN(n7311) );
  ND2D1BWP30P140LVT U10734 ( .A1(n7312), .A2(n7311), .ZN(N8313) );
  AOI22D1BWP30P140LVT U10735 ( .A1(i_data_bus[883]), .A2(n7323), .B1(
        i_data_bus[851]), .B2(n7324), .ZN(n7314) );
  AOI22D1BWP30P140LVT U10736 ( .A1(i_data_bus[819]), .A2(n7326), .B1(
        i_data_bus[787]), .B2(n7325), .ZN(n7313) );
  ND2D1BWP30P140LVT U10737 ( .A1(n7314), .A2(n7313), .ZN(N8312) );
  AOI22D1BWP30P140LVT U10738 ( .A1(i_data_bus[815]), .A2(n7326), .B1(
        i_data_bus[847]), .B2(n7324), .ZN(n7316) );
  AOI22D1BWP30P140LVT U10739 ( .A1(i_data_bus[879]), .A2(n7323), .B1(
        i_data_bus[783]), .B2(n7325), .ZN(n7315) );
  ND2D1BWP30P140LVT U10740 ( .A1(n7316), .A2(n7315), .ZN(N8308) );
  AOI22D1BWP30P140LVT U10741 ( .A1(i_data_bus[812]), .A2(n7326), .B1(
        i_data_bus[876]), .B2(n7323), .ZN(n7318) );
  AOI22D1BWP30P140LVT U10742 ( .A1(i_data_bus[844]), .A2(n7324), .B1(
        i_data_bus[780]), .B2(n7325), .ZN(n7317) );
  ND2D1BWP30P140LVT U10743 ( .A1(n7318), .A2(n7317), .ZN(N8305) );
  AOI22D1BWP30P140LVT U10744 ( .A1(i_data_bus[869]), .A2(n7323), .B1(
        i_data_bus[837]), .B2(n7324), .ZN(n7320) );
  AOI22D1BWP30P140LVT U10745 ( .A1(i_data_bus[805]), .A2(n7326), .B1(
        i_data_bus[773]), .B2(n7325), .ZN(n7319) );
  ND2D1BWP30P140LVT U10746 ( .A1(n7320), .A2(n7319), .ZN(N8298) );
  AOI22D1BWP30P140LVT U10747 ( .A1(i_data_bus[801]), .A2(n7326), .B1(
        i_data_bus[865]), .B2(n7323), .ZN(n7322) );
  AOI22D1BWP30P140LVT U10748 ( .A1(i_data_bus[833]), .A2(n7324), .B1(
        i_data_bus[769]), .B2(n7325), .ZN(n7321) );
  ND2D1BWP30P140LVT U10749 ( .A1(n7322), .A2(n7321), .ZN(N8294) );
  AOI22D1BWP30P140LVT U10750 ( .A1(i_data_bus[832]), .A2(n7324), .B1(
        i_data_bus[864]), .B2(n7323), .ZN(n7328) );
  AOI22D1BWP30P140LVT U10751 ( .A1(i_data_bus[800]), .A2(n7326), .B1(
        i_data_bus[768]), .B2(n7325), .ZN(n7327) );
  ND2D1BWP30P140LVT U10752 ( .A1(n7328), .A2(n7327), .ZN(N8293) );
  AOI22D1BWP30P140LVT U10753 ( .A1(i_data_bus[814]), .A2(n7336), .B1(
        i_data_bus[878]), .B2(n7333), .ZN(n7330) );
  AOI22D1BWP30P140LVT U10754 ( .A1(i_data_bus[846]), .A2(n7334), .B1(
        i_data_bus[782]), .B2(n7335), .ZN(n7329) );
  ND2D1BWP30P140LVT U10755 ( .A1(n7330), .A2(n7329), .ZN(N11031) );
  AOI22D1BWP30P140LVT U10756 ( .A1(i_data_bus[880]), .A2(n7333), .B1(
        i_data_bus[848]), .B2(n7334), .ZN(n7332) );
  AOI22D1BWP30P140LVT U10757 ( .A1(i_data_bus[816]), .A2(n7336), .B1(
        i_data_bus[784]), .B2(n7335), .ZN(n7331) );
  ND2D1BWP30P140LVT U10758 ( .A1(n7332), .A2(n7331), .ZN(N11033) );
  AOI22D1BWP30P140LVT U10759 ( .A1(i_data_bus[854]), .A2(n7334), .B1(
        i_data_bus[886]), .B2(n7333), .ZN(n7338) );
  AOI22D1BWP30P140LVT U10760 ( .A1(i_data_bus[822]), .A2(n7336), .B1(
        i_data_bus[790]), .B2(n7335), .ZN(n7337) );
  ND2D1BWP30P140LVT U10761 ( .A1(n7338), .A2(n7337), .ZN(N11039) );
  AOI22D1BWP30P140LVT U10762 ( .A1(i_data_bus[892]), .A2(n7354), .B1(
        i_data_bus[828]), .B2(n7352), .ZN(n7340) );
  AOI22D1BWP30P140LVT U10763 ( .A1(i_data_bus[860]), .A2(n7351), .B1(
        i_data_bus[796]), .B2(n7353), .ZN(n7339) );
  ND2D1BWP30P140LVT U10764 ( .A1(n7340), .A2(n7339), .ZN(N2873) );
  AOI22D1BWP30P140LVT U10765 ( .A1(i_data_bus[890]), .A2(n7354), .B1(
        i_data_bus[826]), .B2(n7352), .ZN(n7342) );
  AOI22D1BWP30P140LVT U10766 ( .A1(i_data_bus[858]), .A2(n7351), .B1(
        i_data_bus[794]), .B2(n7353), .ZN(n7341) );
  ND2D1BWP30P140LVT U10767 ( .A1(n7342), .A2(n7341), .ZN(N2871) );
  AOI22D1BWP30P140LVT U10768 ( .A1(i_data_bus[880]), .A2(n7354), .B1(
        i_data_bus[848]), .B2(n7351), .ZN(n7344) );
  AOI22D1BWP30P140LVT U10769 ( .A1(i_data_bus[816]), .A2(n7352), .B1(
        i_data_bus[784]), .B2(n7353), .ZN(n7343) );
  ND2D1BWP30P140LVT U10770 ( .A1(n7344), .A2(n7343), .ZN(N2861) );
  AOI22D1BWP30P140LVT U10771 ( .A1(i_data_bus[815]), .A2(n7352), .B1(
        i_data_bus[847]), .B2(n7351), .ZN(n7346) );
  AOI22D1BWP30P140LVT U10772 ( .A1(i_data_bus[879]), .A2(n7354), .B1(
        i_data_bus[783]), .B2(n7353), .ZN(n7345) );
  ND2D1BWP30P140LVT U10773 ( .A1(n7346), .A2(n7345), .ZN(N2860) );
  AOI22D1BWP30P140LVT U10774 ( .A1(i_data_bus[806]), .A2(n7352), .B1(
        i_data_bus[838]), .B2(n7351), .ZN(n7348) );
  AOI22D1BWP30P140LVT U10775 ( .A1(i_data_bus[870]), .A2(n7354), .B1(
        i_data_bus[774]), .B2(n7353), .ZN(n7347) );
  ND2D1BWP30P140LVT U10776 ( .A1(n7348), .A2(n7347), .ZN(N2851) );
  AOI22D1BWP30P140LVT U10777 ( .A1(i_data_bus[869]), .A2(n7354), .B1(
        i_data_bus[837]), .B2(n7351), .ZN(n7350) );
  AOI22D1BWP30P140LVT U10778 ( .A1(i_data_bus[805]), .A2(n7352), .B1(
        i_data_bus[773]), .B2(n7353), .ZN(n7349) );
  ND2D1BWP30P140LVT U10779 ( .A1(n7350), .A2(n7349), .ZN(N2850) );
  AOI22D1BWP30P140LVT U10780 ( .A1(i_data_bus[801]), .A2(n7352), .B1(
        i_data_bus[833]), .B2(n7351), .ZN(n7356) );
  AOI22D1BWP30P140LVT U10781 ( .A1(i_data_bus[865]), .A2(n7354), .B1(
        i_data_bus[769]), .B2(n7353), .ZN(n7355) );
  ND2D1BWP30P140LVT U10782 ( .A1(n7356), .A2(n7355), .ZN(N2846) );
  AOI22D1BWP30P140LVT U10783 ( .A1(i_data_bus[890]), .A2(n7363), .B1(
        i_data_bus[826]), .B2(n7366), .ZN(n7358) );
  AOI22D1BWP30P140LVT U10784 ( .A1(i_data_bus[858]), .A2(n7364), .B1(
        i_data_bus[794]), .B2(n7365), .ZN(n7357) );
  ND2D1BWP30P140LVT U10785 ( .A1(n7358), .A2(n7357), .ZN(N10065) );
  AOI22D1BWP30P140LVT U10786 ( .A1(i_data_bus[883]), .A2(n7363), .B1(
        i_data_bus[851]), .B2(n7364), .ZN(n7360) );
  AOI22D1BWP30P140LVT U10787 ( .A1(i_data_bus[819]), .A2(n7366), .B1(
        i_data_bus[787]), .B2(n7365), .ZN(n7359) );
  ND2D1BWP30P140LVT U10788 ( .A1(n7360), .A2(n7359), .ZN(N10058) );
  AOI22D1BWP30P140LVT U10789 ( .A1(i_data_bus[881]), .A2(n7363), .B1(
        i_data_bus[849]), .B2(n7364), .ZN(n7362) );
  AOI22D1BWP30P140LVT U10790 ( .A1(i_data_bus[817]), .A2(n7366), .B1(
        i_data_bus[785]), .B2(n7365), .ZN(n7361) );
  ND2D1BWP30P140LVT U10791 ( .A1(n7362), .A2(n7361), .ZN(N10056) );
  AOI22D1BWP30P140LVT U10792 ( .A1(i_data_bus[841]), .A2(n7364), .B1(
        i_data_bus[873]), .B2(n7363), .ZN(n7368) );
  AOI22D1BWP30P140LVT U10793 ( .A1(i_data_bus[809]), .A2(n7366), .B1(
        i_data_bus[777]), .B2(n7365), .ZN(n7367) );
  ND2D1BWP30P140LVT U10794 ( .A1(n7368), .A2(n7367), .ZN(N10048) );
  NR4D0BWP30P140LVT U10795 ( .A1(inner_first_stage_valid_reg[49]), .A2(
        inner_first_stage_valid_reg[53]), .A3(inner_first_stage_valid_reg[51]), 
        .A4(inner_first_stage_valid_reg[50]), .ZN(n7373) );
  INR3D2BWP30P140LVT U10796 ( .A1(inner_first_stage_valid_reg[54]), .B1(
        inner_first_stage_valid_reg[55]), .B2(n7370), .ZN(n12160) );
  INR3D2BWP30P140LVT U10797 ( .A1(inner_first_stage_valid_reg[55]), .B1(
        inner_first_stage_valid_reg[54]), .B2(n7370), .ZN(n12159) );
  NR2D1BWP30P140LVT U10798 ( .A1(inner_first_stage_valid_reg[51]), .A2(
        inner_first_stage_valid_reg[50]), .ZN(n7371) );
  NR3D0P7BWP30P140LVT U10799 ( .A1(inner_first_stage_valid_reg[48]), .A2(
        inner_first_stage_valid_reg[54]), .A3(inner_first_stage_valid_reg[55]), 
        .ZN(n7374) );
  INR3D0BWP30P140LVT U10800 ( .A1(n7374), .B1(inner_first_stage_valid_reg[52]), 
        .B2(n11173), .ZN(n7377) );
  INR3D2BWP30P140LVT U10801 ( .A1(inner_first_stage_valid_reg[49]), .B1(
        inner_first_stage_valid_reg[53]), .B2(n7372), .ZN(n12162) );
  INR3D2BWP30P140LVT U10802 ( .A1(inner_first_stage_valid_reg[53]), .B1(
        inner_first_stage_valid_reg[49]), .B2(n7372), .ZN(n12161) );
  NR4D0BWP30P140LVT U10803 ( .A1(n12160), .A2(n12159), .A3(n12162), .A4(n12161), .ZN(n7381) );
  NR2D1BWP30P140LVT U10804 ( .A1(inner_first_stage_valid_reg[49]), .A2(
        inner_first_stage_valid_reg[53]), .ZN(n7378) );
  INR3D2BWP30P140LVT U10805 ( .A1(inner_first_stage_valid_reg[51]), .B1(
        inner_first_stage_valid_reg[50]), .B2(n7379), .ZN(n12158) );
  INR3D2BWP30P140LVT U10806 ( .A1(inner_first_stage_valid_reg[50]), .B1(
        inner_first_stage_valid_reg[51]), .B2(n7379), .ZN(n12157) );
  NR4D0BWP30P140LVT U10807 ( .A1(n12156), .A2(n7376), .A3(n12158), .A4(n12157), 
        .ZN(n7380) );
  AOI22D1BWP30P140LVT U10808 ( .A1(n7425), .A2(i_data_bus[862]), .B1(n7424), 
        .B2(i_data_bus[798]), .ZN(n7383) );
  AOI22D1BWP30P140LVT U10809 ( .A1(n7423), .A2(i_data_bus[830]), .B1(n7422), 
        .B2(i_data_bus[894]), .ZN(n7382) );
  ND2D1BWP30P140LVT U10810 ( .A1(n7383), .A2(n7382), .ZN(N1893) );
  AOI22D1BWP30P140LVT U10811 ( .A1(n7425), .A2(i_data_bus[861]), .B1(n7424), 
        .B2(i_data_bus[797]), .ZN(n7385) );
  AOI22D1BWP30P140LVT U10812 ( .A1(n7423), .A2(i_data_bus[829]), .B1(n7422), 
        .B2(i_data_bus[893]), .ZN(n7384) );
  ND2D1BWP30P140LVT U10813 ( .A1(n7385), .A2(n7384), .ZN(N1892) );
  AOI22D1BWP30P140LVT U10814 ( .A1(n7423), .A2(i_data_bus[828]), .B1(n7424), 
        .B2(i_data_bus[796]), .ZN(n7387) );
  AOI22D1BWP30P140LVT U10815 ( .A1(n7425), .A2(i_data_bus[860]), .B1(n7422), 
        .B2(i_data_bus[892]), .ZN(n7386) );
  ND2D1BWP30P140LVT U10816 ( .A1(n7387), .A2(n7386), .ZN(N1891) );
  AOI22D1BWP30P140LVT U10817 ( .A1(n7423), .A2(i_data_bus[826]), .B1(n7424), 
        .B2(i_data_bus[794]), .ZN(n7389) );
  AOI22D1BWP30P140LVT U10818 ( .A1(n7425), .A2(i_data_bus[858]), .B1(n7422), 
        .B2(i_data_bus[890]), .ZN(n7388) );
  ND2D1BWP30P140LVT U10819 ( .A1(n7389), .A2(n7388), .ZN(N1889) );
  AOI22D1BWP30P140LVT U10820 ( .A1(n7425), .A2(i_data_bus[855]), .B1(n7424), 
        .B2(i_data_bus[791]), .ZN(n7391) );
  AOI22D1BWP30P140LVT U10821 ( .A1(n7423), .A2(i_data_bus[823]), .B1(n7422), 
        .B2(i_data_bus[887]), .ZN(n7390) );
  ND2D1BWP30P140LVT U10822 ( .A1(n7391), .A2(n7390), .ZN(N1886) );
  AOI22D1BWP30P140LVT U10823 ( .A1(n7423), .A2(i_data_bus[822]), .B1(n7424), 
        .B2(i_data_bus[790]), .ZN(n7393) );
  AOI22D1BWP30P140LVT U10824 ( .A1(n7425), .A2(i_data_bus[854]), .B1(n7422), 
        .B2(i_data_bus[886]), .ZN(n7392) );
  ND2D1BWP30P140LVT U10825 ( .A1(n7393), .A2(n7392), .ZN(N1885) );
  AOI22D1BWP30P140LVT U10826 ( .A1(n7425), .A2(i_data_bus[851]), .B1(n7424), 
        .B2(i_data_bus[787]), .ZN(n7395) );
  AOI22D1BWP30P140LVT U10827 ( .A1(n7423), .A2(i_data_bus[819]), .B1(n7422), 
        .B2(i_data_bus[883]), .ZN(n7394) );
  ND2D1BWP30P140LVT U10828 ( .A1(n7395), .A2(n7394), .ZN(N1882) );
  AOI22D1BWP30P140LVT U10829 ( .A1(n7425), .A2(i_data_bus[849]), .B1(n7424), 
        .B2(i_data_bus[785]), .ZN(n7397) );
  AOI22D1BWP30P140LVT U10830 ( .A1(n7423), .A2(i_data_bus[817]), .B1(n7422), 
        .B2(i_data_bus[881]), .ZN(n7396) );
  ND2D1BWP30P140LVT U10831 ( .A1(n7397), .A2(n7396), .ZN(N1880) );
  AOI22D1BWP30P140LVT U10832 ( .A1(n7425), .A2(i_data_bus[848]), .B1(n7424), 
        .B2(i_data_bus[784]), .ZN(n7399) );
  AOI22D1BWP30P140LVT U10833 ( .A1(n7423), .A2(i_data_bus[816]), .B1(n7422), 
        .B2(i_data_bus[880]), .ZN(n7398) );
  ND2D1BWP30P140LVT U10834 ( .A1(n7399), .A2(n7398), .ZN(N1879) );
  AOI22D1BWP30P140LVT U10835 ( .A1(n7425), .A2(i_data_bus[847]), .B1(n7424), 
        .B2(i_data_bus[783]), .ZN(n7401) );
  AOI22D1BWP30P140LVT U10836 ( .A1(n7423), .A2(i_data_bus[815]), .B1(n7422), 
        .B2(i_data_bus[879]), .ZN(n7400) );
  ND2D1BWP30P140LVT U10837 ( .A1(n7401), .A2(n7400), .ZN(N1878) );
  AOI22D1BWP30P140LVT U10838 ( .A1(n7425), .A2(i_data_bus[838]), .B1(n7424), 
        .B2(i_data_bus[774]), .ZN(n7403) );
  AOI22D1BWP30P140LVT U10839 ( .A1(n7423), .A2(i_data_bus[806]), .B1(n7422), 
        .B2(i_data_bus[870]), .ZN(n7402) );
  ND2D1BWP30P140LVT U10840 ( .A1(n7403), .A2(n7402), .ZN(N1869) );
  AOI22D1BWP30P140LVT U10841 ( .A1(n7425), .A2(i_data_bus[837]), .B1(n7424), 
        .B2(i_data_bus[773]), .ZN(n7405) );
  AOI22D1BWP30P140LVT U10842 ( .A1(n7423), .A2(i_data_bus[805]), .B1(n7422), 
        .B2(i_data_bus[869]), .ZN(n7404) );
  ND2D1BWP30P140LVT U10843 ( .A1(n7405), .A2(n7404), .ZN(N1868) );
  AOI22D1BWP30P140LVT U10844 ( .A1(n7425), .A2(i_data_bus[833]), .B1(n7424), 
        .B2(i_data_bus[769]), .ZN(n7407) );
  AOI22D1BWP30P140LVT U10845 ( .A1(n7423), .A2(i_data_bus[801]), .B1(n7422), 
        .B2(i_data_bus[865]), .ZN(n7406) );
  ND2D1BWP30P140LVT U10846 ( .A1(n7407), .A2(n7406), .ZN(N1864) );
  AOI22D1BWP30P140LVT U10847 ( .A1(n7425), .A2(i_data_bus[859]), .B1(n7422), 
        .B2(i_data_bus[891]), .ZN(n7409) );
  AOI22D1BWP30P140LVT U10848 ( .A1(n7423), .A2(i_data_bus[827]), .B1(n7424), 
        .B2(i_data_bus[795]), .ZN(n7408) );
  ND2D1BWP30P140LVT U10849 ( .A1(n7409), .A2(n7408), .ZN(N1890) );
  AOI22D1BWP30P140LVT U10850 ( .A1(n7425), .A2(i_data_bus[857]), .B1(n7422), 
        .B2(i_data_bus[889]), .ZN(n7411) );
  AOI22D1BWP30P140LVT U10851 ( .A1(n7423), .A2(i_data_bus[825]), .B1(n7424), 
        .B2(i_data_bus[793]), .ZN(n7410) );
  ND2D1BWP30P140LVT U10852 ( .A1(n7411), .A2(n7410), .ZN(N1888) );
  AOI22D1BWP30P140LVT U10853 ( .A1(n7423), .A2(i_data_bus[821]), .B1(n7422), 
        .B2(i_data_bus[885]), .ZN(n7413) );
  AOI22D1BWP30P140LVT U10854 ( .A1(n7425), .A2(i_data_bus[853]), .B1(n7424), 
        .B2(i_data_bus[789]), .ZN(n7412) );
  ND2D1BWP30P140LVT U10855 ( .A1(n7413), .A2(n7412), .ZN(N1884) );
  AOI22D1BWP30P140LVT U10856 ( .A1(n7425), .A2(i_data_bus[850]), .B1(n7422), 
        .B2(i_data_bus[882]), .ZN(n7415) );
  AOI22D1BWP30P140LVT U10857 ( .A1(n7423), .A2(i_data_bus[818]), .B1(n7424), 
        .B2(i_data_bus[786]), .ZN(n7414) );
  ND2D1BWP30P140LVT U10858 ( .A1(n7415), .A2(n7414), .ZN(N1881) );
  AOI22D1BWP30P140LVT U10859 ( .A1(n7423), .A2(i_data_bus[811]), .B1(n7422), 
        .B2(i_data_bus[875]), .ZN(n7417) );
  AOI22D1BWP30P140LVT U10860 ( .A1(n7425), .A2(i_data_bus[843]), .B1(n7424), 
        .B2(i_data_bus[779]), .ZN(n7416) );
  ND2D1BWP30P140LVT U10861 ( .A1(n7417), .A2(n7416), .ZN(N1874) );
  AOI22D1BWP30P140LVT U10862 ( .A1(n7423), .A2(i_data_bus[808]), .B1(n7422), 
        .B2(i_data_bus[872]), .ZN(n7419) );
  AOI22D1BWP30P140LVT U10863 ( .A1(n7425), .A2(i_data_bus[840]), .B1(n7424), 
        .B2(i_data_bus[776]), .ZN(n7418) );
  ND2D1BWP30P140LVT U10864 ( .A1(n7419), .A2(n7418), .ZN(N1871) );
  AOI22D1BWP30P140LVT U10865 ( .A1(n7425), .A2(i_data_bus[835]), .B1(n7422), 
        .B2(i_data_bus[867]), .ZN(n7421) );
  AOI22D1BWP30P140LVT U10866 ( .A1(n7423), .A2(i_data_bus[803]), .B1(n7424), 
        .B2(i_data_bus[771]), .ZN(n7420) );
  ND2D1BWP30P140LVT U10867 ( .A1(n7421), .A2(n7420), .ZN(N1866) );
  AOI22D1BWP30P140LVT U10868 ( .A1(n7423), .A2(i_data_bus[802]), .B1(n7422), 
        .B2(i_data_bus[866]), .ZN(n7427) );
  AOI22D1BWP30P140LVT U10869 ( .A1(n7425), .A2(i_data_bus[834]), .B1(n7424), 
        .B2(i_data_bus[770]), .ZN(n7426) );
  ND2D1BWP30P140LVT U10870 ( .A1(n7427), .A2(n7426), .ZN(N1865) );
  AOI22D1BWP30P140LVT U10871 ( .A1(i_data_bus[444]), .A2(n8041), .B1(
        i_data_bus[412]), .B2(n6212), .ZN(n7433) );
  AOI22D1BWP30P140LVT U10872 ( .A1(i_data_bus[508]), .A2(n7443), .B1(
        i_data_bus[476]), .B2(n7434), .ZN(n7432) );
  ND2D1BWP30P140LVT U10873 ( .A1(n7433), .A2(n7432), .ZN(N1231) );
  AOI22D1BWP30P140LVT U10874 ( .A1(i_data_bus[440]), .A2(n8041), .B1(
        i_data_bus[472]), .B2(n7434), .ZN(n7436) );
  AOI22D1BWP30P140LVT U10875 ( .A1(i_data_bus[504]), .A2(n7443), .B1(
        i_data_bus[408]), .B2(n6212), .ZN(n7435) );
  ND2D1BWP30P140LVT U10876 ( .A1(n7436), .A2(n7435), .ZN(N1227) );
  AOI22D1BWP30P140LVT U10877 ( .A1(i_data_bus[435]), .A2(n8041), .B1(
        i_data_bus[499]), .B2(n7443), .ZN(n7438) );
  AOI22D1BWP30P140LVT U10878 ( .A1(i_data_bus[403]), .A2(n6212), .B1(
        i_data_bus[467]), .B2(n7434), .ZN(n7437) );
  ND2D1BWP30P140LVT U10879 ( .A1(n7438), .A2(n7437), .ZN(N1222) );
  AOI22D1BWP30P140LVT U10880 ( .A1(i_data_bus[434]), .A2(n8041), .B1(
        i_data_bus[466]), .B2(n7434), .ZN(n7440) );
  AOI22D1BWP30P140LVT U10881 ( .A1(i_data_bus[498]), .A2(n7443), .B1(
        i_data_bus[402]), .B2(n6212), .ZN(n7439) );
  ND2D1BWP30P140LVT U10882 ( .A1(n7440), .A2(n7439), .ZN(N1221) );
  AOI22D1BWP30P140LVT U10883 ( .A1(i_data_bus[430]), .A2(n8041), .B1(
        i_data_bus[462]), .B2(n7434), .ZN(n7442) );
  AOI22D1BWP30P140LVT U10884 ( .A1(i_data_bus[398]), .A2(n6212), .B1(
        i_data_bus[494]), .B2(n7443), .ZN(n7441) );
  ND2D1BWP30P140LVT U10885 ( .A1(n7442), .A2(n7441), .ZN(N1217) );
  AOI22D1BWP30P140LVT U10886 ( .A1(i_data_bus[429]), .A2(n8041), .B1(
        i_data_bus[493]), .B2(n7443), .ZN(n7445) );
  AOI22D1BWP30P140LVT U10887 ( .A1(i_data_bus[397]), .A2(n6212), .B1(
        i_data_bus[461]), .B2(n7434), .ZN(n7444) );
  ND2D1BWP30P140LVT U10888 ( .A1(n7445), .A2(n7444), .ZN(N1216) );
  AOI22D1BWP30P140LVT U10889 ( .A1(i_data_bus[426]), .A2(n8041), .B1(
        i_data_bus[458]), .B2(n7434), .ZN(n7447) );
  AOI22D1BWP30P140LVT U10890 ( .A1(i_data_bus[490]), .A2(n7443), .B1(
        i_data_bus[394]), .B2(n6212), .ZN(n7446) );
  ND2D1BWP30P140LVT U10891 ( .A1(n7447), .A2(n7446), .ZN(N1213) );
  AOI22D1BWP30P140LVT U10892 ( .A1(i_data_bus[422]), .A2(n8041), .B1(
        i_data_bus[454]), .B2(n7434), .ZN(n7449) );
  AOI22D1BWP30P140LVT U10893 ( .A1(i_data_bus[390]), .A2(n6212), .B1(
        i_data_bus[486]), .B2(n7443), .ZN(n7448) );
  ND2D1BWP30P140LVT U10894 ( .A1(n7449), .A2(n7448), .ZN(N1209) );
  AOI22D1BWP30P140LVT U10895 ( .A1(i_data_bus[421]), .A2(n8041), .B1(
        i_data_bus[389]), .B2(n6212), .ZN(n7451) );
  AOI22D1BWP30P140LVT U10896 ( .A1(i_data_bus[485]), .A2(n7443), .B1(
        i_data_bus[453]), .B2(n7434), .ZN(n7450) );
  ND2D1BWP30P140LVT U10897 ( .A1(n7451), .A2(n7450), .ZN(N1208) );
  NR2D1BWP30P140LVT U10898 ( .A1(inner_first_stage_valid_reg[26]), .A2(
        inner_first_stage_valid_reg[27]), .ZN(n7452) );
  NR3D0P7BWP30P140LVT U10899 ( .A1(inner_first_stage_valid_reg[31]), .A2(
        inner_first_stage_valid_reg[30]), .A3(n11173), .ZN(n7459) );
  INR3D0BWP30P140LVT U10900 ( .A1(n7459), .B1(inner_first_stage_valid_reg[28]), 
        .B2(inner_first_stage_valid_reg[24]), .ZN(n7454) );
  INR3D2BWP30P140LVT U10901 ( .A1(inner_first_stage_valid_reg[25]), .B1(
        inner_first_stage_valid_reg[29]), .B2(n7453), .ZN(n11755) );
  INR3D2BWP30P140LVT U10902 ( .A1(inner_first_stage_valid_reg[29]), .B1(
        inner_first_stage_valid_reg[25]), .B2(n7453), .ZN(n11753) );
  NR2D1BWP30P140LVT U10903 ( .A1(inner_first_stage_valid_reg[25]), .A2(
        inner_first_stage_valid_reg[29]), .ZN(n7455) );
  INR3D2BWP30P140LVT U10904 ( .A1(inner_first_stage_valid_reg[26]), .B1(
        inner_first_stage_valid_reg[27]), .B2(n7456), .ZN(n11754) );
  INR3D2BWP30P140LVT U10905 ( .A1(inner_first_stage_valid_reg[27]), .B1(
        inner_first_stage_valid_reg[26]), .B2(n7456), .ZN(n11752) );
  NR4D0BWP30P140LVT U10906 ( .A1(n11755), .A2(n11753), .A3(n11754), .A4(n11752), .ZN(n7463) );
  NR4D0BWP30P140LVT U10907 ( .A1(inner_first_stage_valid_reg[25]), .A2(
        inner_first_stage_valid_reg[29]), .A3(inner_first_stage_valid_reg[26]), 
        .A4(inner_first_stage_valid_reg[27]), .ZN(n7460) );
  NR2D1BWP30P140LVT U10908 ( .A1(inner_first_stage_valid_reg[28]), .A2(
        inner_first_stage_valid_reg[24]), .ZN(n7457) );
  ND3D1BWP30P140LVT U10909 ( .A1(n12302), .A2(n7460), .A3(n7457), .ZN(n7458)
         );
  INR3D2BWP30P140LVT U10910 ( .A1(inner_first_stage_valid_reg[31]), .B1(
        inner_first_stage_valid_reg[30]), .B2(n7458), .ZN(n11749) );
  INR3D2BWP30P140LVT U10911 ( .A1(inner_first_stage_valid_reg[30]), .B1(
        inner_first_stage_valid_reg[31]), .B2(n7458), .ZN(n11748) );
  INR3D2BWP30P140LVT U10912 ( .A1(inner_first_stage_valid_reg[24]), .B1(
        inner_first_stage_valid_reg[28]), .B2(n7461), .ZN(n11751) );
  INR3D2BWP30P140LVT U10913 ( .A1(inner_first_stage_valid_reg[28]), .B1(
        inner_first_stage_valid_reg[24]), .B2(n7461), .ZN(n11750) );
  NR4D0BWP30P140LVT U10914 ( .A1(n11749), .A2(n11748), .A3(n11751), .A4(n11750), .ZN(n7462) );
  AOI22D1BWP30P140LVT U10915 ( .A1(i_data_bus[387]), .A2(n6212), .B1(
        i_data_bus[483]), .B2(n7443), .ZN(n7465) );
  AOI22D1BWP30P140LVT U10916 ( .A1(i_data_bus[419]), .A2(n8041), .B1(
        i_data_bus[451]), .B2(n7434), .ZN(n7464) );
  ND2D1BWP30P140LVT U10917 ( .A1(n7465), .A2(n7464), .ZN(N1206) );
  AOI22D1BWP30P140LVT U10918 ( .A1(i_data_bus[449]), .A2(n7434), .B1(
        i_data_bus[481]), .B2(n7443), .ZN(n7467) );
  AOI22D1BWP30P140LVT U10919 ( .A1(i_data_bus[417]), .A2(n8041), .B1(
        i_data_bus[385]), .B2(n6212), .ZN(n7466) );
  ND2D1BWP30P140LVT U10920 ( .A1(n7467), .A2(n7466), .ZN(N1204) );
  AOI22D1BWP30P140LVT U10921 ( .A1(i_data_bus[480]), .A2(n7443), .B1(
        i_data_bus[384]), .B2(n6212), .ZN(n7469) );
  AOI22D1BWP30P140LVT U10922 ( .A1(i_data_bus[416]), .A2(n8041), .B1(
        i_data_bus[448]), .B2(n7434), .ZN(n7468) );
  ND2D1BWP30P140LVT U10923 ( .A1(n7469), .A2(n7468), .ZN(N1203) );
  AOI22D1BWP30P140LVT U10924 ( .A1(i_data_bus[414]), .A2(n6212), .B1(
        i_data_bus[478]), .B2(n7434), .ZN(n7471) );
  AOI22D1BWP30P140LVT U10925 ( .A1(i_data_bus[446]), .A2(n8041), .B1(
        i_data_bus[510]), .B2(n7443), .ZN(n7470) );
  ND2D1BWP30P140LVT U10926 ( .A1(n7471), .A2(n7470), .ZN(N1233) );
  AOI22D1BWP30P140LVT U10927 ( .A1(i_data_bus[407]), .A2(n6212), .B1(
        i_data_bus[471]), .B2(n7434), .ZN(n7473) );
  AOI22D1BWP30P140LVT U10928 ( .A1(i_data_bus[439]), .A2(n8041), .B1(
        i_data_bus[503]), .B2(n7443), .ZN(n7472) );
  ND2D1BWP30P140LVT U10929 ( .A1(n7473), .A2(n7472), .ZN(N1226) );
  AOI22D1BWP30P140LVT U10930 ( .A1(i_data_bus[401]), .A2(n6212), .B1(
        i_data_bus[465]), .B2(n7434), .ZN(n7475) );
  AOI22D1BWP30P140LVT U10931 ( .A1(i_data_bus[433]), .A2(n8041), .B1(
        i_data_bus[497]), .B2(n7443), .ZN(n7474) );
  ND2D1BWP30P140LVT U10932 ( .A1(n7475), .A2(n7474), .ZN(N1220) );
  AOI22D1BWP30P140LVT U10933 ( .A1(i_data_bus[492]), .A2(n7443), .B1(
        i_data_bus[460]), .B2(n7434), .ZN(n7477) );
  AOI22D1BWP30P140LVT U10934 ( .A1(i_data_bus[428]), .A2(n8041), .B1(
        i_data_bus[396]), .B2(n6212), .ZN(n7476) );
  ND2D1BWP30P140LVT U10935 ( .A1(n7477), .A2(n7476), .ZN(N1215) );
  AOI22D1BWP30P140LVT U10936 ( .A1(i_data_bus[489]), .A2(n7443), .B1(
        i_data_bus[393]), .B2(n6212), .ZN(n7479) );
  AOI22D1BWP30P140LVT U10937 ( .A1(i_data_bus[425]), .A2(n8041), .B1(
        i_data_bus[457]), .B2(n7434), .ZN(n7478) );
  ND2D1BWP30P140LVT U10938 ( .A1(n7479), .A2(n7478), .ZN(N1212) );
  AOI22D1BWP30P140LVT U10939 ( .A1(i_data_bus[391]), .A2(n6212), .B1(
        i_data_bus[455]), .B2(n7434), .ZN(n7481) );
  AOI22D1BWP30P140LVT U10940 ( .A1(i_data_bus[423]), .A2(n8041), .B1(
        i_data_bus[487]), .B2(n7443), .ZN(n7480) );
  ND2D1BWP30P140LVT U10941 ( .A1(n7481), .A2(n7480), .ZN(N1210) );
  AOI22D1BWP30P140LVT U10942 ( .A1(i_data_bus[452]), .A2(n7434), .B1(
        i_data_bus[484]), .B2(n7443), .ZN(n7483) );
  AOI22D1BWP30P140LVT U10943 ( .A1(i_data_bus[420]), .A2(n8041), .B1(
        i_data_bus[388]), .B2(n6212), .ZN(n7482) );
  ND2D1BWP30P140LVT U10944 ( .A1(n7483), .A2(n7482), .ZN(N1207) );
  INR4D1BWP30P140LVT U10945 ( .A1(i_cmd[243]), .B1(i_cmd[227]), .B2(n7765), 
        .B3(n11053), .ZN(n8207) );
  NR3D0P7BWP30P140LVT U10946 ( .A1(i_cmd[235]), .A2(i_cmd[251]), .A3(
        i_cmd[243]), .ZN(n11052) );
  AOI22D1BWP30P140LVT U10947 ( .A1(i_data_bus[990]), .A2(n8207), .B1(
        i_data_bus[926]), .B2(n8206), .ZN(n7486) );
  NR4D1BWP30P140LVT U10948 ( .A1(i_cmd[235]), .A2(n7771), .A3(n11055), .A4(
        n7484), .ZN(n8205) );
  AOI22D1BWP30P140LVT U10949 ( .A1(i_data_bus[958]), .A2(n8208), .B1(
        i_data_bus[1022]), .B2(n8205), .ZN(n7485) );
  ND2D1BWP30P140LVT U10950 ( .A1(n7486), .A2(n7485), .ZN(N5687) );
  AOI22D1BWP30P140LVT U10951 ( .A1(i_data_bus[971]), .A2(n8207), .B1(
        i_data_bus[907]), .B2(n8206), .ZN(n7488) );
  AOI22D1BWP30P140LVT U10952 ( .A1(i_data_bus[939]), .A2(n8208), .B1(
        i_data_bus[1003]), .B2(n8205), .ZN(n7487) );
  ND2D1BWP30P140LVT U10953 ( .A1(n7488), .A2(n7487), .ZN(N5668) );
  AOI22D1BWP30P140LVT U10954 ( .A1(i_data_bus[968]), .A2(n8207), .B1(
        i_data_bus[936]), .B2(n8208), .ZN(n7490) );
  AOI22D1BWP30P140LVT U10955 ( .A1(i_data_bus[1000]), .A2(n8205), .B1(
        i_data_bus[904]), .B2(n8206), .ZN(n7489) );
  ND2D1BWP30P140LVT U10956 ( .A1(n7490), .A2(n7489), .ZN(N5665) );
  AOI22D1BWP30P140LVT U10957 ( .A1(i_data_bus[961]), .A2(n8207), .B1(
        i_data_bus[929]), .B2(n8208), .ZN(n7492) );
  AOI22D1BWP30P140LVT U10958 ( .A1(i_data_bus[993]), .A2(n8205), .B1(
        i_data_bus[897]), .B2(n8206), .ZN(n7491) );
  ND2D1BWP30P140LVT U10959 ( .A1(n7492), .A2(n7491), .ZN(N5658) );
  AOI22D1BWP30P140LVT U10960 ( .A1(i_data_bus[988]), .A2(n8207), .B1(
        i_data_bus[956]), .B2(n8208), .ZN(n7494) );
  AOI22D1BWP30P140LVT U10961 ( .A1(i_data_bus[1020]), .A2(n8205), .B1(
        i_data_bus[924]), .B2(n8206), .ZN(n7493) );
  ND2D1BWP30P140LVT U10962 ( .A1(n7494), .A2(n7493), .ZN(N5685) );
  AOI22D1BWP30P140LVT U10963 ( .A1(i_data_bus[978]), .A2(n8207), .B1(
        i_data_bus[946]), .B2(n8208), .ZN(n7496) );
  AOI22D1BWP30P140LVT U10964 ( .A1(i_data_bus[914]), .A2(n8206), .B1(
        i_data_bus[1010]), .B2(n8205), .ZN(n7495) );
  ND2D1BWP30P140LVT U10965 ( .A1(n7496), .A2(n7495), .ZN(N5675) );
  AOI22D1BWP30P140LVT U10966 ( .A1(i_data_bus[969]), .A2(n8207), .B1(
        i_data_bus[937]), .B2(n8208), .ZN(n7498) );
  AOI22D1BWP30P140LVT U10967 ( .A1(i_data_bus[905]), .A2(n8206), .B1(
        i_data_bus[1001]), .B2(n8205), .ZN(n7497) );
  ND2D1BWP30P140LVT U10968 ( .A1(n7498), .A2(n7497), .ZN(N5666) );
  AOI22D1BWP30P140LVT U10969 ( .A1(i_data_bus[981]), .A2(n8207), .B1(
        i_data_bus[949]), .B2(n8208), .ZN(n7500) );
  AOI22D1BWP30P140LVT U10970 ( .A1(i_data_bus[917]), .A2(n8206), .B1(
        i_data_bus[1013]), .B2(n8205), .ZN(n7499) );
  ND2D1BWP30P140LVT U10971 ( .A1(n7500), .A2(n7499), .ZN(N5678) );
  AOI22D1BWP30P140LVT U10972 ( .A1(i_data_bus[975]), .A2(n8207), .B1(
        i_data_bus[1007]), .B2(n8205), .ZN(n7502) );
  AOI22D1BWP30P140LVT U10973 ( .A1(i_data_bus[943]), .A2(n8208), .B1(
        i_data_bus[911]), .B2(n8206), .ZN(n7501) );
  ND2D1BWP30P140LVT U10974 ( .A1(n7502), .A2(n7501), .ZN(N5672) );
  AOI22D1BWP30P140LVT U10975 ( .A1(i_data_bus[966]), .A2(n8207), .B1(
        i_data_bus[998]), .B2(n8205), .ZN(n7504) );
  AOI22D1BWP30P140LVT U10976 ( .A1(i_data_bus[934]), .A2(n8208), .B1(
        i_data_bus[902]), .B2(n8206), .ZN(n7503) );
  ND2D1BWP30P140LVT U10977 ( .A1(n7504), .A2(n7503), .ZN(N5663) );
  AOI22D1BWP30P140LVT U10978 ( .A1(i_data_bus[973]), .A2(n8207), .B1(
        i_data_bus[1005]), .B2(n8205), .ZN(n7506) );
  AOI22D1BWP30P140LVT U10979 ( .A1(i_data_bus[909]), .A2(n8206), .B1(
        i_data_bus[941]), .B2(n8208), .ZN(n7505) );
  ND2D1BWP30P140LVT U10980 ( .A1(n7506), .A2(n7505), .ZN(N5670) );
  AOI22D1BWP30P140LVT U10981 ( .A1(i_data_bus[970]), .A2(n8207), .B1(
        i_data_bus[1002]), .B2(n8205), .ZN(n7508) );
  AOI22D1BWP30P140LVT U10982 ( .A1(i_data_bus[906]), .A2(n8206), .B1(
        i_data_bus[938]), .B2(n8208), .ZN(n7507) );
  ND2D1BWP30P140LVT U10983 ( .A1(n7508), .A2(n7507), .ZN(N5667) );
  AOI22D1BWP30P140LVT U10984 ( .A1(i_data_bus[965]), .A2(n8207), .B1(
        i_data_bus[997]), .B2(n8205), .ZN(n7510) );
  AOI22D1BWP30P140LVT U10985 ( .A1(i_data_bus[901]), .A2(n8206), .B1(
        i_data_bus[933]), .B2(n8208), .ZN(n7509) );
  ND2D1BWP30P140LVT U10986 ( .A1(n7510), .A2(n7509), .ZN(N5662) );
  AOI22D1BWP30P140LVT U10987 ( .A1(i_data_bus[979]), .A2(n8207), .B1(
        i_data_bus[1011]), .B2(n8205), .ZN(n7512) );
  AOI22D1BWP30P140LVT U10988 ( .A1(i_data_bus[915]), .A2(n8206), .B1(
        i_data_bus[947]), .B2(n8208), .ZN(n7511) );
  ND2D1BWP30P140LVT U10989 ( .A1(n7512), .A2(n7511), .ZN(N5676) );
  OR2D1BWP30P140LVT U10990 ( .A1(i_cmd[237]), .A2(i_cmd[253]), .Z(n10972) );
  INR4D1BWP30P140LVT U10991 ( .A1(i_cmd[245]), .B1(i_cmd[229]), .B2(n7765), 
        .B3(n10972), .ZN(n8232) );
  INR4D1BWP30P140LVT U10992 ( .A1(i_cmd[237]), .B1(i_cmd[253]), .B2(n7769), 
        .B3(n7513), .ZN(n8231) );
  AOI22D1BWP30P140LVT U10993 ( .A1(i_data_bus[987]), .A2(n8232), .B1(
        i_data_bus[955]), .B2(n8231), .ZN(n7515) );
  NR3D0P7BWP30P140LVT U10994 ( .A1(i_cmd[237]), .A2(i_cmd[253]), .A3(
        i_cmd[245]), .ZN(n10968) );
  INR4D1BWP30P140LVT U10995 ( .A1(i_cmd[253]), .B1(i_cmd[237]), .B2(n7771), 
        .B3(n7513), .ZN(n8230) );
  AOI22D1BWP30P140LVT U10996 ( .A1(i_data_bus[923]), .A2(n8233), .B1(
        i_data_bus[1019]), .B2(n8230), .ZN(n7514) );
  ND2D1BWP30P140LVT U10997 ( .A1(n7515), .A2(n7514), .ZN(N8408) );
  AOI22D1BWP30P140LVT U10998 ( .A1(i_data_bus[961]), .A2(n8232), .B1(
        i_data_bus[929]), .B2(n8231), .ZN(n7517) );
  AOI22D1BWP30P140LVT U10999 ( .A1(i_data_bus[993]), .A2(n8230), .B1(
        i_data_bus[897]), .B2(n8233), .ZN(n7516) );
  ND2D1BWP30P140LVT U11000 ( .A1(n7517), .A2(n7516), .ZN(N8382) );
  AOI22D1BWP30P140LVT U11001 ( .A1(i_data_bus[986]), .A2(n8232), .B1(
        i_data_bus[1018]), .B2(n8230), .ZN(n7519) );
  AOI22D1BWP30P140LVT U11002 ( .A1(i_data_bus[922]), .A2(n8233), .B1(
        i_data_bus[954]), .B2(n8231), .ZN(n7518) );
  ND2D1BWP30P140LVT U11003 ( .A1(n7519), .A2(n7518), .ZN(N8407) );
  AOI22D1BWP30P140LVT U11004 ( .A1(i_data_bus[969]), .A2(n8232), .B1(
        i_data_bus[1001]), .B2(n8230), .ZN(n7521) );
  AOI22D1BWP30P140LVT U11005 ( .A1(i_data_bus[905]), .A2(n8233), .B1(
        i_data_bus[937]), .B2(n8231), .ZN(n7520) );
  ND2D1BWP30P140LVT U11006 ( .A1(n7521), .A2(n7520), .ZN(N8390) );
  AOI22D1BWP30P140LVT U11007 ( .A1(i_data_bus[968]), .A2(n8232), .B1(
        i_data_bus[1000]), .B2(n8230), .ZN(n7523) );
  AOI22D1BWP30P140LVT U11008 ( .A1(i_data_bus[904]), .A2(n8233), .B1(
        i_data_bus[936]), .B2(n8231), .ZN(n7522) );
  ND2D1BWP30P140LVT U11009 ( .A1(n7523), .A2(n7522), .ZN(N8389) );
  AOI22D1BWP30P140LVT U11010 ( .A1(i_data_bus[971]), .A2(n8232), .B1(
        i_data_bus[1003]), .B2(n8230), .ZN(n7525) );
  AOI22D1BWP30P140LVT U11011 ( .A1(i_data_bus[939]), .A2(n8231), .B1(
        i_data_bus[907]), .B2(n8233), .ZN(n7524) );
  ND2D1BWP30P140LVT U11012 ( .A1(n7525), .A2(n7524), .ZN(N8392) );
  AOI22D1BWP30P140LVT U11013 ( .A1(i_data_bus[980]), .A2(n8232), .B1(
        i_data_bus[916]), .B2(n8233), .ZN(n7527) );
  AOI22D1BWP30P140LVT U11014 ( .A1(i_data_bus[1012]), .A2(n8230), .B1(
        i_data_bus[948]), .B2(n8231), .ZN(n7526) );
  ND2D1BWP30P140LVT U11015 ( .A1(n7527), .A2(n7526), .ZN(N8401) );
  AOI22D1BWP30P140LVT U11016 ( .A1(i_data_bus[981]), .A2(n8232), .B1(
        i_data_bus[917]), .B2(n8233), .ZN(n7529) );
  AOI22D1BWP30P140LVT U11017 ( .A1(i_data_bus[949]), .A2(n8231), .B1(
        i_data_bus[1013]), .B2(n8230), .ZN(n7528) );
  ND2D1BWP30P140LVT U11018 ( .A1(n7529), .A2(n7528), .ZN(N8402) );
  INR4D1BWP30P140LVT U11019 ( .A1(i_cmd[247]), .B1(i_cmd[231]), .B2(n7765), 
        .B3(n10914), .ZN(n8257) );
  AOI22D1BWP30P140LVT U11020 ( .A1(i_data_bus[979]), .A2(n8257), .B1(
        i_data_bus[947]), .B2(n8256), .ZN(n7534) );
  NR3D0P7BWP30P140LVT U11021 ( .A1(i_cmd[247]), .A2(i_cmd[255]), .A3(
        i_cmd[239]), .ZN(n10910) );
  NR4D1BWP30P140LVT U11022 ( .A1(i_cmd[239]), .A2(n7532), .A3(n7771), .A4(
        n7531), .ZN(n8255) );
  AOI22D1BWP30P140LVT U11023 ( .A1(i_data_bus[915]), .A2(n8258), .B1(
        i_data_bus[1011]), .B2(n8255), .ZN(n7533) );
  ND2D1BWP30P140LVT U11024 ( .A1(n7534), .A2(n7533), .ZN(N11124) );
  AOI22D1BWP30P140LVT U11025 ( .A1(i_data_bus[969]), .A2(n8257), .B1(
        i_data_bus[937]), .B2(n8256), .ZN(n7536) );
  AOI22D1BWP30P140LVT U11026 ( .A1(i_data_bus[905]), .A2(n8258), .B1(
        i_data_bus[1001]), .B2(n8255), .ZN(n7535) );
  ND2D1BWP30P140LVT U11027 ( .A1(n7536), .A2(n7535), .ZN(N11114) );
  AOI22D1BWP30P140LVT U11028 ( .A1(i_data_bus[988]), .A2(n8257), .B1(
        i_data_bus[956]), .B2(n8256), .ZN(n7538) );
  AOI22D1BWP30P140LVT U11029 ( .A1(i_data_bus[1020]), .A2(n8255), .B1(
        i_data_bus[924]), .B2(n8258), .ZN(n7537) );
  ND2D1BWP30P140LVT U11030 ( .A1(n7538), .A2(n7537), .ZN(N11133) );
  AOI22D1BWP30P140LVT U11031 ( .A1(i_data_bus[977]), .A2(n8257), .B1(
        i_data_bus[1009]), .B2(n8255), .ZN(n7540) );
  AOI22D1BWP30P140LVT U11032 ( .A1(i_data_bus[913]), .A2(n8258), .B1(
        i_data_bus[945]), .B2(n8256), .ZN(n7539) );
  ND2D1BWP30P140LVT U11033 ( .A1(n7540), .A2(n7539), .ZN(N11122) );
  AOI22D1BWP30P140LVT U11034 ( .A1(i_data_bus[968]), .A2(n8257), .B1(
        i_data_bus[1000]), .B2(n8255), .ZN(n7542) );
  AOI22D1BWP30P140LVT U11035 ( .A1(i_data_bus[904]), .A2(n8258), .B1(
        i_data_bus[936]), .B2(n8256), .ZN(n7541) );
  ND2D1BWP30P140LVT U11036 ( .A1(n7542), .A2(n7541), .ZN(N11113) );
  AOI22D1BWP30P140LVT U11037 ( .A1(i_data_bus[974]), .A2(n8257), .B1(
        i_data_bus[910]), .B2(n8258), .ZN(n7544) );
  AOI22D1BWP30P140LVT U11038 ( .A1(i_data_bus[1006]), .A2(n8255), .B1(
        i_data_bus[942]), .B2(n8256), .ZN(n7543) );
  ND2D1BWP30P140LVT U11039 ( .A1(n7544), .A2(n7543), .ZN(N11119) );
  AOI22D1BWP30P140LVT U11040 ( .A1(i_data_bus[980]), .A2(n8257), .B1(
        i_data_bus[916]), .B2(n8258), .ZN(n7546) );
  AOI22D1BWP30P140LVT U11041 ( .A1(i_data_bus[1012]), .A2(n8255), .B1(
        i_data_bus[948]), .B2(n8256), .ZN(n7545) );
  ND2D1BWP30P140LVT U11042 ( .A1(n7546), .A2(n7545), .ZN(N11125) );
  AOI22D1BWP30P140LVT U11043 ( .A1(i_data_bus[991]), .A2(n8257), .B1(
        i_data_bus[927]), .B2(n8258), .ZN(n7548) );
  AOI22D1BWP30P140LVT U11044 ( .A1(i_data_bus[959]), .A2(n8256), .B1(
        i_data_bus[1023]), .B2(n8255), .ZN(n7547) );
  ND2D1BWP30P140LVT U11045 ( .A1(n7548), .A2(n7547), .ZN(N11136) );
  AOI22D1BWP30P140LVT U11046 ( .A1(i_data_bus[971]), .A2(n8257), .B1(
        i_data_bus[907]), .B2(n8258), .ZN(n7550) );
  AOI22D1BWP30P140LVT U11047 ( .A1(i_data_bus[939]), .A2(n8256), .B1(
        i_data_bus[1003]), .B2(n8255), .ZN(n7549) );
  ND2D1BWP30P140LVT U11048 ( .A1(n7550), .A2(n7549), .ZN(N11116) );
  INR4D1BWP30P140LVT U11049 ( .A1(i_cmd[242]), .B1(i_cmd[226]), .B2(n7765), 
        .B3(n7551), .ZN(n8353) );
  NR4D1BWP30P140LVT U11050 ( .A1(i_cmd[234]), .A2(n7771), .A3(n7552), .A4(
        n7554), .ZN(n8352) );
  AOI22D1BWP30P140LVT U11051 ( .A1(i_data_bus[983]), .A2(n8353), .B1(
        i_data_bus[1015]), .B2(n8352), .ZN(n7557) );
  AOI22D1BWP30P140LVT U11052 ( .A1(i_data_bus[919]), .A2(n8354), .B1(
        i_data_bus[951]), .B2(n8351), .ZN(n7556) );
  ND2D1BWP30P140LVT U11053 ( .A1(n7557), .A2(n7556), .ZN(N4830) );
  AOI22D1BWP30P140LVT U11054 ( .A1(i_data_bus[960]), .A2(n8353), .B1(
        i_data_bus[992]), .B2(n8352), .ZN(n7559) );
  AOI22D1BWP30P140LVT U11055 ( .A1(i_data_bus[896]), .A2(n8354), .B1(
        i_data_bus[928]), .B2(n8351), .ZN(n7558) );
  ND2D1BWP30P140LVT U11056 ( .A1(n7559), .A2(n7558), .ZN(N4807) );
  OR2D1BWP30P140LVT U11057 ( .A1(i_cmd[254]), .A2(i_cmd[238]), .Z(n10943) );
  INR4D1BWP30P140LVT U11058 ( .A1(i_cmd[246]), .B1(i_cmd[230]), .B2(n7765), 
        .B3(n10943), .ZN(n8341) );
  INR4D1BWP30P140LVT U11059 ( .A1(i_cmd[238]), .B1(i_cmd[254]), .B2(n7769), 
        .B3(n7560), .ZN(n8340) );
  AOI22D1BWP30P140LVT U11060 ( .A1(i_data_bus[978]), .A2(n8341), .B1(
        i_data_bus[946]), .B2(n8340), .ZN(n7562) );
  NR3D0P7BWP30P140LVT U11061 ( .A1(i_cmd[246]), .A2(i_cmd[238]), .A3(
        i_cmd[254]), .ZN(n10939) );
  INR4D1BWP30P140LVT U11062 ( .A1(i_cmd[254]), .B1(i_cmd[238]), .B2(n7771), 
        .B3(n7560), .ZN(n8339) );
  AOI22D1BWP30P140LVT U11063 ( .A1(i_data_bus[914]), .A2(n8342), .B1(
        i_data_bus[1010]), .B2(n8339), .ZN(n7561) );
  ND2D1BWP30P140LVT U11064 ( .A1(n7562), .A2(n7561), .ZN(N10273) );
  AOI22D1BWP30P140LVT U11065 ( .A1(i_data_bus[967]), .A2(n8353), .B1(
        i_data_bus[999]), .B2(n8352), .ZN(n7564) );
  AOI22D1BWP30P140LVT U11066 ( .A1(i_data_bus[935]), .A2(n8351), .B1(
        i_data_bus[903]), .B2(n8354), .ZN(n7563) );
  ND2D1BWP30P140LVT U11067 ( .A1(n7564), .A2(n7563), .ZN(N4814) );
  AOI22D1BWP30P140LVT U11068 ( .A1(i_data_bus[961]), .A2(n8353), .B1(
        i_data_bus[993]), .B2(n8352), .ZN(n7566) );
  AOI22D1BWP30P140LVT U11069 ( .A1(i_data_bus[929]), .A2(n8351), .B1(
        i_data_bus[897]), .B2(n8354), .ZN(n7565) );
  ND2D1BWP30P140LVT U11070 ( .A1(n7566), .A2(n7565), .ZN(N4808) );
  AOI22D1BWP30P140LVT U11071 ( .A1(i_data_bus[988]), .A2(n8341), .B1(
        i_data_bus[956]), .B2(n8340), .ZN(n7568) );
  AOI22D1BWP30P140LVT U11072 ( .A1(i_data_bus[1020]), .A2(n8339), .B1(
        i_data_bus[924]), .B2(n8342), .ZN(n7567) );
  ND2D1BWP30P140LVT U11073 ( .A1(n7568), .A2(n7567), .ZN(N10283) );
  AOI22D1BWP30P140LVT U11074 ( .A1(i_data_bus[967]), .A2(n8341), .B1(
        i_data_bus[935]), .B2(n8340), .ZN(n7570) );
  AOI22D1BWP30P140LVT U11075 ( .A1(i_data_bus[999]), .A2(n8339), .B1(
        i_data_bus[903]), .B2(n8342), .ZN(n7569) );
  ND2D1BWP30P140LVT U11076 ( .A1(n7570), .A2(n7569), .ZN(N10262) );
  AOI22D1BWP30P140LVT U11077 ( .A1(i_data_bus[961]), .A2(n8341), .B1(
        i_data_bus[929]), .B2(n8340), .ZN(n7572) );
  AOI22D1BWP30P140LVT U11078 ( .A1(i_data_bus[993]), .A2(n8339), .B1(
        i_data_bus[897]), .B2(n8342), .ZN(n7571) );
  ND2D1BWP30P140LVT U11079 ( .A1(n7572), .A2(n7571), .ZN(N10256) );
  AOI22D1BWP30P140LVT U11080 ( .A1(i_data_bus[984]), .A2(n8341), .B1(
        i_data_bus[1016]), .B2(n8339), .ZN(n7574) );
  AOI22D1BWP30P140LVT U11081 ( .A1(i_data_bus[920]), .A2(n8342), .B1(
        i_data_bus[952]), .B2(n8340), .ZN(n7573) );
  ND2D1BWP30P140LVT U11082 ( .A1(n7574), .A2(n7573), .ZN(N10279) );
  AOI22D1BWP30P140LVT U11083 ( .A1(i_data_bus[973]), .A2(n8341), .B1(
        i_data_bus[1005]), .B2(n8339), .ZN(n7576) );
  AOI22D1BWP30P140LVT U11084 ( .A1(i_data_bus[909]), .A2(n8342), .B1(
        i_data_bus[941]), .B2(n8340), .ZN(n7575) );
  ND2D1BWP30P140LVT U11085 ( .A1(n7576), .A2(n7575), .ZN(N10268) );
  AOI22D1BWP30P140LVT U11086 ( .A1(i_data_bus[968]), .A2(n8341), .B1(
        i_data_bus[1000]), .B2(n8339), .ZN(n7578) );
  AOI22D1BWP30P140LVT U11087 ( .A1(i_data_bus[904]), .A2(n8342), .B1(
        i_data_bus[936]), .B2(n8340), .ZN(n7577) );
  ND2D1BWP30P140LVT U11088 ( .A1(n7578), .A2(n7577), .ZN(N10263) );
  AOI22D1BWP30P140LVT U11089 ( .A1(i_data_bus[968]), .A2(n8353), .B1(
        i_data_bus[904]), .B2(n8354), .ZN(n7580) );
  AOI22D1BWP30P140LVT U11090 ( .A1(i_data_bus[1000]), .A2(n8352), .B1(
        i_data_bus[936]), .B2(n8351), .ZN(n7579) );
  ND2D1BWP30P140LVT U11091 ( .A1(n7580), .A2(n7579), .ZN(N4815) );
  AOI22D1BWP30P140LVT U11092 ( .A1(i_data_bus[971]), .A2(n8341), .B1(
        i_data_bus[907]), .B2(n8342), .ZN(n7582) );
  AOI22D1BWP30P140LVT U11093 ( .A1(i_data_bus[939]), .A2(n8340), .B1(
        i_data_bus[1003]), .B2(n8339), .ZN(n7581) );
  ND2D1BWP30P140LVT U11094 ( .A1(n7582), .A2(n7581), .ZN(N10266) );
  INR4D1BWP30P140LVT U11095 ( .A1(i_cmd[241]), .B1(i_cmd[225]), .B2(n11114), 
        .B3(n7765), .ZN(n8721) );
  NR4D1BWP30P140LVT U11096 ( .A1(i_cmd[233]), .A2(n11116), .A3(n7583), .A4(
        n7771), .ZN(n8719) );
  AOI22D1BWP30P140LVT U11097 ( .A1(i_data_bus[960]), .A2(n8721), .B1(
        i_data_bus[992]), .B2(n8719), .ZN(n7585) );
  NR3D0P7BWP30P140LVT U11098 ( .A1(i_cmd[241]), .A2(i_cmd[233]), .A3(
        i_cmd[249]), .ZN(n11113) );
  AOI22D1BWP30P140LVT U11099 ( .A1(i_data_bus[896]), .A2(n8722), .B1(
        i_data_bus[928]), .B2(n8720), .ZN(n7584) );
  ND2D1BWP30P140LVT U11100 ( .A1(n7585), .A2(n7584), .ZN(N2933) );
  INR4D1BWP30P140LVT U11101 ( .A1(i_cmd[115]), .B1(i_cmd[99]), .B2(n8443), 
        .B3(n11076), .ZN(n7911) );
  NR4D1BWP30P140LVT U11102 ( .A1(i_cmd[107]), .A2(n8447), .A3(n11078), .A4(
        n7586), .ZN(n7909) );
  AOI22D1BWP30P140LVT U11103 ( .A1(i_data_bus[452]), .A2(n7911), .B1(
        i_data_bus[484]), .B2(n7909), .ZN(n7588) );
  NR4D1BWP30P140LVT U11104 ( .A1(i_cmd[123]), .A2(n11079), .A3(n8445), .A4(
        n7586), .ZN(n7910) );
  NR3D0P7BWP30P140LVT U11105 ( .A1(i_cmd[107]), .A2(i_cmd[123]), .A3(
        i_cmd[115]), .ZN(n11075) );
  AOI22D1BWP30P140LVT U11106 ( .A1(i_data_bus[420]), .A2(n7910), .B1(
        i_data_bus[388]), .B2(n6215), .ZN(n7587) );
  ND2D1BWP30P140LVT U11107 ( .A1(n7588), .A2(n7587), .ZN(N5309) );
  AOI22D1BWP30P140LVT U11108 ( .A1(n8721), .A2(i_data_bus[962]), .B1(n8719), 
        .B2(i_data_bus[994]), .ZN(n7590) );
  AOI22D1BWP30P140LVT U11109 ( .A1(n8722), .A2(i_data_bus[898]), .B1(n8720), 
        .B2(i_data_bus[930]), .ZN(n7589) );
  ND2D1BWP30P140LVT U11110 ( .A1(n7590), .A2(n7589), .ZN(N2935) );
  AOI22D1BWP30P140LVT U11111 ( .A1(n8721), .A2(i_data_bus[965]), .B1(n8719), 
        .B2(i_data_bus[997]), .ZN(n7592) );
  AOI22D1BWP30P140LVT U11112 ( .A1(n8722), .A2(i_data_bus[901]), .B1(n8720), 
        .B2(i_data_bus[933]), .ZN(n7591) );
  ND2D1BWP30P140LVT U11113 ( .A1(n7592), .A2(n7591), .ZN(N2938) );
  AOI22D1BWP30P140LVT U11114 ( .A1(n8721), .A2(i_data_bus[970]), .B1(n8719), 
        .B2(i_data_bus[1002]), .ZN(n7594) );
  AOI22D1BWP30P140LVT U11115 ( .A1(n8722), .A2(i_data_bus[906]), .B1(n8720), 
        .B2(i_data_bus[938]), .ZN(n7593) );
  ND2D1BWP30P140LVT U11116 ( .A1(n7594), .A2(n7593), .ZN(N2943) );
  AOI22D1BWP30P140LVT U11117 ( .A1(n8721), .A2(i_data_bus[986]), .B1(n8719), 
        .B2(i_data_bus[1018]), .ZN(n7596) );
  AOI22D1BWP30P140LVT U11118 ( .A1(n8722), .A2(i_data_bus[922]), .B1(n8720), 
        .B2(i_data_bus[954]), .ZN(n7595) );
  ND2D1BWP30P140LVT U11119 ( .A1(n7596), .A2(n7595), .ZN(N2959) );
  AOI22D1BWP30P140LVT U11120 ( .A1(n8721), .A2(i_data_bus[985]), .B1(n8719), 
        .B2(i_data_bus[1017]), .ZN(n7598) );
  AOI22D1BWP30P140LVT U11121 ( .A1(n8722), .A2(i_data_bus[921]), .B1(n8720), 
        .B2(i_data_bus[953]), .ZN(n7597) );
  ND2D1BWP30P140LVT U11122 ( .A1(n7598), .A2(n7597), .ZN(N2958) );
  AOI22D1BWP30P140LVT U11123 ( .A1(n8721), .A2(i_data_bus[984]), .B1(n8719), 
        .B2(i_data_bus[1016]), .ZN(n7600) );
  AOI22D1BWP30P140LVT U11124 ( .A1(n8722), .A2(i_data_bus[920]), .B1(n8720), 
        .B2(i_data_bus[952]), .ZN(n7599) );
  ND2D1BWP30P140LVT U11125 ( .A1(n7600), .A2(n7599), .ZN(N2957) );
  AOI22D1BWP30P140LVT U11126 ( .A1(n8721), .A2(i_data_bus[983]), .B1(n8719), 
        .B2(i_data_bus[1015]), .ZN(n7602) );
  AOI22D1BWP30P140LVT U11127 ( .A1(n8722), .A2(i_data_bus[919]), .B1(n8720), 
        .B2(i_data_bus[951]), .ZN(n7601) );
  ND2D1BWP30P140LVT U11128 ( .A1(n7602), .A2(n7601), .ZN(N2956) );
  AOI22D1BWP30P140LVT U11129 ( .A1(i_data_bus[1006]), .A2(n8205), .B1(
        i_data_bus[942]), .B2(n8208), .ZN(n7604) );
  AOI22D1BWP30P140LVT U11130 ( .A1(i_data_bus[974]), .A2(n8207), .B1(
        i_data_bus[910]), .B2(n8206), .ZN(n7603) );
  ND2D1BWP30P140LVT U11131 ( .A1(n7604), .A2(n7603), .ZN(N5671) );
  AOI22D1BWP30P140LVT U11132 ( .A1(i_data_bus[908]), .A2(n8206), .B1(
        i_data_bus[1004]), .B2(n8205), .ZN(n7606) );
  AOI22D1BWP30P140LVT U11133 ( .A1(i_data_bus[972]), .A2(n8207), .B1(
        i_data_bus[940]), .B2(n8208), .ZN(n7605) );
  ND2D1BWP30P140LVT U11134 ( .A1(n7606), .A2(n7605), .ZN(N5669) );
  AOI22D1BWP30P140LVT U11135 ( .A1(i_data_bus[923]), .A2(n8206), .B1(
        i_data_bus[955]), .B2(n8208), .ZN(n7608) );
  AOI22D1BWP30P140LVT U11136 ( .A1(i_data_bus[987]), .A2(n8207), .B1(
        i_data_bus[1019]), .B2(n8205), .ZN(n7607) );
  ND2D1BWP30P140LVT U11137 ( .A1(n7608), .A2(n7607), .ZN(N5684) );
  AOI22D1BWP30P140LVT U11138 ( .A1(i_data_bus[935]), .A2(n8208), .B1(
        i_data_bus[903]), .B2(n8206), .ZN(n7610) );
  AOI22D1BWP30P140LVT U11139 ( .A1(i_data_bus[967]), .A2(n8207), .B1(
        i_data_bus[999]), .B2(n8205), .ZN(n7609) );
  ND2D1BWP30P140LVT U11140 ( .A1(n7610), .A2(n7609), .ZN(N5664) );
  AOI22D1BWP30P140LVT U11141 ( .A1(i_data_bus[920]), .A2(n8206), .B1(
        i_data_bus[952]), .B2(n8208), .ZN(n7612) );
  AOI22D1BWP30P140LVT U11142 ( .A1(i_data_bus[984]), .A2(n8207), .B1(
        i_data_bus[1016]), .B2(n8205), .ZN(n7611) );
  ND2D1BWP30P140LVT U11143 ( .A1(n7612), .A2(n7611), .ZN(N5681) );
  AOI22D1BWP30P140LVT U11144 ( .A1(i_data_bus[909]), .A2(n8233), .B1(
        i_data_bus[1005]), .B2(n8230), .ZN(n7614) );
  AOI22D1BWP30P140LVT U11145 ( .A1(i_data_bus[973]), .A2(n8232), .B1(
        i_data_bus[941]), .B2(n8231), .ZN(n7613) );
  ND2D1BWP30P140LVT U11146 ( .A1(n7614), .A2(n7613), .ZN(N8394) );
  AOI22D1BWP30P140LVT U11147 ( .A1(i_data_bus[956]), .A2(n8231), .B1(
        i_data_bus[924]), .B2(n8233), .ZN(n7616) );
  AOI22D1BWP30P140LVT U11148 ( .A1(i_data_bus[988]), .A2(n8232), .B1(
        i_data_bus[1020]), .B2(n8230), .ZN(n7615) );
  ND2D1BWP30P140LVT U11149 ( .A1(n7616), .A2(n7615), .ZN(N8409) );
  AOI22D1BWP30P140LVT U11150 ( .A1(i_data_bus[920]), .A2(n8233), .B1(
        i_data_bus[952]), .B2(n8231), .ZN(n7618) );
  AOI22D1BWP30P140LVT U11151 ( .A1(i_data_bus[984]), .A2(n8232), .B1(
        i_data_bus[1016]), .B2(n8230), .ZN(n7617) );
  ND2D1BWP30P140LVT U11152 ( .A1(n7618), .A2(n7617), .ZN(N8405) );
  AOI22D1BWP30P140LVT U11153 ( .A1(i_data_bus[908]), .A2(n8233), .B1(
        i_data_bus[940]), .B2(n8231), .ZN(n7620) );
  AOI22D1BWP30P140LVT U11154 ( .A1(i_data_bus[972]), .A2(n8232), .B1(
        i_data_bus[1004]), .B2(n8230), .ZN(n7619) );
  ND2D1BWP30P140LVT U11155 ( .A1(n7620), .A2(n7619), .ZN(N8393) );
  AOI22D1BWP30P140LVT U11156 ( .A1(i_data_bus[906]), .A2(n8233), .B1(
        i_data_bus[938]), .B2(n8231), .ZN(n7622) );
  AOI22D1BWP30P140LVT U11157 ( .A1(i_data_bus[970]), .A2(n8232), .B1(
        i_data_bus[1002]), .B2(n8230), .ZN(n7621) );
  ND2D1BWP30P140LVT U11158 ( .A1(n7622), .A2(n7621), .ZN(N8391) );
  AOI22D1BWP30P140LVT U11159 ( .A1(i_data_bus[935]), .A2(n8231), .B1(
        i_data_bus[903]), .B2(n8233), .ZN(n7624) );
  AOI22D1BWP30P140LVT U11160 ( .A1(i_data_bus[967]), .A2(n8232), .B1(
        i_data_bus[999]), .B2(n8230), .ZN(n7623) );
  ND2D1BWP30P140LVT U11161 ( .A1(n7624), .A2(n7623), .ZN(N8388) );
  AOI22D1BWP30P140LVT U11162 ( .A1(i_data_bus[901]), .A2(n8233), .B1(
        i_data_bus[933]), .B2(n8231), .ZN(n7626) );
  AOI22D1BWP30P140LVT U11163 ( .A1(i_data_bus[965]), .A2(n8232), .B1(
        i_data_bus[997]), .B2(n8230), .ZN(n7625) );
  ND2D1BWP30P140LVT U11164 ( .A1(n7626), .A2(n7625), .ZN(N8386) );
  NR4D1BWP30P140LVT U11165 ( .A1(i_cmd[109]), .A2(n10994), .A3(n8447), .A4(
        n7627), .ZN(n7826) );
  NR4D1BWP30P140LVT U11166 ( .A1(i_cmd[125]), .A2(n8445), .A3(n10993), .A4(
        n7627), .ZN(n7824) );
  AOI22D1BWP30P140LVT U11167 ( .A1(i_data_bus[506]), .A2(n7826), .B1(
        i_data_bus[442]), .B2(n7824), .ZN(n7629) );
  INR4D1BWP30P140LVT U11168 ( .A1(i_cmd[117]), .B1(i_cmd[101]), .B2(n8443), 
        .B3(n10991), .ZN(n7825) );
  NR3D0P7BWP30P140LVT U11169 ( .A1(i_cmd[117]), .A2(i_cmd[125]), .A3(
        i_cmd[109]), .ZN(n10990) );
  AOI22D1BWP30P140LVT U11170 ( .A1(i_data_bus[474]), .A2(n7825), .B1(
        i_data_bus[410]), .B2(n6214), .ZN(n7628) );
  ND2D1BWP30P140LVT U11171 ( .A1(n7629), .A2(n7628), .ZN(N8055) );
  AOI22D1BWP30P140LVT U11172 ( .A1(i_data_bus[958]), .A2(n8231), .B1(
        i_data_bus[1022]), .B2(n8230), .ZN(n7631) );
  AOI22D1BWP30P140LVT U11173 ( .A1(i_data_bus[990]), .A2(n8232), .B1(
        i_data_bus[926]), .B2(n8233), .ZN(n7630) );
  ND2D1BWP30P140LVT U11174 ( .A1(n7631), .A2(n7630), .ZN(N8411) );
  AOI22D1BWP30P140LVT U11175 ( .A1(i_data_bus[943]), .A2(n8231), .B1(
        i_data_bus[1007]), .B2(n8230), .ZN(n7633) );
  AOI22D1BWP30P140LVT U11176 ( .A1(i_data_bus[975]), .A2(n8232), .B1(
        i_data_bus[911]), .B2(n8233), .ZN(n7632) );
  ND2D1BWP30P140LVT U11177 ( .A1(n7633), .A2(n7632), .ZN(N8396) );
  AOI22D1BWP30P140LVT U11178 ( .A1(i_data_bus[932]), .A2(n8231), .B1(
        i_data_bus[996]), .B2(n8230), .ZN(n7635) );
  AOI22D1BWP30P140LVT U11179 ( .A1(i_data_bus[964]), .A2(n8232), .B1(
        i_data_bus[900]), .B2(n8233), .ZN(n7634) );
  ND2D1BWP30P140LVT U11180 ( .A1(n7635), .A2(n7634), .ZN(N8385) );
  AOI22D1BWP30P140LVT U11181 ( .A1(i_data_bus[999]), .A2(n8255), .B1(
        i_data_bus[903]), .B2(n8258), .ZN(n7637) );
  AOI22D1BWP30P140LVT U11182 ( .A1(i_data_bus[967]), .A2(n8257), .B1(
        i_data_bus[935]), .B2(n8256), .ZN(n7636) );
  ND2D1BWP30P140LVT U11183 ( .A1(n7637), .A2(n7636), .ZN(N11112) );
  AOI22D1BWP30P140LVT U11184 ( .A1(i_data_bus[920]), .A2(n8258), .B1(
        i_data_bus[952]), .B2(n8256), .ZN(n7639) );
  AOI22D1BWP30P140LVT U11185 ( .A1(i_data_bus[984]), .A2(n8257), .B1(
        i_data_bus[1016]), .B2(n8255), .ZN(n7638) );
  ND2D1BWP30P140LVT U11186 ( .A1(n7639), .A2(n7638), .ZN(N11129) );
  AOI22D1BWP30P140LVT U11187 ( .A1(i_data_bus[929]), .A2(n8256), .B1(
        i_data_bus[897]), .B2(n8258), .ZN(n7641) );
  AOI22D1BWP30P140LVT U11188 ( .A1(i_data_bus[961]), .A2(n8257), .B1(
        i_data_bus[993]), .B2(n8255), .ZN(n7640) );
  ND2D1BWP30P140LVT U11189 ( .A1(n7641), .A2(n7640), .ZN(N11106) );
  AOI22D1BWP30P140LVT U11190 ( .A1(i_data_bus[919]), .A2(n8258), .B1(
        i_data_bus[951]), .B2(n8256), .ZN(n7643) );
  AOI22D1BWP30P140LVT U11191 ( .A1(i_data_bus[983]), .A2(n8257), .B1(
        i_data_bus[1015]), .B2(n8255), .ZN(n7642) );
  ND2D1BWP30P140LVT U11192 ( .A1(n7643), .A2(n7642), .ZN(N11128) );
  AOI22D1BWP30P140LVT U11193 ( .A1(i_data_bus[923]), .A2(n8258), .B1(
        i_data_bus[955]), .B2(n8256), .ZN(n7645) );
  AOI22D1BWP30P140LVT U11194 ( .A1(i_data_bus[987]), .A2(n8257), .B1(
        i_data_bus[1019]), .B2(n8255), .ZN(n7644) );
  ND2D1BWP30P140LVT U11195 ( .A1(n7645), .A2(n7644), .ZN(N11132) );
  AOI22D1BWP30P140LVT U11196 ( .A1(i_data_bus[949]), .A2(n8256), .B1(
        i_data_bus[1013]), .B2(n8255), .ZN(n7647) );
  AOI22D1BWP30P140LVT U11197 ( .A1(i_data_bus[981]), .A2(n8257), .B1(
        i_data_bus[917]), .B2(n8258), .ZN(n7646) );
  ND2D1BWP30P140LVT U11198 ( .A1(n7647), .A2(n7646), .ZN(N11126) );
  AOI22D1BWP30P140LVT U11199 ( .A1(i_data_bus[943]), .A2(n8256), .B1(
        i_data_bus[1007]), .B2(n8255), .ZN(n7649) );
  AOI22D1BWP30P140LVT U11200 ( .A1(i_data_bus[975]), .A2(n8257), .B1(
        i_data_bus[911]), .B2(n8258), .ZN(n7648) );
  ND2D1BWP30P140LVT U11201 ( .A1(n7649), .A2(n7648), .ZN(N11120) );
  AOI22D1BWP30P140LVT U11202 ( .A1(i_data_bus[1020]), .A2(n8352), .B1(
        i_data_bus[924]), .B2(n8354), .ZN(n7651) );
  AOI22D1BWP30P140LVT U11203 ( .A1(i_data_bus[988]), .A2(n8353), .B1(
        i_data_bus[956]), .B2(n8351), .ZN(n7650) );
  ND2D1BWP30P140LVT U11204 ( .A1(n7651), .A2(n7650), .ZN(N4835) );
  AOI22D1BWP30P140LVT U11205 ( .A1(i_data_bus[905]), .A2(n8354), .B1(
        i_data_bus[1001]), .B2(n8352), .ZN(n7653) );
  AOI22D1BWP30P140LVT U11206 ( .A1(i_data_bus[969]), .A2(n8353), .B1(
        i_data_bus[937]), .B2(n8351), .ZN(n7652) );
  ND2D1BWP30P140LVT U11207 ( .A1(n7653), .A2(n7652), .ZN(N4816) );
  AOI22D1BWP30P140LVT U11208 ( .A1(i_data_bus[923]), .A2(n8354), .B1(
        i_data_bus[955]), .B2(n8351), .ZN(n7655) );
  AOI22D1BWP30P140LVT U11209 ( .A1(i_data_bus[987]), .A2(n8353), .B1(
        i_data_bus[1019]), .B2(n8352), .ZN(n7654) );
  ND2D1BWP30P140LVT U11210 ( .A1(n7655), .A2(n7654), .ZN(N4834) );
  AOI22D1BWP30P140LVT U11211 ( .A1(i_data_bus[920]), .A2(n8354), .B1(
        i_data_bus[952]), .B2(n8351), .ZN(n7657) );
  AOI22D1BWP30P140LVT U11212 ( .A1(i_data_bus[984]), .A2(n8353), .B1(
        i_data_bus[1016]), .B2(n8352), .ZN(n7656) );
  ND2D1BWP30P140LVT U11213 ( .A1(n7657), .A2(n7656), .ZN(N4831) );
  AOI22D1BWP30P140LVT U11214 ( .A1(i_data_bus[913]), .A2(n8354), .B1(
        i_data_bus[945]), .B2(n8351), .ZN(n7659) );
  AOI22D1BWP30P140LVT U11215 ( .A1(i_data_bus[977]), .A2(n8353), .B1(
        i_data_bus[1009]), .B2(n8352), .ZN(n7658) );
  ND2D1BWP30P140LVT U11216 ( .A1(n7659), .A2(n7658), .ZN(N4824) );
  AOI22D1BWP30P140LVT U11217 ( .A1(i_data_bus[908]), .A2(n8354), .B1(
        i_data_bus[940]), .B2(n8351), .ZN(n7661) );
  AOI22D1BWP30P140LVT U11218 ( .A1(i_data_bus[972]), .A2(n8353), .B1(
        i_data_bus[1004]), .B2(n8352), .ZN(n7660) );
  ND2D1BWP30P140LVT U11219 ( .A1(n7661), .A2(n7660), .ZN(N4819) );
  AOI22D1BWP30P140LVT U11220 ( .A1(i_data_bus[906]), .A2(n8354), .B1(
        i_data_bus[938]), .B2(n8351), .ZN(n7663) );
  AOI22D1BWP30P140LVT U11221 ( .A1(i_data_bus[970]), .A2(n8353), .B1(
        i_data_bus[1002]), .B2(n8352), .ZN(n7662) );
  ND2D1BWP30P140LVT U11222 ( .A1(n7663), .A2(n7662), .ZN(N4817) );
  AOI22D1BWP30P140LVT U11223 ( .A1(i_data_bus[913]), .A2(n8342), .B1(
        i_data_bus[1009]), .B2(n8339), .ZN(n7665) );
  AOI22D1BWP30P140LVT U11224 ( .A1(i_data_bus[977]), .A2(n8341), .B1(
        i_data_bus[945]), .B2(n8340), .ZN(n7664) );
  ND2D1BWP30P140LVT U11225 ( .A1(n7665), .A2(n7664), .ZN(N10272) );
  AOI22D1BWP30P140LVT U11226 ( .A1(i_data_bus[949]), .A2(n8340), .B1(
        i_data_bus[917]), .B2(n8342), .ZN(n7667) );
  AOI22D1BWP30P140LVT U11227 ( .A1(i_data_bus[981]), .A2(n8341), .B1(
        i_data_bus[1013]), .B2(n8339), .ZN(n7666) );
  ND2D1BWP30P140LVT U11228 ( .A1(n7667), .A2(n7666), .ZN(N10276) );
  AOI22D1BWP30P140LVT U11229 ( .A1(i_data_bus[908]), .A2(n8342), .B1(
        i_data_bus[940]), .B2(n8340), .ZN(n7669) );
  AOI22D1BWP30P140LVT U11230 ( .A1(i_data_bus[972]), .A2(n8341), .B1(
        i_data_bus[1004]), .B2(n8339), .ZN(n7668) );
  ND2D1BWP30P140LVT U11231 ( .A1(n7669), .A2(n7668), .ZN(N10267) );
  AOI22D1BWP30P140LVT U11232 ( .A1(i_data_bus[905]), .A2(n8342), .B1(
        i_data_bus[937]), .B2(n8340), .ZN(n7671) );
  AOI22D1BWP30P140LVT U11233 ( .A1(i_data_bus[969]), .A2(n8341), .B1(
        i_data_bus[1001]), .B2(n8339), .ZN(n7670) );
  ND2D1BWP30P140LVT U11234 ( .A1(n7671), .A2(n7670), .ZN(N10264) );
  AOI22D1BWP30P140LVT U11235 ( .A1(i_data_bus[901]), .A2(n8342), .B1(
        i_data_bus[933]), .B2(n8340), .ZN(n7673) );
  AOI22D1BWP30P140LVT U11236 ( .A1(i_data_bus[965]), .A2(n8341), .B1(
        i_data_bus[997]), .B2(n8339), .ZN(n7672) );
  ND2D1BWP30P140LVT U11237 ( .A1(n7673), .A2(n7672), .ZN(N10260) );
  AOI22D1BWP30P140LVT U11238 ( .A1(i_data_bus[934]), .A2(n8340), .B1(
        i_data_bus[998]), .B2(n8339), .ZN(n7675) );
  AOI22D1BWP30P140LVT U11239 ( .A1(i_data_bus[966]), .A2(n8341), .B1(
        i_data_bus[902]), .B2(n8342), .ZN(n7674) );
  ND2D1BWP30P140LVT U11240 ( .A1(n7675), .A2(n7674), .ZN(N10261) );
  AOI22D1BWP30P140LVT U11241 ( .A1(i_data_bus[958]), .A2(n8351), .B1(
        i_data_bus[1022]), .B2(n8352), .ZN(n7677) );
  AOI22D1BWP30P140LVT U11242 ( .A1(i_data_bus[990]), .A2(n8353), .B1(
        i_data_bus[926]), .B2(n8354), .ZN(n7676) );
  ND2D1BWP30P140LVT U11243 ( .A1(n7677), .A2(n7676), .ZN(N4837) );
  AOI22D1BWP30P140LVT U11244 ( .A1(i_data_bus[949]), .A2(n8351), .B1(
        i_data_bus[1013]), .B2(n8352), .ZN(n7679) );
  AOI22D1BWP30P140LVT U11245 ( .A1(i_data_bus[981]), .A2(n8353), .B1(
        i_data_bus[917]), .B2(n8354), .ZN(n7678) );
  ND2D1BWP30P140LVT U11246 ( .A1(n7679), .A2(n7678), .ZN(N4828) );
  AOI22D1BWP30P140LVT U11247 ( .A1(i_data_bus[485]), .A2(n7909), .B1(
        i_data_bus[453]), .B2(n7911), .ZN(n7681) );
  AOI22D1BWP30P140LVT U11248 ( .A1(i_data_bus[421]), .A2(n7910), .B1(
        i_data_bus[389]), .B2(n6215), .ZN(n7680) );
  ND2D1BWP30P140LVT U11249 ( .A1(n7681), .A2(n7680), .ZN(N5310) );
  AOI22D1BWP30P140LVT U11250 ( .A1(i_data_bus[490]), .A2(n7909), .B1(
        i_data_bus[458]), .B2(n7911), .ZN(n7683) );
  AOI22D1BWP30P140LVT U11251 ( .A1(i_data_bus[426]), .A2(n7910), .B1(
        i_data_bus[394]), .B2(n6215), .ZN(n7682) );
  ND2D1BWP30P140LVT U11252 ( .A1(n7683), .A2(n7682), .ZN(N5315) );
  AOI22D1BWP30P140LVT U11253 ( .A1(i_data_bus[416]), .A2(n7824), .B1(
        i_data_bus[480]), .B2(n7826), .ZN(n7685) );
  AOI22D1BWP30P140LVT U11254 ( .A1(i_data_bus[448]), .A2(n7825), .B1(
        i_data_bus[384]), .B2(n6214), .ZN(n7684) );
  ND2D1BWP30P140LVT U11255 ( .A1(n7685), .A2(n7684), .ZN(N8029) );
  AOI22D1BWP30P140LVT U11256 ( .A1(i_data_bus[508]), .A2(n7826), .B1(
        i_data_bus[476]), .B2(n7825), .ZN(n7687) );
  AOI22D1BWP30P140LVT U11257 ( .A1(i_data_bus[444]), .A2(n7824), .B1(
        i_data_bus[412]), .B2(n6214), .ZN(n7686) );
  ND2D1BWP30P140LVT U11258 ( .A1(n7687), .A2(n7686), .ZN(N8057) );
  AOI22D1BWP30P140LVT U11259 ( .A1(i_data_bus[451]), .A2(n7911), .B1(
        i_data_bus[387]), .B2(n6215), .ZN(n7689) );
  AOI22D1BWP30P140LVT U11260 ( .A1(i_data_bus[419]), .A2(n7910), .B1(
        i_data_bus[483]), .B2(n7909), .ZN(n7688) );
  ND2D1BWP30P140LVT U11261 ( .A1(n7689), .A2(n7688), .ZN(N5308) );
  AOI22D1BWP30P140LVT U11262 ( .A1(i_data_bus[498]), .A2(n7826), .B1(
        i_data_bus[466]), .B2(n7825), .ZN(n7691) );
  AOI22D1BWP30P140LVT U11263 ( .A1(i_data_bus[434]), .A2(n7824), .B1(
        i_data_bus[402]), .B2(n6214), .ZN(n7690) );
  ND2D1BWP30P140LVT U11264 ( .A1(n7691), .A2(n7690), .ZN(N8047) );
  AOI22D1BWP30P140LVT U11265 ( .A1(i_data_bus[412]), .A2(n6215), .B1(
        i_data_bus[476]), .B2(n7911), .ZN(n7693) );
  AOI22D1BWP30P140LVT U11266 ( .A1(i_data_bus[444]), .A2(n7910), .B1(
        i_data_bus[508]), .B2(n7909), .ZN(n7692) );
  ND2D1BWP30P140LVT U11267 ( .A1(n7693), .A2(n7692), .ZN(N5333) );
  AOI22D1BWP30P140LVT U11268 ( .A1(i_data_bus[396]), .A2(n6215), .B1(
        i_data_bus[460]), .B2(n7911), .ZN(n7695) );
  AOI22D1BWP30P140LVT U11269 ( .A1(i_data_bus[428]), .A2(n7910), .B1(
        i_data_bus[492]), .B2(n7909), .ZN(n7694) );
  ND2D1BWP30P140LVT U11270 ( .A1(n7695), .A2(n7694), .ZN(N5317) );
  AOI22D1BWP30P140LVT U11271 ( .A1(i_data_bus[416]), .A2(n7910), .B1(
        i_data_bus[384]), .B2(n6215), .ZN(n7697) );
  AOI22D1BWP30P140LVT U11272 ( .A1(i_data_bus[448]), .A2(n7911), .B1(
        i_data_bus[480]), .B2(n7909), .ZN(n7696) );
  ND2D1BWP30P140LVT U11273 ( .A1(n7697), .A2(n7696), .ZN(N5305) );
  AOI22D1BWP30P140LVT U11274 ( .A1(i_data_bus[457]), .A2(n7911), .B1(
        i_data_bus[393]), .B2(n6215), .ZN(n7699) );
  AOI22D1BWP30P140LVT U11275 ( .A1(i_data_bus[425]), .A2(n7910), .B1(
        i_data_bus[489]), .B2(n7909), .ZN(n7698) );
  ND2D1BWP30P140LVT U11276 ( .A1(n7699), .A2(n7698), .ZN(N5314) );
  AOI22D1BWP30P140LVT U11277 ( .A1(n8722), .A2(i_data_bus[904]), .B1(n8720), 
        .B2(i_data_bus[936]), .ZN(n7701) );
  AOI22D1BWP30P140LVT U11278 ( .A1(n8721), .A2(i_data_bus[968]), .B1(n8719), 
        .B2(i_data_bus[1000]), .ZN(n7700) );
  ND2D1BWP30P140LVT U11279 ( .A1(n7701), .A2(n7700), .ZN(N2941) );
  AOI22D1BWP30P140LVT U11280 ( .A1(n8722), .A2(i_data_bus[910]), .B1(n8720), 
        .B2(i_data_bus[942]), .ZN(n7703) );
  AOI22D1BWP30P140LVT U11281 ( .A1(n8721), .A2(i_data_bus[974]), .B1(n8719), 
        .B2(i_data_bus[1006]), .ZN(n7702) );
  ND2D1BWP30P140LVT U11282 ( .A1(n7703), .A2(n7702), .ZN(N2947) );
  AOI22D1BWP30P140LVT U11283 ( .A1(n8722), .A2(i_data_bus[924]), .B1(n8720), 
        .B2(i_data_bus[956]), .ZN(n7705) );
  AOI22D1BWP30P140LVT U11284 ( .A1(n8721), .A2(i_data_bus[988]), .B1(n8719), 
        .B2(i_data_bus[1020]), .ZN(n7704) );
  ND2D1BWP30P140LVT U11285 ( .A1(n7705), .A2(n7704), .ZN(N2961) );
  AOI22D1BWP30P140LVT U11286 ( .A1(i_data_bus[479]), .A2(n7825), .B1(
        i_data_bus[415]), .B2(n6214), .ZN(n7707) );
  AOI22D1BWP30P140LVT U11287 ( .A1(i_data_bus[511]), .A2(n7826), .B1(
        i_data_bus[447]), .B2(n7824), .ZN(n7706) );
  ND2D1BWP30P140LVT U11288 ( .A1(n7707), .A2(n7706), .ZN(N8060) );
  AOI22D1BWP30P140LVT U11289 ( .A1(i_data_bus[414]), .A2(n6214), .B1(
        i_data_bus[510]), .B2(n7826), .ZN(n7709) );
  AOI22D1BWP30P140LVT U11290 ( .A1(i_data_bus[478]), .A2(n7825), .B1(
        i_data_bus[446]), .B2(n7824), .ZN(n7708) );
  ND2D1BWP30P140LVT U11291 ( .A1(n7709), .A2(n7708), .ZN(N8059) );
  AOI22D1BWP30P140LVT U11292 ( .A1(i_data_bus[509]), .A2(n7826), .B1(
        i_data_bus[477]), .B2(n7825), .ZN(n7711) );
  AOI22D1BWP30P140LVT U11293 ( .A1(i_data_bus[413]), .A2(n6214), .B1(
        i_data_bus[445]), .B2(n7824), .ZN(n7710) );
  ND2D1BWP30P140LVT U11294 ( .A1(n7711), .A2(n7710), .ZN(N8058) );
  AOI22D1BWP30P140LVT U11295 ( .A1(i_data_bus[507]), .A2(n7826), .B1(
        i_data_bus[475]), .B2(n7825), .ZN(n7713) );
  AOI22D1BWP30P140LVT U11296 ( .A1(i_data_bus[411]), .A2(n6214), .B1(
        i_data_bus[443]), .B2(n7824), .ZN(n7712) );
  ND2D1BWP30P140LVT U11297 ( .A1(n7713), .A2(n7712), .ZN(N8056) );
  AOI22D1BWP30P140LVT U11298 ( .A1(i_data_bus[505]), .A2(n7826), .B1(
        i_data_bus[473]), .B2(n7825), .ZN(n7715) );
  AOI22D1BWP30P140LVT U11299 ( .A1(i_data_bus[409]), .A2(n6214), .B1(
        i_data_bus[441]), .B2(n7824), .ZN(n7714) );
  ND2D1BWP30P140LVT U11300 ( .A1(n7715), .A2(n7714), .ZN(N8054) );
  AOI22D1BWP30P140LVT U11301 ( .A1(i_data_bus[501]), .A2(n7826), .B1(
        i_data_bus[469]), .B2(n7825), .ZN(n7717) );
  AOI22D1BWP30P140LVT U11302 ( .A1(i_data_bus[405]), .A2(n6214), .B1(
        i_data_bus[437]), .B2(n7824), .ZN(n7716) );
  ND2D1BWP30P140LVT U11303 ( .A1(n7717), .A2(n7716), .ZN(N8050) );
  AOI22D1BWP30P140LVT U11304 ( .A1(i_data_bus[496]), .A2(n7826), .B1(
        i_data_bus[464]), .B2(n7825), .ZN(n7719) );
  AOI22D1BWP30P140LVT U11305 ( .A1(i_data_bus[400]), .A2(n6214), .B1(
        i_data_bus[432]), .B2(n7824), .ZN(n7718) );
  ND2D1BWP30P140LVT U11306 ( .A1(n7719), .A2(n7718), .ZN(N8045) );
  AOI22D1BWP30P140LVT U11307 ( .A1(i_data_bus[495]), .A2(n7826), .B1(
        i_data_bus[399]), .B2(n6214), .ZN(n7721) );
  AOI22D1BWP30P140LVT U11308 ( .A1(i_data_bus[463]), .A2(n7825), .B1(
        i_data_bus[431]), .B2(n7824), .ZN(n7720) );
  ND2D1BWP30P140LVT U11309 ( .A1(n7721), .A2(n7720), .ZN(N8044) );
  AOI22D1BWP30P140LVT U11310 ( .A1(i_data_bus[395]), .A2(n6214), .B1(
        i_data_bus[491]), .B2(n7826), .ZN(n7723) );
  AOI22D1BWP30P140LVT U11311 ( .A1(i_data_bus[459]), .A2(n7825), .B1(
        i_data_bus[427]), .B2(n7824), .ZN(n7722) );
  ND2D1BWP30P140LVT U11312 ( .A1(n7723), .A2(n7722), .ZN(N8040) );
  AOI22D1BWP30P140LVT U11313 ( .A1(i_data_bus[456]), .A2(n7825), .B1(
        i_data_bus[392]), .B2(n6214), .ZN(n7725) );
  AOI22D1BWP30P140LVT U11314 ( .A1(i_data_bus[488]), .A2(n7826), .B1(
        i_data_bus[424]), .B2(n7824), .ZN(n7724) );
  ND2D1BWP30P140LVT U11315 ( .A1(n7725), .A2(n7724), .ZN(N8037) );
  AOI22D1BWP30P140LVT U11316 ( .A1(i_data_bus[388]), .A2(n6214), .B1(
        i_data_bus[484]), .B2(n7826), .ZN(n7727) );
  AOI22D1BWP30P140LVT U11317 ( .A1(i_data_bus[452]), .A2(n7825), .B1(
        i_data_bus[420]), .B2(n7824), .ZN(n7726) );
  ND2D1BWP30P140LVT U11318 ( .A1(n7727), .A2(n7726), .ZN(N8033) );
  AOI22D1BWP30P140LVT U11319 ( .A1(i_data_bus[386]), .A2(n6214), .B1(
        i_data_bus[450]), .B2(n7825), .ZN(n7729) );
  AOI22D1BWP30P140LVT U11320 ( .A1(i_data_bus[482]), .A2(n7826), .B1(
        i_data_bus[418]), .B2(n7824), .ZN(n7728) );
  ND2D1BWP30P140LVT U11321 ( .A1(n7729), .A2(n7728), .ZN(N8031) );
  AOI22D1BWP30P140LVT U11322 ( .A1(i_data_bus[481]), .A2(n7826), .B1(
        i_data_bus[385]), .B2(n6214), .ZN(n7731) );
  AOI22D1BWP30P140LVT U11323 ( .A1(i_data_bus[449]), .A2(n7825), .B1(
        i_data_bus[417]), .B2(n7824), .ZN(n7730) );
  ND2D1BWP30P140LVT U11324 ( .A1(n7731), .A2(n7730), .ZN(N8030) );
  AOI22D1BWP30P140LVT U11325 ( .A1(i_data_bus[974]), .A2(n9544), .B1(
        i_data_bus[910]), .B2(n6226), .ZN(n7737) );
  AOI22D1BWP30P140LVT U11326 ( .A1(i_data_bus[1006]), .A2(n9543), .B1(
        i_data_bus[942]), .B2(n9545), .ZN(n7736) );
  ND2D1BWP30P140LVT U11327 ( .A1(n7737), .A2(n7736), .ZN(N2097) );
  AOI22D1BWP30P140LVT U11328 ( .A1(i_data_bus[961]), .A2(n9544), .B1(
        i_data_bus[897]), .B2(n6226), .ZN(n7739) );
  AOI22D1BWP30P140LVT U11329 ( .A1(i_data_bus[929]), .A2(n9545), .B1(
        i_data_bus[993]), .B2(n9543), .ZN(n7738) );
  ND2D1BWP30P140LVT U11330 ( .A1(n7739), .A2(n7738), .ZN(N2084) );
  AOI22D1BWP30P140LVT U11331 ( .A1(i_data_bus[975]), .A2(n9544), .B1(
        i_data_bus[911]), .B2(n6226), .ZN(n7741) );
  AOI22D1BWP30P140LVT U11332 ( .A1(i_data_bus[943]), .A2(n9545), .B1(
        i_data_bus[1007]), .B2(n9543), .ZN(n7740) );
  ND2D1BWP30P140LVT U11333 ( .A1(n7741), .A2(n7740), .ZN(N2098) );
  AOI22D1BWP30P140LVT U11334 ( .A1(i_data_bus[967]), .A2(n9544), .B1(
        i_data_bus[935]), .B2(n9545), .ZN(n7743) );
  AOI22D1BWP30P140LVT U11335 ( .A1(i_data_bus[999]), .A2(n9543), .B1(
        i_data_bus[903]), .B2(n6226), .ZN(n7742) );
  ND2D1BWP30P140LVT U11336 ( .A1(n7743), .A2(n7742), .ZN(N2090) );
  AOI22D1BWP30P140LVT U11337 ( .A1(i_data_bus[988]), .A2(n9544), .B1(
        i_data_bus[956]), .B2(n9545), .ZN(n7745) );
  AOI22D1BWP30P140LVT U11338 ( .A1(i_data_bus[1020]), .A2(n9543), .B1(
        i_data_bus[924]), .B2(n6226), .ZN(n7744) );
  ND2D1BWP30P140LVT U11339 ( .A1(n7745), .A2(n7744), .ZN(N2111) );
  AOI22D1BWP30P140LVT U11340 ( .A1(i_data_bus[479]), .A2(n7911), .B1(
        i_data_bus[447]), .B2(n7910), .ZN(n7747) );
  AOI22D1BWP30P140LVT U11341 ( .A1(i_data_bus[511]), .A2(n7909), .B1(
        i_data_bus[415]), .B2(n6215), .ZN(n7746) );
  ND2D1BWP30P140LVT U11342 ( .A1(n7747), .A2(n7746), .ZN(N5336) );
  AOI22D1BWP30P140LVT U11343 ( .A1(i_data_bus[507]), .A2(n7909), .B1(
        i_data_bus[443]), .B2(n7910), .ZN(n7749) );
  AOI22D1BWP30P140LVT U11344 ( .A1(i_data_bus[475]), .A2(n7911), .B1(
        i_data_bus[411]), .B2(n6215), .ZN(n7748) );
  ND2D1BWP30P140LVT U11345 ( .A1(n7749), .A2(n7748), .ZN(N5332) );
  AOI22D1BWP30P140LVT U11346 ( .A1(i_data_bus[488]), .A2(n7909), .B1(
        i_data_bus[424]), .B2(n7910), .ZN(n7751) );
  AOI22D1BWP30P140LVT U11347 ( .A1(i_data_bus[456]), .A2(n7911), .B1(
        i_data_bus[392]), .B2(n6215), .ZN(n7750) );
  ND2D1BWP30P140LVT U11348 ( .A1(n7751), .A2(n7750), .ZN(N5313) );
  AOI22D1BWP30P140LVT U11349 ( .A1(i_data_bus[962]), .A2(n9544), .B1(
        i_data_bus[994]), .B2(n9543), .ZN(n7753) );
  AOI22D1BWP30P140LVT U11350 ( .A1(i_data_bus[898]), .A2(n6226), .B1(
        i_data_bus[930]), .B2(n9545), .ZN(n7752) );
  ND2D1BWP30P140LVT U11351 ( .A1(n7753), .A2(n7752), .ZN(N2085) );
  AOI22D1BWP30P140LVT U11352 ( .A1(i_data_bus[395]), .A2(n6215), .B1(
        i_data_bus[427]), .B2(n7910), .ZN(n7755) );
  AOI22D1BWP30P140LVT U11353 ( .A1(i_data_bus[459]), .A2(n7911), .B1(
        i_data_bus[491]), .B2(n7909), .ZN(n7754) );
  ND2D1BWP30P140LVT U11354 ( .A1(n7755), .A2(n7754), .ZN(N5316) );
  AOI22D1BWP30P140LVT U11355 ( .A1(i_data_bus[391]), .A2(n6215), .B1(
        i_data_bus[423]), .B2(n7910), .ZN(n7757) );
  AOI22D1BWP30P140LVT U11356 ( .A1(i_data_bus[455]), .A2(n7911), .B1(
        i_data_bus[487]), .B2(n7909), .ZN(n7756) );
  ND2D1BWP30P140LVT U11357 ( .A1(n7757), .A2(n7756), .ZN(N5312) );
  AOI22D1BWP30P140LVT U11358 ( .A1(i_data_bus[414]), .A2(n6215), .B1(
        i_data_bus[446]), .B2(n7910), .ZN(n7759) );
  AOI22D1BWP30P140LVT U11359 ( .A1(i_data_bus[478]), .A2(n7911), .B1(
        i_data_bus[510]), .B2(n7909), .ZN(n7758) );
  ND2D1BWP30P140LVT U11360 ( .A1(n7759), .A2(n7758), .ZN(N5335) );
  AOI22D1BWP30P140LVT U11361 ( .A1(i_data_bus[471]), .A2(n7911), .B1(
        i_data_bus[439]), .B2(n7910), .ZN(n7761) );
  AOI22D1BWP30P140LVT U11362 ( .A1(i_data_bus[407]), .A2(n6215), .B1(
        i_data_bus[503]), .B2(n7909), .ZN(n7760) );
  ND2D1BWP30P140LVT U11363 ( .A1(n7761), .A2(n7760), .ZN(N5328) );
  AOI22D1BWP30P140LVT U11364 ( .A1(i_data_bus[399]), .A2(n6215), .B1(
        i_data_bus[431]), .B2(n7910), .ZN(n7763) );
  AOI22D1BWP30P140LVT U11365 ( .A1(i_data_bus[463]), .A2(n7911), .B1(
        i_data_bus[495]), .B2(n7909), .ZN(n7762) );
  ND2D1BWP30P140LVT U11366 ( .A1(n7763), .A2(n7762), .ZN(N5320) );
  AOI22D1BWP30P140LVT U11367 ( .A1(i_data_bus[981]), .A2(n9662), .B1(
        i_data_bus[917]), .B2(n9661), .ZN(n7773) );
  AOI22D1BWP30P140LVT U11368 ( .A1(i_data_bus[949]), .A2(n9660), .B1(
        i_data_bus[1013]), .B2(n9663), .ZN(n7772) );
  ND2D1BWP30P140LVT U11369 ( .A1(n7773), .A2(n7772), .ZN(N7552) );
  AOI22D1BWP30P140LVT U11370 ( .A1(i_data_bus[972]), .A2(n9662), .B1(
        i_data_bus[940]), .B2(n9660), .ZN(n7775) );
  AOI22D1BWP30P140LVT U11371 ( .A1(i_data_bus[908]), .A2(n9661), .B1(
        i_data_bus[1004]), .B2(n9663), .ZN(n7774) );
  ND2D1BWP30P140LVT U11372 ( .A1(n7775), .A2(n7774), .ZN(N7543) );
  AOI22D1BWP30P140LVT U11373 ( .A1(i_data_bus[969]), .A2(n9662), .B1(
        i_data_bus[937]), .B2(n9660), .ZN(n7777) );
  AOI22D1BWP30P140LVT U11374 ( .A1(i_data_bus[905]), .A2(n9661), .B1(
        i_data_bus[1001]), .B2(n9663), .ZN(n7776) );
  ND2D1BWP30P140LVT U11375 ( .A1(n7777), .A2(n7776), .ZN(N7540) );
  AOI22D1BWP30P140LVT U11376 ( .A1(i_data_bus[973]), .A2(n9662), .B1(
        i_data_bus[1005]), .B2(n9663), .ZN(n7779) );
  AOI22D1BWP30P140LVT U11377 ( .A1(i_data_bus[909]), .A2(n9661), .B1(
        i_data_bus[941]), .B2(n9660), .ZN(n7778) );
  ND2D1BWP30P140LVT U11378 ( .A1(n7779), .A2(n7778), .ZN(N7544) );
  AOI22D1BWP30P140LVT U11379 ( .A1(i_data_bus[390]), .A2(n6215), .B1(
        i_data_bus[422]), .B2(n7910), .ZN(n7781) );
  AOI22D1BWP30P140LVT U11380 ( .A1(i_data_bus[486]), .A2(n7909), .B1(
        i_data_bus[454]), .B2(n7911), .ZN(n7780) );
  ND2D1BWP30P140LVT U11381 ( .A1(n7781), .A2(n7780), .ZN(N5311) );
  AOI22D1BWP30P140LVT U11382 ( .A1(i_data_bus[409]), .A2(n6215), .B1(
        i_data_bus[505]), .B2(n7909), .ZN(n7783) );
  AOI22D1BWP30P140LVT U11383 ( .A1(i_data_bus[441]), .A2(n7910), .B1(
        i_data_bus[473]), .B2(n7911), .ZN(n7782) );
  ND2D1BWP30P140LVT U11384 ( .A1(n7783), .A2(n7782), .ZN(N5330) );
  AOI22D1BWP30P140LVT U11385 ( .A1(i_data_bus[504]), .A2(n7909), .B1(
        i_data_bus[408]), .B2(n6215), .ZN(n7785) );
  AOI22D1BWP30P140LVT U11386 ( .A1(i_data_bus[440]), .A2(n7910), .B1(
        i_data_bus[472]), .B2(n7911), .ZN(n7784) );
  ND2D1BWP30P140LVT U11387 ( .A1(n7785), .A2(n7784), .ZN(N5329) );
  AOI22D1BWP30P140LVT U11388 ( .A1(i_data_bus[404]), .A2(n6215), .B1(
        i_data_bus[500]), .B2(n7909), .ZN(n7787) );
  AOI22D1BWP30P140LVT U11389 ( .A1(i_data_bus[436]), .A2(n7910), .B1(
        i_data_bus[468]), .B2(n7911), .ZN(n7786) );
  ND2D1BWP30P140LVT U11390 ( .A1(n7787), .A2(n7786), .ZN(N5325) );
  AOI22D1BWP30P140LVT U11391 ( .A1(i_data_bus[434]), .A2(n7910), .B1(
        i_data_bus[402]), .B2(n6215), .ZN(n7789) );
  AOI22D1BWP30P140LVT U11392 ( .A1(i_data_bus[498]), .A2(n7909), .B1(
        i_data_bus[466]), .B2(n7911), .ZN(n7788) );
  ND2D1BWP30P140LVT U11393 ( .A1(n7789), .A2(n7788), .ZN(N5323) );
  AOI22D1BWP30P140LVT U11394 ( .A1(i_data_bus[400]), .A2(n6215), .B1(
        i_data_bus[432]), .B2(n7910), .ZN(n7791) );
  AOI22D1BWP30P140LVT U11395 ( .A1(i_data_bus[496]), .A2(n7909), .B1(
        i_data_bus[464]), .B2(n7911), .ZN(n7790) );
  ND2D1BWP30P140LVT U11396 ( .A1(n7791), .A2(n7790), .ZN(N5321) );
  AOI22D1BWP30P140LVT U11397 ( .A1(i_data_bus[430]), .A2(n7910), .B1(
        i_data_bus[494]), .B2(n7909), .ZN(n7793) );
  AOI22D1BWP30P140LVT U11398 ( .A1(i_data_bus[398]), .A2(n6215), .B1(
        i_data_bus[462]), .B2(n7911), .ZN(n7792) );
  ND2D1BWP30P140LVT U11399 ( .A1(n7793), .A2(n7792), .ZN(N5319) );
  AOI22D1BWP30P140LVT U11400 ( .A1(i_data_bus[482]), .A2(n7909), .B1(
        i_data_bus[418]), .B2(n7910), .ZN(n7795) );
  AOI22D1BWP30P140LVT U11401 ( .A1(i_data_bus[386]), .A2(n6215), .B1(
        i_data_bus[450]), .B2(n7911), .ZN(n7794) );
  ND2D1BWP30P140LVT U11402 ( .A1(n7795), .A2(n7794), .ZN(N5307) );
  AOI22D1BWP30P140LVT U11403 ( .A1(i_data_bus[407]), .A2(n6214), .B1(
        i_data_bus[471]), .B2(n7825), .ZN(n7797) );
  AOI22D1BWP30P140LVT U11404 ( .A1(i_data_bus[439]), .A2(n7824), .B1(
        i_data_bus[503]), .B2(n7826), .ZN(n7796) );
  ND2D1BWP30P140LVT U11405 ( .A1(n7797), .A2(n7796), .ZN(N8052) );
  AOI22D1BWP30P140LVT U11406 ( .A1(i_data_bus[404]), .A2(n6214), .B1(
        i_data_bus[468]), .B2(n7825), .ZN(n7799) );
  AOI22D1BWP30P140LVT U11407 ( .A1(i_data_bus[436]), .A2(n7824), .B1(
        i_data_bus[500]), .B2(n7826), .ZN(n7798) );
  ND2D1BWP30P140LVT U11408 ( .A1(n7799), .A2(n7798), .ZN(N8049) );
  AOI22D1BWP30P140LVT U11409 ( .A1(i_data_bus[465]), .A2(n7825), .B1(
        i_data_bus[433]), .B2(n7824), .ZN(n7801) );
  AOI22D1BWP30P140LVT U11410 ( .A1(i_data_bus[401]), .A2(n6214), .B1(
        i_data_bus[497]), .B2(n7826), .ZN(n7800) );
  ND2D1BWP30P140LVT U11411 ( .A1(n7801), .A2(n7800), .ZN(N8046) );
  AOI22D1BWP30P140LVT U11412 ( .A1(i_data_bus[461]), .A2(n7825), .B1(
        i_data_bus[429]), .B2(n7824), .ZN(n7803) );
  AOI22D1BWP30P140LVT U11413 ( .A1(i_data_bus[397]), .A2(n6214), .B1(
        i_data_bus[493]), .B2(n7826), .ZN(n7802) );
  ND2D1BWP30P140LVT U11414 ( .A1(n7803), .A2(n7802), .ZN(N8042) );
  AOI22D1BWP30P140LVT U11415 ( .A1(i_data_bus[457]), .A2(n7825), .B1(
        i_data_bus[393]), .B2(n6214), .ZN(n7805) );
  AOI22D1BWP30P140LVT U11416 ( .A1(i_data_bus[425]), .A2(n7824), .B1(
        i_data_bus[489]), .B2(n7826), .ZN(n7804) );
  ND2D1BWP30P140LVT U11417 ( .A1(n7805), .A2(n7804), .ZN(N8038) );
  AOI22D1BWP30P140LVT U11418 ( .A1(i_data_bus[391]), .A2(n6214), .B1(
        i_data_bus[423]), .B2(n7824), .ZN(n7807) );
  AOI22D1BWP30P140LVT U11419 ( .A1(i_data_bus[455]), .A2(n7825), .B1(
        i_data_bus[487]), .B2(n7826), .ZN(n7806) );
  ND2D1BWP30P140LVT U11420 ( .A1(n7807), .A2(n7806), .ZN(N8036) );
  AOI22D1BWP30P140LVT U11421 ( .A1(i_data_bus[390]), .A2(n6214), .B1(
        i_data_bus[454]), .B2(n7825), .ZN(n7809) );
  AOI22D1BWP30P140LVT U11422 ( .A1(i_data_bus[422]), .A2(n7824), .B1(
        i_data_bus[486]), .B2(n7826), .ZN(n7808) );
  ND2D1BWP30P140LVT U11423 ( .A1(n7809), .A2(n7808), .ZN(N8035) );
  AOI22D1BWP30P140LVT U11424 ( .A1(i_data_bus[451]), .A2(n7825), .B1(
        i_data_bus[387]), .B2(n6214), .ZN(n7811) );
  AOI22D1BWP30P140LVT U11425 ( .A1(i_data_bus[419]), .A2(n7824), .B1(
        i_data_bus[483]), .B2(n7826), .ZN(n7810) );
  ND2D1BWP30P140LVT U11426 ( .A1(n7811), .A2(n7810), .ZN(N8032) );
  AOI22D1BWP30P140LVT U11427 ( .A1(i_data_bus[440]), .A2(n7824), .B1(
        i_data_bus[504]), .B2(n7826), .ZN(n7813) );
  AOI22D1BWP30P140LVT U11428 ( .A1(i_data_bus[408]), .A2(n6214), .B1(
        i_data_bus[472]), .B2(n7825), .ZN(n7812) );
  ND2D1BWP30P140LVT U11429 ( .A1(n7813), .A2(n7812), .ZN(N8053) );
  AOI22D1BWP30P140LVT U11430 ( .A1(i_data_bus[502]), .A2(n7826), .B1(
        i_data_bus[406]), .B2(n6214), .ZN(n7815) );
  AOI22D1BWP30P140LVT U11431 ( .A1(i_data_bus[438]), .A2(n7824), .B1(
        i_data_bus[470]), .B2(n7825), .ZN(n7814) );
  ND2D1BWP30P140LVT U11432 ( .A1(n7815), .A2(n7814), .ZN(N8051) );
  AOI22D1BWP30P140LVT U11433 ( .A1(i_data_bus[435]), .A2(n7824), .B1(
        i_data_bus[499]), .B2(n7826), .ZN(n7817) );
  AOI22D1BWP30P140LVT U11434 ( .A1(i_data_bus[403]), .A2(n6214), .B1(
        i_data_bus[467]), .B2(n7825), .ZN(n7816) );
  ND2D1BWP30P140LVT U11435 ( .A1(n7817), .A2(n7816), .ZN(N8048) );
  AOI22D1BWP30P140LVT U11436 ( .A1(i_data_bus[398]), .A2(n6214), .B1(
        i_data_bus[494]), .B2(n7826), .ZN(n7819) );
  AOI22D1BWP30P140LVT U11437 ( .A1(i_data_bus[430]), .A2(n7824), .B1(
        i_data_bus[462]), .B2(n7825), .ZN(n7818) );
  ND2D1BWP30P140LVT U11438 ( .A1(n7819), .A2(n7818), .ZN(N8043) );
  AOI22D1BWP30P140LVT U11439 ( .A1(i_data_bus[428]), .A2(n7824), .B1(
        i_data_bus[396]), .B2(n6214), .ZN(n7821) );
  AOI22D1BWP30P140LVT U11440 ( .A1(i_data_bus[492]), .A2(n7826), .B1(
        i_data_bus[460]), .B2(n7825), .ZN(n7820) );
  ND2D1BWP30P140LVT U11441 ( .A1(n7821), .A2(n7820), .ZN(N8041) );
  AOI22D1BWP30P140LVT U11442 ( .A1(i_data_bus[426]), .A2(n7824), .B1(
        i_data_bus[394]), .B2(n6214), .ZN(n7823) );
  AOI22D1BWP30P140LVT U11443 ( .A1(i_data_bus[490]), .A2(n7826), .B1(
        i_data_bus[458]), .B2(n7825), .ZN(n7822) );
  ND2D1BWP30P140LVT U11444 ( .A1(n7823), .A2(n7822), .ZN(N8039) );
  AOI22D1BWP30P140LVT U11445 ( .A1(i_data_bus[421]), .A2(n7824), .B1(
        i_data_bus[389]), .B2(n6214), .ZN(n7828) );
  AOI22D1BWP30P140LVT U11446 ( .A1(i_data_bus[485]), .A2(n7826), .B1(
        i_data_bus[453]), .B2(n7825), .ZN(n7827) );
  ND2D1BWP30P140LVT U11447 ( .A1(n7828), .A2(n7827), .ZN(N8034) );
  NR4D1BWP30P140LVT U11448 ( .A1(i_cmd[154]), .A2(n7829), .A3(n10696), .A4(
        n7831), .ZN(n10002) );
  AOI22D1BWP30P140LVT U11449 ( .A1(i_data_bus[569]), .A2(n10002), .B1(
        i_data_bus[537]), .B2(n6222), .ZN(n7835) );
  NR4D1BWP30P140LVT U11450 ( .A1(i_cmd[138]), .A2(n10694), .A3(n7832), .A4(
        n7831), .ZN(n10003) );
  INR4D1BWP30P140LVT U11451 ( .A1(i_cmd[146]), .B1(i_cmd[130]), .B2(n10692), 
        .B3(n7833), .ZN(n10001) );
  AOI22D1BWP30P140LVT U11452 ( .A1(i_data_bus[633]), .A2(n10003), .B1(
        i_data_bus[601]), .B2(n10001), .ZN(n7834) );
  ND2D1BWP30P140LVT U11453 ( .A1(n7835), .A2(n7834), .ZN(N4184) );
  AOI22D1BWP30P140LVT U11454 ( .A1(i_data_bus[560]), .A2(n10002), .B1(
        i_data_bus[528]), .B2(n6222), .ZN(n7837) );
  AOI22D1BWP30P140LVT U11455 ( .A1(i_data_bus[624]), .A2(n10003), .B1(
        i_data_bus[592]), .B2(n10001), .ZN(n7836) );
  ND2D1BWP30P140LVT U11456 ( .A1(n7837), .A2(n7836), .ZN(N4175) );
  AOI22D1BWP30P140LVT U11457 ( .A1(i_data_bus[555]), .A2(n10002), .B1(
        i_data_bus[523]), .B2(n6222), .ZN(n7839) );
  AOI22D1BWP30P140LVT U11458 ( .A1(i_data_bus[619]), .A2(n10003), .B1(
        i_data_bus[587]), .B2(n10001), .ZN(n7838) );
  ND2D1BWP30P140LVT U11459 ( .A1(n7839), .A2(n7838), .ZN(N4170) );
  AOI22D1BWP30P140LVT U11460 ( .A1(i_data_bus[545]), .A2(n10002), .B1(
        i_data_bus[513]), .B2(n6222), .ZN(n7841) );
  AOI22D1BWP30P140LVT U11461 ( .A1(i_data_bus[609]), .A2(n10003), .B1(
        i_data_bus[577]), .B2(n10001), .ZN(n7840) );
  ND2D1BWP30P140LVT U11462 ( .A1(n7841), .A2(n7840), .ZN(N4160) );
  OR2D1BWP30P140LVT U11463 ( .A1(i_cmd[106]), .A2(i_cmd[122]), .Z(n11105) );
  INR4D1BWP30P140LVT U11464 ( .A1(i_cmd[114]), .B1(i_cmd[98]), .B2(n8443), 
        .B3(n11105), .ZN(n8195) );
  INR4D1BWP30P140LVT U11465 ( .A1(i_cmd[122]), .B1(i_cmd[106]), .B2(n7842), 
        .B3(n8447), .ZN(n8194) );
  AOI22D1BWP30P140LVT U11466 ( .A1(n8195), .A2(i_data_bus[473]), .B1(n8194), 
        .B2(i_data_bus[505]), .ZN(n7844) );
  INR4D1BWP30P140LVT U11467 ( .A1(i_cmd[106]), .B1(i_cmd[122]), .B2(n8445), 
        .B3(n7842), .ZN(n8196) );
  NR3D0P7BWP30P140LVT U11468 ( .A1(i_cmd[106]), .A2(i_cmd[122]), .A3(
        i_cmd[114]), .ZN(n11101) );
  AOI22D1BWP30P140LVT U11469 ( .A1(n8196), .A2(i_data_bus[441]), .B1(n6224), 
        .B2(i_data_bus[409]), .ZN(n7843) );
  ND2D1BWP30P140LVT U11470 ( .A1(n7844), .A2(n7843), .ZN(N3968) );
  AOI22D1BWP30P140LVT U11471 ( .A1(n8195), .A2(i_data_bus[468]), .B1(n8194), 
        .B2(i_data_bus[500]), .ZN(n7846) );
  AOI22D1BWP30P140LVT U11472 ( .A1(n8196), .A2(i_data_bus[436]), .B1(n6224), 
        .B2(i_data_bus[404]), .ZN(n7845) );
  ND2D1BWP30P140LVT U11473 ( .A1(n7846), .A2(n7845), .ZN(N3963) );
  AOI22D1BWP30P140LVT U11474 ( .A1(n8195), .A2(i_data_bus[462]), .B1(n8194), 
        .B2(i_data_bus[494]), .ZN(n7848) );
  AOI22D1BWP30P140LVT U11475 ( .A1(n8196), .A2(i_data_bus[430]), .B1(n6224), 
        .B2(i_data_bus[398]), .ZN(n7847) );
  ND2D1BWP30P140LVT U11476 ( .A1(n7848), .A2(n7847), .ZN(N3957) );
  AOI22D1BWP30P140LVT U11477 ( .A1(n8195), .A2(i_data_bus[455]), .B1(n8194), 
        .B2(i_data_bus[487]), .ZN(n7850) );
  AOI22D1BWP30P140LVT U11478 ( .A1(n8196), .A2(i_data_bus[423]), .B1(n6224), 
        .B2(i_data_bus[391]), .ZN(n7849) );
  ND2D1BWP30P140LVT U11479 ( .A1(n7850), .A2(n7849), .ZN(N3950) );
  AOI22D1BWP30P140LVT U11480 ( .A1(n8195), .A2(i_data_bus[454]), .B1(n8194), 
        .B2(i_data_bus[486]), .ZN(n7852) );
  AOI22D1BWP30P140LVT U11481 ( .A1(n8196), .A2(i_data_bus[422]), .B1(n6224), 
        .B2(i_data_bus[390]), .ZN(n7851) );
  ND2D1BWP30P140LVT U11482 ( .A1(n7852), .A2(n7851), .ZN(N3949) );
  AOI22D1BWP30P140LVT U11483 ( .A1(n8196), .A2(i_data_bus[446]), .B1(n8194), 
        .B2(i_data_bus[510]), .ZN(n7854) );
  AOI22D1BWP30P140LVT U11484 ( .A1(n8195), .A2(i_data_bus[478]), .B1(n6224), 
        .B2(i_data_bus[414]), .ZN(n7853) );
  ND2D1BWP30P140LVT U11485 ( .A1(n7854), .A2(n7853), .ZN(N3973) );
  AOI22D1BWP30P140LVT U11486 ( .A1(n8196), .A2(i_data_bus[439]), .B1(n8194), 
        .B2(i_data_bus[503]), .ZN(n7856) );
  AOI22D1BWP30P140LVT U11487 ( .A1(n8195), .A2(i_data_bus[471]), .B1(n6224), 
        .B2(i_data_bus[407]), .ZN(n7855) );
  ND2D1BWP30P140LVT U11488 ( .A1(n7856), .A2(n7855), .ZN(N3966) );
  AOI22D1BWP30P140LVT U11489 ( .A1(n8196), .A2(i_data_bus[435]), .B1(n8194), 
        .B2(i_data_bus[499]), .ZN(n7858) );
  AOI22D1BWP30P140LVT U11490 ( .A1(n8195), .A2(i_data_bus[467]), .B1(n6224), 
        .B2(i_data_bus[403]), .ZN(n7857) );
  ND2D1BWP30P140LVT U11491 ( .A1(n7858), .A2(n7857), .ZN(N3962) );
  AOI22D1BWP30P140LVT U11492 ( .A1(n8196), .A2(i_data_bus[433]), .B1(n8194), 
        .B2(i_data_bus[497]), .ZN(n7860) );
  AOI22D1BWP30P140LVT U11493 ( .A1(n8195), .A2(i_data_bus[465]), .B1(n6224), 
        .B2(i_data_bus[401]), .ZN(n7859) );
  ND2D1BWP30P140LVT U11494 ( .A1(n7860), .A2(n7859), .ZN(N3960) );
  AOI22D1BWP30P140LVT U11495 ( .A1(n8196), .A2(i_data_bus[429]), .B1(n8194), 
        .B2(i_data_bus[493]), .ZN(n7862) );
  AOI22D1BWP30P140LVT U11496 ( .A1(n8195), .A2(i_data_bus[461]), .B1(n6224), 
        .B2(i_data_bus[397]), .ZN(n7861) );
  ND2D1BWP30P140LVT U11497 ( .A1(n7862), .A2(n7861), .ZN(N3956) );
  AOI22D1BWP30P140LVT U11498 ( .A1(n8196), .A2(i_data_bus[427]), .B1(n8194), 
        .B2(i_data_bus[491]), .ZN(n7864) );
  AOI22D1BWP30P140LVT U11499 ( .A1(n8195), .A2(i_data_bus[459]), .B1(n6224), 
        .B2(i_data_bus[395]), .ZN(n7863) );
  ND2D1BWP30P140LVT U11500 ( .A1(n7864), .A2(n7863), .ZN(N3954) );
  AOI22D1BWP30P140LVT U11501 ( .A1(n8196), .A2(i_data_bus[418]), .B1(n8194), 
        .B2(i_data_bus[482]), .ZN(n7866) );
  AOI22D1BWP30P140LVT U11502 ( .A1(n8195), .A2(i_data_bus[450]), .B1(n6224), 
        .B2(i_data_bus[386]), .ZN(n7865) );
  ND2D1BWP30P140LVT U11503 ( .A1(n7866), .A2(n7865), .ZN(N3945) );
  NR4D1BWP30P140LVT U11504 ( .A1(i_cmd[158]), .A2(n10953), .A3(n10696), .A4(
        n7867), .ZN(n10253) );
  NR3D0P7BWP30P140LVT U11505 ( .A1(i_cmd[142]), .A2(i_cmd[158]), .A3(
        i_cmd[150]), .ZN(n10949) );
  AOI22D1BWP30P140LVT U11506 ( .A1(i_data_bus[555]), .A2(n10253), .B1(
        i_data_bus[523]), .B2(n10245), .ZN(n7869) );
  NR4D1BWP30P140LVT U11507 ( .A1(i_cmd[142]), .A2(n10694), .A3(n10952), .A4(
        n7867), .ZN(n10254) );
  INR4D1BWP30P140LVT U11508 ( .A1(i_cmd[150]), .B1(i_cmd[134]), .B2(n10692), 
        .B3(n10950), .ZN(n10252) );
  AOI22D1BWP30P140LVT U11509 ( .A1(i_data_bus[619]), .A2(n10254), .B1(
        i_data_bus[587]), .B2(n10252), .ZN(n7868) );
  ND2D1BWP30P140LVT U11510 ( .A1(n7869), .A2(n7868), .ZN(N9618) );
  INR4D1BWP30P140LVT U11511 ( .A1(i_cmd[139]), .B1(i_cmd[155]), .B2(n10696), 
        .B3(n7870), .ZN(n9935) );
  OR2D1BWP30P140LVT U11512 ( .A1(i_cmd[139]), .A2(i_cmd[155]), .Z(n11074) );
  INR4D1BWP30P140LVT U11513 ( .A1(i_cmd[147]), .B1(i_cmd[131]), .B2(n10692), 
        .B3(n11074), .ZN(n9936) );
  AOI22D1BWP30P140LVT U11514 ( .A1(i_data_bus[573]), .A2(n9935), .B1(
        i_data_bus[605]), .B2(n9936), .ZN(n7872) );
  INR4D1BWP30P140LVT U11515 ( .A1(i_cmd[155]), .B1(i_cmd[139]), .B2(n10694), 
        .B3(n7870), .ZN(n9933) );
  NR3D0P7BWP30P140LVT U11516 ( .A1(i_cmd[139]), .A2(i_cmd[155]), .A3(
        i_cmd[147]), .ZN(n11070) );
  AOI22D1BWP30P140LVT U11517 ( .A1(i_data_bus[637]), .A2(n9933), .B1(
        i_data_bus[541]), .B2(n9934), .ZN(n7871) );
  ND2D1BWP30P140LVT U11518 ( .A1(n7872), .A2(n7871), .ZN(N5422) );
  AOI22D1BWP30P140LVT U11519 ( .A1(i_data_bus[1000]), .A2(n9543), .B1(
        i_data_bus[936]), .B2(n9545), .ZN(n7874) );
  AOI22D1BWP30P140LVT U11520 ( .A1(i_data_bus[968]), .A2(n9544), .B1(
        i_data_bus[904]), .B2(n6226), .ZN(n7873) );
  ND2D1BWP30P140LVT U11521 ( .A1(n7874), .A2(n7873), .ZN(N2091) );
  AOI22D1BWP30P140LVT U11522 ( .A1(i_data_bus[959]), .A2(n9545), .B1(
        i_data_bus[1023]), .B2(n9543), .ZN(n7876) );
  AOI22D1BWP30P140LVT U11523 ( .A1(i_data_bus[991]), .A2(n9544), .B1(
        i_data_bus[927]), .B2(n6226), .ZN(n7875) );
  ND2D1BWP30P140LVT U11524 ( .A1(n7876), .A2(n7875), .ZN(N2114) );
  AOI22D1BWP30P140LVT U11525 ( .A1(i_data_bus[949]), .A2(n9545), .B1(
        i_data_bus[1013]), .B2(n9543), .ZN(n7878) );
  AOI22D1BWP30P140LVT U11526 ( .A1(i_data_bus[981]), .A2(n9544), .B1(
        i_data_bus[917]), .B2(n6226), .ZN(n7877) );
  ND2D1BWP30P140LVT U11527 ( .A1(n7878), .A2(n7877), .ZN(N2104) );
  AOI22D1BWP30P140LVT U11528 ( .A1(i_data_bus[386]), .A2(n6212), .B1(
        i_data_bus[418]), .B2(n8041), .ZN(n7880) );
  AOI22D1BWP30P140LVT U11529 ( .A1(i_data_bus[450]), .A2(n7434), .B1(
        i_data_bus[482]), .B2(n7443), .ZN(n7879) );
  ND2D1BWP30P140LVT U11530 ( .A1(n7880), .A2(n7879), .ZN(N1205) );
  AOI22D1BWP30P140LVT U11531 ( .A1(i_data_bus[479]), .A2(n7434), .B1(
        i_data_bus[447]), .B2(n8041), .ZN(n7882) );
  AOI22D1BWP30P140LVT U11532 ( .A1(i_data_bus[511]), .A2(n7443), .B1(
        i_data_bus[415]), .B2(n6212), .ZN(n7881) );
  ND2D1BWP30P140LVT U11533 ( .A1(n7882), .A2(n7881), .ZN(N1234) );
  AOI22D1BWP30P140LVT U11534 ( .A1(i_data_bus[477]), .A2(n7434), .B1(
        i_data_bus[445]), .B2(n8041), .ZN(n7884) );
  AOI22D1BWP30P140LVT U11535 ( .A1(i_data_bus[413]), .A2(n6212), .B1(
        i_data_bus[509]), .B2(n7443), .ZN(n7883) );
  ND2D1BWP30P140LVT U11536 ( .A1(n7884), .A2(n7883), .ZN(N1232) );
  AOI22D1BWP30P140LVT U11537 ( .A1(i_data_bus[506]), .A2(n7443), .B1(
        i_data_bus[442]), .B2(n8041), .ZN(n7886) );
  AOI22D1BWP30P140LVT U11538 ( .A1(i_data_bus[474]), .A2(n7434), .B1(
        i_data_bus[410]), .B2(n6212), .ZN(n7885) );
  ND2D1BWP30P140LVT U11539 ( .A1(n7886), .A2(n7885), .ZN(N1229) );
  AOI22D1BWP30P140LVT U11540 ( .A1(i_data_bus[409]), .A2(n6212), .B1(
        i_data_bus[441]), .B2(n8041), .ZN(n7888) );
  AOI22D1BWP30P140LVT U11541 ( .A1(i_data_bus[505]), .A2(n7443), .B1(
        i_data_bus[473]), .B2(n7434), .ZN(n7887) );
  ND2D1BWP30P140LVT U11542 ( .A1(n7888), .A2(n7887), .ZN(N1228) );
  AOI22D1BWP30P140LVT U11543 ( .A1(i_data_bus[400]), .A2(n6212), .B1(
        i_data_bus[432]), .B2(n8041), .ZN(n7890) );
  AOI22D1BWP30P140LVT U11544 ( .A1(i_data_bus[496]), .A2(n7443), .B1(
        i_data_bus[464]), .B2(n7434), .ZN(n7889) );
  ND2D1BWP30P140LVT U11545 ( .A1(n7890), .A2(n7889), .ZN(N1219) );
  AOI22D1BWP30P140LVT U11546 ( .A1(i_data_bus[463]), .A2(n7434), .B1(
        i_data_bus[431]), .B2(n8041), .ZN(n7892) );
  AOI22D1BWP30P140LVT U11547 ( .A1(i_data_bus[495]), .A2(n7443), .B1(
        i_data_bus[399]), .B2(n6212), .ZN(n7891) );
  ND2D1BWP30P140LVT U11548 ( .A1(n7892), .A2(n7891), .ZN(N1218) );
  AOI22D1BWP30P140LVT U11549 ( .A1(i_data_bus[488]), .A2(n7443), .B1(
        i_data_bus[424]), .B2(n8041), .ZN(n7894) );
  AOI22D1BWP30P140LVT U11550 ( .A1(i_data_bus[456]), .A2(n7434), .B1(
        i_data_bus[392]), .B2(n6212), .ZN(n7893) );
  ND2D1BWP30P140LVT U11551 ( .A1(n7894), .A2(n7893), .ZN(N1211) );
  AOI22D1BWP30P140LVT U11552 ( .A1(i_data_bus[509]), .A2(n7909), .B1(
        i_data_bus[477]), .B2(n7911), .ZN(n7896) );
  AOI22D1BWP30P140LVT U11553 ( .A1(i_data_bus[413]), .A2(n6215), .B1(
        i_data_bus[445]), .B2(n7910), .ZN(n7895) );
  ND2D1BWP30P140LVT U11554 ( .A1(n7896), .A2(n7895), .ZN(N5334) );
  AOI22D1BWP30P140LVT U11555 ( .A1(i_data_bus[474]), .A2(n7911), .B1(
        i_data_bus[410]), .B2(n6215), .ZN(n7898) );
  AOI22D1BWP30P140LVT U11556 ( .A1(i_data_bus[506]), .A2(n7909), .B1(
        i_data_bus[442]), .B2(n7910), .ZN(n7897) );
  ND2D1BWP30P140LVT U11557 ( .A1(n7898), .A2(n7897), .ZN(N5331) );
  AOI22D1BWP30P140LVT U11558 ( .A1(i_data_bus[406]), .A2(n6215), .B1(
        i_data_bus[470]), .B2(n7911), .ZN(n7900) );
  AOI22D1BWP30P140LVT U11559 ( .A1(i_data_bus[502]), .A2(n7909), .B1(
        i_data_bus[438]), .B2(n7910), .ZN(n7899) );
  ND2D1BWP30P140LVT U11560 ( .A1(n7900), .A2(n7899), .ZN(N5327) );
  AOI22D1BWP30P140LVT U11561 ( .A1(i_data_bus[469]), .A2(n7911), .B1(
        i_data_bus[405]), .B2(n6215), .ZN(n7902) );
  AOI22D1BWP30P140LVT U11562 ( .A1(i_data_bus[501]), .A2(n7909), .B1(
        i_data_bus[437]), .B2(n7910), .ZN(n7901) );
  ND2D1BWP30P140LVT U11563 ( .A1(n7902), .A2(n7901), .ZN(N5326) );
  AOI22D1BWP30P140LVT U11564 ( .A1(i_data_bus[403]), .A2(n6215), .B1(
        i_data_bus[499]), .B2(n7909), .ZN(n7904) );
  AOI22D1BWP30P140LVT U11565 ( .A1(i_data_bus[467]), .A2(n7911), .B1(
        i_data_bus[435]), .B2(n7910), .ZN(n7903) );
  ND2D1BWP30P140LVT U11566 ( .A1(n7904), .A2(n7903), .ZN(N5324) );
  AOI22D1BWP30P140LVT U11567 ( .A1(i_data_bus[401]), .A2(n6215), .B1(
        i_data_bus[497]), .B2(n7909), .ZN(n7906) );
  AOI22D1BWP30P140LVT U11568 ( .A1(i_data_bus[465]), .A2(n7911), .B1(
        i_data_bus[433]), .B2(n7910), .ZN(n7905) );
  ND2D1BWP30P140LVT U11569 ( .A1(n7906), .A2(n7905), .ZN(N5322) );
  AOI22D1BWP30P140LVT U11570 ( .A1(i_data_bus[397]), .A2(n6215), .B1(
        i_data_bus[493]), .B2(n7909), .ZN(n7908) );
  AOI22D1BWP30P140LVT U11571 ( .A1(i_data_bus[461]), .A2(n7911), .B1(
        i_data_bus[429]), .B2(n7910), .ZN(n7907) );
  ND2D1BWP30P140LVT U11572 ( .A1(n7908), .A2(n7907), .ZN(N5318) );
  AOI22D1BWP30P140LVT U11573 ( .A1(i_data_bus[481]), .A2(n7909), .B1(
        i_data_bus[385]), .B2(n6215), .ZN(n7913) );
  AOI22D1BWP30P140LVT U11574 ( .A1(i_data_bus[449]), .A2(n7911), .B1(
        i_data_bus[417]), .B2(n7910), .ZN(n7912) );
  ND2D1BWP30P140LVT U11575 ( .A1(n7913), .A2(n7912), .ZN(N5306) );
  NR4D1BWP30P140LVT U11576 ( .A1(i_cmd[156]), .A2(n7914), .A3(n10696), .A4(
        n11030), .ZN(n10184) );
  INR4D1BWP30P140LVT U11577 ( .A1(i_cmd[148]), .B1(i_cmd[132]), .B2(n10692), 
        .B3(n11027), .ZN(n10183) );
  AOI22D1BWP30P140LVT U11578 ( .A1(i_data_bus[573]), .A2(n10184), .B1(
        i_data_bus[605]), .B2(n10183), .ZN(n7916) );
  NR4D1BWP30P140LVT U11579 ( .A1(i_cmd[140]), .A2(n7914), .A3(n10694), .A4(
        n11029), .ZN(n10185) );
  NR3D0P7BWP30P140LVT U11580 ( .A1(i_cmd[148]), .A2(i_cmd[140]), .A3(
        i_cmd[156]), .ZN(n11026) );
  AOI22D1BWP30P140LVT U11581 ( .A1(i_data_bus[637]), .A2(n10185), .B1(
        i_data_bus[541]), .B2(n10182), .ZN(n7915) );
  ND2D1BWP30P140LVT U11582 ( .A1(n7916), .A2(n7915), .ZN(N6912) );
  AOI22D1BWP30P140LVT U11583 ( .A1(i_data_bus[560]), .A2(n10184), .B1(
        i_data_bus[592]), .B2(n10183), .ZN(n7918) );
  AOI22D1BWP30P140LVT U11584 ( .A1(i_data_bus[624]), .A2(n10185), .B1(
        i_data_bus[528]), .B2(n10182), .ZN(n7917) );
  ND2D1BWP30P140LVT U11585 ( .A1(n7918), .A2(n7917), .ZN(N6899) );
  AOI22D1BWP30P140LVT U11586 ( .A1(i_data_bus[915]), .A2(n6226), .B1(
        i_data_bus[1011]), .B2(n9543), .ZN(n7920) );
  AOI22D1BWP30P140LVT U11587 ( .A1(i_data_bus[979]), .A2(n9544), .B1(
        i_data_bus[947]), .B2(n9545), .ZN(n7919) );
  ND2D1BWP30P140LVT U11588 ( .A1(n7920), .A2(n7919), .ZN(N2102) );
  AOI22D1BWP30P140LVT U11589 ( .A1(i_data_bus[934]), .A2(n9545), .B1(
        i_data_bus[902]), .B2(n6226), .ZN(n7922) );
  AOI22D1BWP30P140LVT U11590 ( .A1(i_data_bus[966]), .A2(n9544), .B1(
        i_data_bus[998]), .B2(n9543), .ZN(n7921) );
  ND2D1BWP30P140LVT U11591 ( .A1(n7922), .A2(n7921), .ZN(N2089) );
  AOI22D1BWP30P140LVT U11592 ( .A1(i_data_bus[923]), .A2(n6226), .B1(
        i_data_bus[955]), .B2(n9545), .ZN(n7924) );
  AOI22D1BWP30P140LVT U11593 ( .A1(i_data_bus[987]), .A2(n9544), .B1(
        i_data_bus[1019]), .B2(n9543), .ZN(n7923) );
  ND2D1BWP30P140LVT U11594 ( .A1(n7924), .A2(n7923), .ZN(N2110) );
  AOI22D1BWP30P140LVT U11595 ( .A1(i_data_bus[939]), .A2(n9545), .B1(
        i_data_bus[907]), .B2(n6226), .ZN(n7926) );
  AOI22D1BWP30P140LVT U11596 ( .A1(i_data_bus[971]), .A2(n9544), .B1(
        i_data_bus[1003]), .B2(n9543), .ZN(n7925) );
  ND2D1BWP30P140LVT U11597 ( .A1(n7926), .A2(n7925), .ZN(N2094) );
  AOI22D1BWP30P140LVT U11598 ( .A1(i_data_bus[555]), .A2(n9935), .B1(
        i_data_bus[523]), .B2(n9934), .ZN(n7928) );
  AOI22D1BWP30P140LVT U11599 ( .A1(i_data_bus[619]), .A2(n9933), .B1(
        i_data_bus[587]), .B2(n9936), .ZN(n7927) );
  ND2D1BWP30P140LVT U11600 ( .A1(n7928), .A2(n7927), .ZN(N5404) );
  AOI22D1BWP30P140LVT U11601 ( .A1(i_data_bus[567]), .A2(n10184), .B1(
        i_data_bus[535]), .B2(n10182), .ZN(n7930) );
  AOI22D1BWP30P140LVT U11602 ( .A1(i_data_bus[631]), .A2(n10185), .B1(
        i_data_bus[599]), .B2(n10183), .ZN(n7929) );
  ND2D1BWP30P140LVT U11603 ( .A1(n7930), .A2(n7929), .ZN(N6906) );
  AOI22D1BWP30P140LVT U11604 ( .A1(i_data_bus[545]), .A2(n10184), .B1(
        i_data_bus[513]), .B2(n10182), .ZN(n7932) );
  AOI22D1BWP30P140LVT U11605 ( .A1(i_data_bus[609]), .A2(n10185), .B1(
        i_data_bus[577]), .B2(n10183), .ZN(n7931) );
  ND2D1BWP30P140LVT U11606 ( .A1(n7932), .A2(n7931), .ZN(N6884) );
  AOI22D1BWP30P140LVT U11607 ( .A1(i_data_bus[935]), .A2(n9660), .B1(
        i_data_bus[999]), .B2(n9663), .ZN(n7934) );
  AOI22D1BWP30P140LVT U11608 ( .A1(i_data_bus[967]), .A2(n9662), .B1(
        i_data_bus[903]), .B2(n9661), .ZN(n7933) );
  ND2D1BWP30P140LVT U11609 ( .A1(n7934), .A2(n7933), .ZN(N7538) );
  AOI22D1BWP30P140LVT U11610 ( .A1(i_data_bus[449]), .A2(n8124), .B1(
        i_data_bus[481]), .B2(n8123), .ZN(n7940) );
  AOI22D1BWP30P140LVT U11611 ( .A1(i_data_bus[417]), .A2(n8125), .B1(
        i_data_bus[385]), .B2(n8122), .ZN(n7939) );
  ND2D1BWP30P140LVT U11612 ( .A1(n7940), .A2(n7939), .ZN(N2582) );
  AOI22D1BWP30P140LVT U11613 ( .A1(i_data_bus[993]), .A2(n9663), .B1(
        i_data_bus[897]), .B2(n9661), .ZN(n7942) );
  AOI22D1BWP30P140LVT U11614 ( .A1(i_data_bus[961]), .A2(n9662), .B1(
        i_data_bus[929]), .B2(n9660), .ZN(n7941) );
  ND2D1BWP30P140LVT U11615 ( .A1(n7942), .A2(n7941), .ZN(N7532) );
  AOI22D1BWP30P140LVT U11616 ( .A1(i_data_bus[956]), .A2(n9660), .B1(
        i_data_bus[924]), .B2(n9661), .ZN(n7944) );
  AOI22D1BWP30P140LVT U11617 ( .A1(i_data_bus[988]), .A2(n9662), .B1(
        i_data_bus[1020]), .B2(n9663), .ZN(n7943) );
  ND2D1BWP30P140LVT U11618 ( .A1(n7944), .A2(n7943), .ZN(N7559) );
  AOI22D1BWP30P140LVT U11619 ( .A1(i_data_bus[920]), .A2(n9661), .B1(
        i_data_bus[952]), .B2(n9660), .ZN(n7946) );
  AOI22D1BWP30P140LVT U11620 ( .A1(i_data_bus[984]), .A2(n9662), .B1(
        i_data_bus[1016]), .B2(n9663), .ZN(n7945) );
  ND2D1BWP30P140LVT U11621 ( .A1(n7946), .A2(n7945), .ZN(N7555) );
  AOI22D1BWP30P140LVT U11622 ( .A1(i_data_bus[915]), .A2(n9661), .B1(
        i_data_bus[947]), .B2(n9660), .ZN(n7948) );
  AOI22D1BWP30P140LVT U11623 ( .A1(i_data_bus[979]), .A2(n9662), .B1(
        i_data_bus[1011]), .B2(n9663), .ZN(n7947) );
  ND2D1BWP30P140LVT U11624 ( .A1(n7948), .A2(n7947), .ZN(N7550) );
  AOI22D1BWP30P140LVT U11625 ( .A1(i_data_bus[913]), .A2(n9661), .B1(
        i_data_bus[945]), .B2(n9660), .ZN(n7950) );
  AOI22D1BWP30P140LVT U11626 ( .A1(i_data_bus[977]), .A2(n9662), .B1(
        i_data_bus[1009]), .B2(n9663), .ZN(n7949) );
  ND2D1BWP30P140LVT U11627 ( .A1(n7950), .A2(n7949), .ZN(N7548) );
  AOI22D1BWP30P140LVT U11628 ( .A1(i_data_bus[904]), .A2(n9661), .B1(
        i_data_bus[936]), .B2(n9660), .ZN(n7952) );
  AOI22D1BWP30P140LVT U11629 ( .A1(i_data_bus[968]), .A2(n9662), .B1(
        i_data_bus[1000]), .B2(n9663), .ZN(n7951) );
  ND2D1BWP30P140LVT U11630 ( .A1(n7952), .A2(n7951), .ZN(N7539) );
  AOI22D1BWP30P140LVT U11631 ( .A1(i_data_bus[506]), .A2(n8123), .B1(
        i_data_bus[442]), .B2(n8125), .ZN(n7954) );
  AOI22D1BWP30P140LVT U11632 ( .A1(i_data_bus[474]), .A2(n8124), .B1(
        i_data_bus[410]), .B2(n8122), .ZN(n7953) );
  ND2D1BWP30P140LVT U11633 ( .A1(n7954), .A2(n7953), .ZN(N2607) );
  AOI22D1BWP30P140LVT U11634 ( .A1(i_data_bus[475]), .A2(n8124), .B1(
        i_data_bus[443]), .B2(n8125), .ZN(n7956) );
  AOI22D1BWP30P140LVT U11635 ( .A1(i_data_bus[507]), .A2(n8123), .B1(
        i_data_bus[411]), .B2(n8122), .ZN(n7955) );
  ND2D1BWP30P140LVT U11636 ( .A1(n7956), .A2(n7955), .ZN(N2608) );
  AOI22D1BWP30P140LVT U11637 ( .A1(i_data_bus[560]), .A2(n10253), .B1(
        i_data_bus[528]), .B2(n10245), .ZN(n7958) );
  AOI22D1BWP30P140LVT U11638 ( .A1(i_data_bus[624]), .A2(n10254), .B1(
        i_data_bus[592]), .B2(n10252), .ZN(n7957) );
  ND2D1BWP30P140LVT U11639 ( .A1(n7958), .A2(n7957), .ZN(N9623) );
  AOI22D1BWP30P140LVT U11640 ( .A1(i_data_bus[498]), .A2(n8123), .B1(
        i_data_bus[466]), .B2(n8124), .ZN(n7960) );
  AOI22D1BWP30P140LVT U11641 ( .A1(i_data_bus[434]), .A2(n8125), .B1(
        i_data_bus[402]), .B2(n8122), .ZN(n7959) );
  ND2D1BWP30P140LVT U11642 ( .A1(n7960), .A2(n7959), .ZN(N2599) );
  INR4D1BWP30P140LVT U11643 ( .A1(i_cmd[141]), .B1(i_cmd[157]), .B2(n10696), 
        .B3(n7961), .ZN(n10271) );
  NR3D0P7BWP30P140LVT U11644 ( .A1(i_cmd[141]), .A2(i_cmd[157]), .A3(
        i_cmd[149]), .ZN(n10985) );
  AOI22D1BWP30P140LVT U11645 ( .A1(i_data_bus[560]), .A2(n10271), .B1(
        i_data_bus[528]), .B2(n10272), .ZN(n7963) );
  INR4D1BWP30P140LVT U11646 ( .A1(i_cmd[157]), .B1(i_cmd[141]), .B2(n10694), 
        .B3(n7961), .ZN(n10270) );
  OR2D1BWP30P140LVT U11647 ( .A1(i_cmd[141]), .A2(i_cmd[157]), .Z(n10989) );
  INR4D1BWP30P140LVT U11648 ( .A1(i_cmd[149]), .B1(i_cmd[133]), .B2(n10692), 
        .B3(n10989), .ZN(n10269) );
  AOI22D1BWP30P140LVT U11649 ( .A1(i_data_bus[624]), .A2(n10270), .B1(
        i_data_bus[592]), .B2(n10269), .ZN(n7962) );
  ND2D1BWP30P140LVT U11650 ( .A1(n7963), .A2(n7962), .ZN(N8133) );
  AOI22D1BWP30P140LVT U11651 ( .A1(i_data_bus[559]), .A2(n10271), .B1(
        i_data_bus[527]), .B2(n10272), .ZN(n7965) );
  AOI22D1BWP30P140LVT U11652 ( .A1(i_data_bus[623]), .A2(n10270), .B1(
        i_data_bus[591]), .B2(n10269), .ZN(n7964) );
  ND2D1BWP30P140LVT U11653 ( .A1(n7965), .A2(n7964), .ZN(N8132) );
  AOI22D1BWP30P140LVT U11654 ( .A1(i_data_bus[633]), .A2(n9933), .B1(
        i_data_bus[601]), .B2(n9936), .ZN(n7967) );
  AOI22D1BWP30P140LVT U11655 ( .A1(i_data_bus[569]), .A2(n9935), .B1(
        i_data_bus[537]), .B2(n9934), .ZN(n7966) );
  ND2D1BWP30P140LVT U11656 ( .A1(n7967), .A2(n7966), .ZN(N5418) );
  AOI22D1BWP30P140LVT U11657 ( .A1(i_data_bus[631]), .A2(n10003), .B1(
        i_data_bus[599]), .B2(n10001), .ZN(n7969) );
  AOI22D1BWP30P140LVT U11658 ( .A1(i_data_bus[567]), .A2(n10002), .B1(
        i_data_bus[535]), .B2(n6222), .ZN(n7968) );
  ND2D1BWP30P140LVT U11659 ( .A1(n7969), .A2(n7968), .ZN(N4182) );
  AOI22D1BWP30P140LVT U11660 ( .A1(i_data_bus[624]), .A2(n9933), .B1(
        i_data_bus[528]), .B2(n9934), .ZN(n7971) );
  AOI22D1BWP30P140LVT U11661 ( .A1(i_data_bus[560]), .A2(n9935), .B1(
        i_data_bus[592]), .B2(n9936), .ZN(n7970) );
  ND2D1BWP30P140LVT U11662 ( .A1(n7971), .A2(n7970), .ZN(N5409) );
  AOI22D1BWP30P140LVT U11663 ( .A1(i_data_bus[615]), .A2(n9933), .B1(
        i_data_bus[519]), .B2(n9934), .ZN(n7973) );
  AOI22D1BWP30P140LVT U11664 ( .A1(i_data_bus[551]), .A2(n9935), .B1(
        i_data_bus[583]), .B2(n9936), .ZN(n7972) );
  ND2D1BWP30P140LVT U11665 ( .A1(n7973), .A2(n7972), .ZN(N5400) );
  AOI22D1BWP30P140LVT U11666 ( .A1(i_data_bus[609]), .A2(n9933), .B1(
        i_data_bus[513]), .B2(n9934), .ZN(n7975) );
  AOI22D1BWP30P140LVT U11667 ( .A1(i_data_bus[545]), .A2(n9935), .B1(
        i_data_bus[577]), .B2(n9936), .ZN(n7974) );
  ND2D1BWP30P140LVT U11668 ( .A1(n7975), .A2(n7974), .ZN(N5394) );
  AOI22D1BWP30P140LVT U11669 ( .A1(i_data_bus[615]), .A2(n10003), .B1(
        i_data_bus[519]), .B2(n6222), .ZN(n7977) );
  AOI22D1BWP30P140LVT U11670 ( .A1(i_data_bus[551]), .A2(n10002), .B1(
        i_data_bus[583]), .B2(n10001), .ZN(n7976) );
  ND2D1BWP30P140LVT U11671 ( .A1(n7977), .A2(n7976), .ZN(N4166) );
  NR4D1BWP30P140LVT U11672 ( .A1(i_cmd[137]), .A2(n10694), .A3(n11128), .A4(
        n7978), .ZN(n10011) );
  NR3D0P7BWP30P140LVT U11673 ( .A1(i_cmd[137]), .A2(i_cmd[153]), .A3(
        i_cmd[145]), .ZN(n11125) );
  AOI22D1BWP30P140LVT U11674 ( .A1(i_data_bus[615]), .A2(n10011), .B1(
        i_data_bus[519]), .B2(n10006), .ZN(n7980) );
  NR4D1BWP30P140LVT U11675 ( .A1(i_cmd[153]), .A2(n11129), .A3(n10696), .A4(
        n7978), .ZN(n10012) );
  INR4D1BWP30P140LVT U11676 ( .A1(i_cmd[145]), .B1(i_cmd[129]), .B2(n10692), 
        .B3(n11126), .ZN(n10013) );
  AOI22D1BWP30P140LVT U11677 ( .A1(i_data_bus[551]), .A2(n10012), .B1(
        i_data_bus[583]), .B2(n10013), .ZN(n7979) );
  ND2D1BWP30P140LVT U11678 ( .A1(n7980), .A2(n7979), .ZN(N2676) );
  AOI22D1BWP30P140LVT U11679 ( .A1(i_data_bus[609]), .A2(n10011), .B1(
        i_data_bus[513]), .B2(n10006), .ZN(n7982) );
  AOI22D1BWP30P140LVT U11680 ( .A1(i_data_bus[545]), .A2(n10012), .B1(
        i_data_bus[577]), .B2(n10013), .ZN(n7981) );
  ND2D1BWP30P140LVT U11681 ( .A1(n7982), .A2(n7981), .ZN(N2670) );
  AOI22D1BWP30P140LVT U11682 ( .A1(i_data_bus[623]), .A2(n10185), .B1(
        i_data_bus[591]), .B2(n10183), .ZN(n7984) );
  AOI22D1BWP30P140LVT U11683 ( .A1(i_data_bus[559]), .A2(n10184), .B1(
        i_data_bus[527]), .B2(n10182), .ZN(n7983) );
  ND2D1BWP30P140LVT U11684 ( .A1(n7984), .A2(n7983), .ZN(N6898) );
  AOI22D1BWP30P140LVT U11685 ( .A1(n8196), .A2(i_data_bus[447]), .B1(n6224), 
        .B2(i_data_bus[415]), .ZN(n7986) );
  AOI22D1BWP30P140LVT U11686 ( .A1(n8195), .A2(i_data_bus[479]), .B1(n8194), 
        .B2(i_data_bus[511]), .ZN(n7985) );
  ND2D1BWP30P140LVT U11687 ( .A1(n7986), .A2(n7985), .ZN(N3974) );
  AOI22D1BWP30P140LVT U11688 ( .A1(n8195), .A2(i_data_bus[476]), .B1(n6224), 
        .B2(i_data_bus[412]), .ZN(n7988) );
  AOI22D1BWP30P140LVT U11689 ( .A1(n8196), .A2(i_data_bus[444]), .B1(n8194), 
        .B2(i_data_bus[508]), .ZN(n7987) );
  ND2D1BWP30P140LVT U11690 ( .A1(n7988), .A2(n7987), .ZN(N3971) );
  AOI22D1BWP30P140LVT U11691 ( .A1(n8196), .A2(i_data_bus[443]), .B1(n6224), 
        .B2(i_data_bus[411]), .ZN(n7990) );
  AOI22D1BWP30P140LVT U11692 ( .A1(n8195), .A2(i_data_bus[475]), .B1(n8194), 
        .B2(i_data_bus[507]), .ZN(n7989) );
  ND2D1BWP30P140LVT U11693 ( .A1(n7990), .A2(n7989), .ZN(N3970) );
  AOI22D1BWP30P140LVT U11694 ( .A1(n8196), .A2(i_data_bus[442]), .B1(n6224), 
        .B2(i_data_bus[410]), .ZN(n7992) );
  AOI22D1BWP30P140LVT U11695 ( .A1(n8195), .A2(i_data_bus[474]), .B1(n8194), 
        .B2(i_data_bus[506]), .ZN(n7991) );
  ND2D1BWP30P140LVT U11696 ( .A1(n7992), .A2(n7991), .ZN(N3969) );
  AOI22D1BWP30P140LVT U11697 ( .A1(n8195), .A2(i_data_bus[472]), .B1(n6224), 
        .B2(i_data_bus[408]), .ZN(n7994) );
  AOI22D1BWP30P140LVT U11698 ( .A1(n8196), .A2(i_data_bus[440]), .B1(n8194), 
        .B2(i_data_bus[504]), .ZN(n7993) );
  ND2D1BWP30P140LVT U11699 ( .A1(n7994), .A2(n7993), .ZN(N3967) );
  AOI22D1BWP30P140LVT U11700 ( .A1(n8195), .A2(i_data_bus[470]), .B1(n6224), 
        .B2(i_data_bus[406]), .ZN(n7996) );
  AOI22D1BWP30P140LVT U11701 ( .A1(n8196), .A2(i_data_bus[438]), .B1(n8194), 
        .B2(i_data_bus[502]), .ZN(n7995) );
  ND2D1BWP30P140LVT U11702 ( .A1(n7996), .A2(n7995), .ZN(N3965) );
  AOI22D1BWP30P140LVT U11703 ( .A1(n8196), .A2(i_data_bus[437]), .B1(n6224), 
        .B2(i_data_bus[405]), .ZN(n7998) );
  AOI22D1BWP30P140LVT U11704 ( .A1(n8195), .A2(i_data_bus[469]), .B1(n8194), 
        .B2(i_data_bus[501]), .ZN(n7997) );
  ND2D1BWP30P140LVT U11705 ( .A1(n7998), .A2(n7997), .ZN(N3964) );
  AOI22D1BWP30P140LVT U11706 ( .A1(n8195), .A2(i_data_bus[466]), .B1(n6224), 
        .B2(i_data_bus[402]), .ZN(n8000) );
  AOI22D1BWP30P140LVT U11707 ( .A1(n8196), .A2(i_data_bus[434]), .B1(n8194), 
        .B2(i_data_bus[498]), .ZN(n7999) );
  ND2D1BWP30P140LVT U11708 ( .A1(n8000), .A2(n7999), .ZN(N3961) );
  AOI22D1BWP30P140LVT U11709 ( .A1(n8196), .A2(i_data_bus[431]), .B1(n6224), 
        .B2(i_data_bus[399]), .ZN(n8002) );
  AOI22D1BWP30P140LVT U11710 ( .A1(n8195), .A2(i_data_bus[463]), .B1(n8194), 
        .B2(i_data_bus[495]), .ZN(n8001) );
  ND2D1BWP30P140LVT U11711 ( .A1(n8002), .A2(n8001), .ZN(N3958) );
  AOI22D1BWP30P140LVT U11712 ( .A1(n8195), .A2(i_data_bus[460]), .B1(n6224), 
        .B2(i_data_bus[396]), .ZN(n8004) );
  AOI22D1BWP30P140LVT U11713 ( .A1(n8196), .A2(i_data_bus[428]), .B1(n8194), 
        .B2(i_data_bus[492]), .ZN(n8003) );
  ND2D1BWP30P140LVT U11714 ( .A1(n8004), .A2(n8003), .ZN(N3955) );
  AOI22D1BWP30P140LVT U11715 ( .A1(n8195), .A2(i_data_bus[458]), .B1(n6224), 
        .B2(i_data_bus[394]), .ZN(n8006) );
  AOI22D1BWP30P140LVT U11716 ( .A1(n8196), .A2(i_data_bus[426]), .B1(n8194), 
        .B2(i_data_bus[490]), .ZN(n8005) );
  ND2D1BWP30P140LVT U11717 ( .A1(n8006), .A2(n8005), .ZN(N3953) );
  AOI22D1BWP30P140LVT U11718 ( .A1(n8196), .A2(i_data_bus[424]), .B1(n6224), 
        .B2(i_data_bus[392]), .ZN(n8008) );
  AOI22D1BWP30P140LVT U11719 ( .A1(n8195), .A2(i_data_bus[456]), .B1(n8194), 
        .B2(i_data_bus[488]), .ZN(n8007) );
  ND2D1BWP30P140LVT U11720 ( .A1(n8008), .A2(n8007), .ZN(N3951) );
  AOI22D1BWP30P140LVT U11721 ( .A1(n8195), .A2(i_data_bus[453]), .B1(n6224), 
        .B2(i_data_bus[389]), .ZN(n8010) );
  AOI22D1BWP30P140LVT U11722 ( .A1(n8196), .A2(i_data_bus[421]), .B1(n8194), 
        .B2(i_data_bus[485]), .ZN(n8009) );
  ND2D1BWP30P140LVT U11723 ( .A1(n8010), .A2(n8009), .ZN(N3948) );
  AOI22D1BWP30P140LVT U11724 ( .A1(n8196), .A2(i_data_bus[445]), .B1(n8195), 
        .B2(i_data_bus[477]), .ZN(n8012) );
  AOI22D1BWP30P140LVT U11725 ( .A1(n8194), .A2(i_data_bus[509]), .B1(n6224), 
        .B2(i_data_bus[413]), .ZN(n8011) );
  ND2D1BWP30P140LVT U11726 ( .A1(n8012), .A2(n8011), .ZN(N3972) );
  AOI22D1BWP30P140LVT U11727 ( .A1(n8196), .A2(i_data_bus[432]), .B1(n8195), 
        .B2(i_data_bus[464]), .ZN(n8014) );
  AOI22D1BWP30P140LVT U11728 ( .A1(n8194), .A2(i_data_bus[496]), .B1(n6224), 
        .B2(i_data_bus[400]), .ZN(n8013) );
  ND2D1BWP30P140LVT U11729 ( .A1(n8014), .A2(n8013), .ZN(N3959) );
  AOI22D1BWP30P140LVT U11730 ( .A1(i_data_bus[633]), .A2(n10011), .B1(
        i_data_bus[601]), .B2(n10013), .ZN(n8016) );
  AOI22D1BWP30P140LVT U11731 ( .A1(i_data_bus[569]), .A2(n10012), .B1(
        i_data_bus[537]), .B2(n10006), .ZN(n8015) );
  ND2D1BWP30P140LVT U11732 ( .A1(n8016), .A2(n8015), .ZN(N2694) );
  AOI22D1BWP30P140LVT U11733 ( .A1(i_data_bus[631]), .A2(n10270), .B1(
        i_data_bus[535]), .B2(n10272), .ZN(n8018) );
  AOI22D1BWP30P140LVT U11734 ( .A1(i_data_bus[567]), .A2(n10271), .B1(
        i_data_bus[599]), .B2(n10269), .ZN(n8017) );
  ND2D1BWP30P140LVT U11735 ( .A1(n8018), .A2(n8017), .ZN(N8140) );
  AOI22D1BWP30P140LVT U11736 ( .A1(i_data_bus[620]), .A2(n10270), .B1(
        i_data_bus[524]), .B2(n10272), .ZN(n8020) );
  AOI22D1BWP30P140LVT U11737 ( .A1(i_data_bus[556]), .A2(n10271), .B1(
        i_data_bus[588]), .B2(n10269), .ZN(n8019) );
  ND2D1BWP30P140LVT U11738 ( .A1(n8020), .A2(n8019), .ZN(N8129) );
  AOI22D1BWP30P140LVT U11739 ( .A1(i_data_bus[615]), .A2(n10270), .B1(
        i_data_bus[519]), .B2(n10272), .ZN(n8022) );
  AOI22D1BWP30P140LVT U11740 ( .A1(i_data_bus[551]), .A2(n10271), .B1(
        i_data_bus[583]), .B2(n10269), .ZN(n8021) );
  ND2D1BWP30P140LVT U11741 ( .A1(n8022), .A2(n8021), .ZN(N8124) );
  AOI22D1BWP30P140LVT U11742 ( .A1(i_data_bus[560]), .A2(n10012), .B1(
        i_data_bus[592]), .B2(n10013), .ZN(n8024) );
  AOI22D1BWP30P140LVT U11743 ( .A1(i_data_bus[624]), .A2(n10011), .B1(
        i_data_bus[528]), .B2(n10006), .ZN(n8023) );
  ND2D1BWP30P140LVT U11744 ( .A1(n8024), .A2(n8023), .ZN(N2685) );
  AOI22D1BWP30P140LVT U11745 ( .A1(i_data_bus[556]), .A2(n10012), .B1(
        i_data_bus[588]), .B2(n10013), .ZN(n8026) );
  AOI22D1BWP30P140LVT U11746 ( .A1(i_data_bus[620]), .A2(n10011), .B1(
        i_data_bus[524]), .B2(n10006), .ZN(n8025) );
  ND2D1BWP30P140LVT U11747 ( .A1(n8026), .A2(n8025), .ZN(N2681) );
  AOI22D1BWP30P140LVT U11748 ( .A1(i_data_bus[637]), .A2(n10254), .B1(
        i_data_bus[541]), .B2(n10245), .ZN(n8028) );
  AOI22D1BWP30P140LVT U11749 ( .A1(i_data_bus[573]), .A2(n10253), .B1(
        i_data_bus[605]), .B2(n10252), .ZN(n8027) );
  ND2D1BWP30P140LVT U11750 ( .A1(n8028), .A2(n8027), .ZN(N9636) );
  AOI22D1BWP30P140LVT U11751 ( .A1(i_data_bus[623]), .A2(n10254), .B1(
        i_data_bus[527]), .B2(n10245), .ZN(n8030) );
  AOI22D1BWP30P140LVT U11752 ( .A1(i_data_bus[559]), .A2(n10253), .B1(
        i_data_bus[591]), .B2(n10252), .ZN(n8029) );
  ND2D1BWP30P140LVT U11753 ( .A1(n8030), .A2(n8029), .ZN(N9622) );
  AOI22D1BWP30P140LVT U11754 ( .A1(i_data_bus[609]), .A2(n10254), .B1(
        i_data_bus[513]), .B2(n10245), .ZN(n8032) );
  AOI22D1BWP30P140LVT U11755 ( .A1(i_data_bus[545]), .A2(n10253), .B1(
        i_data_bus[577]), .B2(n10252), .ZN(n8031) );
  ND2D1BWP30P140LVT U11756 ( .A1(n8032), .A2(n8031), .ZN(N9608) );
  AOI22D1BWP30P140LVT U11757 ( .A1(i_data_bus[475]), .A2(n7434), .B1(
        i_data_bus[411]), .B2(n6212), .ZN(n8034) );
  AOI22D1BWP30P140LVT U11758 ( .A1(i_data_bus[507]), .A2(n7443), .B1(
        i_data_bus[443]), .B2(n8041), .ZN(n8033) );
  ND2D1BWP30P140LVT U11759 ( .A1(n8034), .A2(n8033), .ZN(N1230) );
  AOI22D1BWP30P140LVT U11760 ( .A1(i_data_bus[500]), .A2(n7443), .B1(
        i_data_bus[468]), .B2(n7434), .ZN(n8036) );
  AOI22D1BWP30P140LVT U11761 ( .A1(i_data_bus[404]), .A2(n6212), .B1(
        i_data_bus[436]), .B2(n8041), .ZN(n8035) );
  ND2D1BWP30P140LVT U11762 ( .A1(n8036), .A2(n8035), .ZN(N1223) );
  AOI22D1BWP30P140LVT U11763 ( .A1(i_data_bus[406]), .A2(n6212), .B1(
        i_data_bus[470]), .B2(n7434), .ZN(n8038) );
  AOI22D1BWP30P140LVT U11764 ( .A1(i_data_bus[502]), .A2(n7443), .B1(
        i_data_bus[438]), .B2(n8041), .ZN(n8037) );
  ND2D1BWP30P140LVT U11765 ( .A1(n8038), .A2(n8037), .ZN(N1225) );
  AOI22D1BWP30P140LVT U11766 ( .A1(i_data_bus[501]), .A2(n7443), .B1(
        i_data_bus[405]), .B2(n6212), .ZN(n8040) );
  AOI22D1BWP30P140LVT U11767 ( .A1(i_data_bus[469]), .A2(n7434), .B1(
        i_data_bus[437]), .B2(n8041), .ZN(n8039) );
  ND2D1BWP30P140LVT U11768 ( .A1(n8040), .A2(n8039), .ZN(N1224) );
  AOI22D1BWP30P140LVT U11769 ( .A1(i_data_bus[459]), .A2(n7434), .B1(
        i_data_bus[491]), .B2(n7443), .ZN(n8043) );
  AOI22D1BWP30P140LVT U11770 ( .A1(i_data_bus[395]), .A2(n6212), .B1(
        i_data_bus[427]), .B2(n8041), .ZN(n8042) );
  ND2D1BWP30P140LVT U11771 ( .A1(n8043), .A2(n8042), .ZN(N1214) );
  AOI22D1BWP30P140LVT U11772 ( .A1(i_data_bus[620]), .A2(n10254), .B1(
        i_data_bus[588]), .B2(n10252), .ZN(n8045) );
  AOI22D1BWP30P140LVT U11773 ( .A1(i_data_bus[556]), .A2(n10253), .B1(
        i_data_bus[524]), .B2(n10245), .ZN(n8044) );
  ND2D1BWP30P140LVT U11774 ( .A1(n8045), .A2(n8044), .ZN(N9619) );
  AOI22D1BWP30P140LVT U11775 ( .A1(i_data_bus[545]), .A2(n10271), .B1(
        i_data_bus[577]), .B2(n10269), .ZN(n8047) );
  AOI22D1BWP30P140LVT U11776 ( .A1(i_data_bus[609]), .A2(n10270), .B1(
        i_data_bus[513]), .B2(n10272), .ZN(n8046) );
  ND2D1BWP30P140LVT U11777 ( .A1(n8047), .A2(n8046), .ZN(N8118) );
  AOI22D1BWP30P140LVT U11778 ( .A1(i_data_bus[478]), .A2(n8124), .B1(
        i_data_bus[446]), .B2(n8125), .ZN(n8049) );
  AOI22D1BWP30P140LVT U11779 ( .A1(i_data_bus[414]), .A2(n8122), .B1(
        i_data_bus[510]), .B2(n8123), .ZN(n8048) );
  ND2D1BWP30P140LVT U11780 ( .A1(n8049), .A2(n8048), .ZN(N2611) );
  AOI22D1BWP30P140LVT U11781 ( .A1(i_data_bus[403]), .A2(n8122), .B1(
        i_data_bus[467]), .B2(n8124), .ZN(n8051) );
  AOI22D1BWP30P140LVT U11782 ( .A1(i_data_bus[435]), .A2(n8125), .B1(
        i_data_bus[499]), .B2(n8123), .ZN(n8050) );
  ND2D1BWP30P140LVT U11783 ( .A1(n8051), .A2(n8050), .ZN(N2600) );
  AOI22D1BWP30P140LVT U11784 ( .A1(i_data_bus[401]), .A2(n8122), .B1(
        i_data_bus[433]), .B2(n8125), .ZN(n8053) );
  AOI22D1BWP30P140LVT U11785 ( .A1(i_data_bus[465]), .A2(n8124), .B1(
        i_data_bus[497]), .B2(n8123), .ZN(n8052) );
  ND2D1BWP30P140LVT U11786 ( .A1(n8053), .A2(n8052), .ZN(N2598) );
  AOI22D1BWP30P140LVT U11787 ( .A1(i_data_bus[398]), .A2(n8122), .B1(
        i_data_bus[462]), .B2(n8124), .ZN(n8055) );
  AOI22D1BWP30P140LVT U11788 ( .A1(i_data_bus[430]), .A2(n8125), .B1(
        i_data_bus[494]), .B2(n8123), .ZN(n8054) );
  ND2D1BWP30P140LVT U11789 ( .A1(n8055), .A2(n8054), .ZN(N2595) );
  AOI22D1BWP30P140LVT U11790 ( .A1(i_data_bus[397]), .A2(n8122), .B1(
        i_data_bus[429]), .B2(n8125), .ZN(n8057) );
  AOI22D1BWP30P140LVT U11791 ( .A1(i_data_bus[461]), .A2(n8124), .B1(
        i_data_bus[493]), .B2(n8123), .ZN(n8056) );
  ND2D1BWP30P140LVT U11792 ( .A1(n8057), .A2(n8056), .ZN(N2594) );
  AOI22D1BWP30P140LVT U11793 ( .A1(i_data_bus[425]), .A2(n8125), .B1(
        i_data_bus[393]), .B2(n8122), .ZN(n8059) );
  AOI22D1BWP30P140LVT U11794 ( .A1(i_data_bus[457]), .A2(n8124), .B1(
        i_data_bus[489]), .B2(n8123), .ZN(n8058) );
  ND2D1BWP30P140LVT U11795 ( .A1(n8059), .A2(n8058), .ZN(N2590) );
  AOI22D1BWP30P140LVT U11796 ( .A1(i_data_bus[423]), .A2(n8125), .B1(
        i_data_bus[455]), .B2(n8124), .ZN(n8061) );
  AOI22D1BWP30P140LVT U11797 ( .A1(i_data_bus[391]), .A2(n8122), .B1(
        i_data_bus[487]), .B2(n8123), .ZN(n8060) );
  ND2D1BWP30P140LVT U11798 ( .A1(n8061), .A2(n8060), .ZN(N2588) );
  AOI22D1BWP30P140LVT U11799 ( .A1(i_data_bus[451]), .A2(n8124), .B1(
        i_data_bus[387]), .B2(n8122), .ZN(n8063) );
  AOI22D1BWP30P140LVT U11800 ( .A1(i_data_bus[419]), .A2(n8125), .B1(
        i_data_bus[483]), .B2(n8123), .ZN(n8062) );
  ND2D1BWP30P140LVT U11801 ( .A1(n8063), .A2(n8062), .ZN(N2584) );
  AOI22D1BWP30P140LVT U11802 ( .A1(i_data_bus[416]), .A2(n8125), .B1(
        i_data_bus[384]), .B2(n8122), .ZN(n8065) );
  AOI22D1BWP30P140LVT U11803 ( .A1(i_data_bus[448]), .A2(n8124), .B1(
        i_data_bus[480]), .B2(n8123), .ZN(n8064) );
  ND2D1BWP30P140LVT U11804 ( .A1(n8065), .A2(n8064), .ZN(N2581) );
  AOI22D1BWP30P140LVT U11805 ( .A1(i_data_bus[1012]), .A2(n8205), .B1(
        i_data_bus[980]), .B2(n8207), .ZN(n8067) );
  AOI22D1BWP30P140LVT U11806 ( .A1(i_data_bus[948]), .A2(n8208), .B1(
        i_data_bus[916]), .B2(n8206), .ZN(n8066) );
  ND2D1BWP30P140LVT U11807 ( .A1(n8067), .A2(n8066), .ZN(N5677) );
  AOI22D1BWP30P140LVT U11808 ( .A1(i_data_bus[1008]), .A2(n8205), .B1(
        i_data_bus[976]), .B2(n8207), .ZN(n8069) );
  AOI22D1BWP30P140LVT U11809 ( .A1(i_data_bus[944]), .A2(n8208), .B1(
        i_data_bus[912]), .B2(n8206), .ZN(n8068) );
  ND2D1BWP30P140LVT U11810 ( .A1(n8069), .A2(n8068), .ZN(N5673) );
  AOI22D1BWP30P140LVT U11811 ( .A1(i_data_bus[932]), .A2(n8208), .B1(
        i_data_bus[964]), .B2(n8207), .ZN(n8071) );
  AOI22D1BWP30P140LVT U11812 ( .A1(i_data_bus[996]), .A2(n8205), .B1(
        i_data_bus[900]), .B2(n8206), .ZN(n8070) );
  ND2D1BWP30P140LVT U11813 ( .A1(n8071), .A2(n8070), .ZN(N5661) );
  AOI22D1BWP30P140LVT U11814 ( .A1(i_data_bus[619]), .A2(n10270), .B1(
        i_data_bus[587]), .B2(n10269), .ZN(n8073) );
  AOI22D1BWP30P140LVT U11815 ( .A1(i_data_bus[555]), .A2(n10271), .B1(
        i_data_bus[523]), .B2(n10272), .ZN(n8072) );
  ND2D1BWP30P140LVT U11816 ( .A1(n8073), .A2(n8072), .ZN(N8128) );
  AOI22D1BWP30P140LVT U11817 ( .A1(i_data_bus[959]), .A2(n8208), .B1(
        i_data_bus[991]), .B2(n8207), .ZN(n8075) );
  AOI22D1BWP30P140LVT U11818 ( .A1(i_data_bus[1023]), .A2(n8205), .B1(
        i_data_bus[927]), .B2(n8206), .ZN(n8074) );
  ND2D1BWP30P140LVT U11819 ( .A1(n8075), .A2(n8074), .ZN(N5688) );
  AOI22D1BWP30P140LVT U11820 ( .A1(i_data_bus[1014]), .A2(n8205), .B1(
        i_data_bus[982]), .B2(n8207), .ZN(n8077) );
  AOI22D1BWP30P140LVT U11821 ( .A1(i_data_bus[918]), .A2(n8206), .B1(
        i_data_bus[950]), .B2(n8208), .ZN(n8076) );
  ND2D1BWP30P140LVT U11822 ( .A1(n8077), .A2(n8076), .ZN(N5679) );
  AOI22D1BWP30P140LVT U11823 ( .A1(i_data_bus[922]), .A2(n8206), .B1(
        i_data_bus[986]), .B2(n8207), .ZN(n8079) );
  AOI22D1BWP30P140LVT U11824 ( .A1(i_data_bus[954]), .A2(n8208), .B1(
        i_data_bus[1018]), .B2(n8205), .ZN(n8078) );
  ND2D1BWP30P140LVT U11825 ( .A1(n8079), .A2(n8078), .ZN(N5683) );
  AOI22D1BWP30P140LVT U11826 ( .A1(i_data_bus[931]), .A2(n8208), .B1(
        i_data_bus[963]), .B2(n8207), .ZN(n8081) );
  AOI22D1BWP30P140LVT U11827 ( .A1(i_data_bus[899]), .A2(n8206), .B1(
        i_data_bus[995]), .B2(n8205), .ZN(n8080) );
  ND2D1BWP30P140LVT U11828 ( .A1(n8081), .A2(n8080), .ZN(N5660) );
  AOI22D1BWP30P140LVT U11829 ( .A1(i_data_bus[913]), .A2(n8206), .B1(
        i_data_bus[977]), .B2(n8207), .ZN(n8083) );
  AOI22D1BWP30P140LVT U11830 ( .A1(i_data_bus[945]), .A2(n8208), .B1(
        i_data_bus[1009]), .B2(n8205), .ZN(n8082) );
  ND2D1BWP30P140LVT U11831 ( .A1(n8083), .A2(n8082), .ZN(N5674) );
  AOI22D1BWP30P140LVT U11832 ( .A1(i_data_bus[919]), .A2(n8206), .B1(
        i_data_bus[983]), .B2(n8207), .ZN(n8085) );
  AOI22D1BWP30P140LVT U11833 ( .A1(i_data_bus[951]), .A2(n8208), .B1(
        i_data_bus[1015]), .B2(n8205), .ZN(n8084) );
  ND2D1BWP30P140LVT U11834 ( .A1(n8085), .A2(n8084), .ZN(N5680) );
  AOI22D1BWP30P140LVT U11835 ( .A1(i_data_bus[511]), .A2(n8123), .B1(
        i_data_bus[415]), .B2(n8122), .ZN(n8087) );
  AOI22D1BWP30P140LVT U11836 ( .A1(i_data_bus[479]), .A2(n8124), .B1(
        i_data_bus[447]), .B2(n8125), .ZN(n8086) );
  ND2D1BWP30P140LVT U11837 ( .A1(n8087), .A2(n8086), .ZN(N2612) );
  AOI22D1BWP30P140LVT U11838 ( .A1(i_data_bus[509]), .A2(n8123), .B1(
        i_data_bus[477]), .B2(n8124), .ZN(n8089) );
  AOI22D1BWP30P140LVT U11839 ( .A1(i_data_bus[413]), .A2(n8122), .B1(
        i_data_bus[445]), .B2(n8125), .ZN(n8088) );
  ND2D1BWP30P140LVT U11840 ( .A1(n8089), .A2(n8088), .ZN(N2610) );
  AOI22D1BWP30P140LVT U11841 ( .A1(i_data_bus[469]), .A2(n8124), .B1(
        i_data_bus[405]), .B2(n8122), .ZN(n8091) );
  AOI22D1BWP30P140LVT U11842 ( .A1(i_data_bus[501]), .A2(n8123), .B1(
        i_data_bus[437]), .B2(n8125), .ZN(n8090) );
  ND2D1BWP30P140LVT U11843 ( .A1(n8091), .A2(n8090), .ZN(N2602) );
  AOI22D1BWP30P140LVT U11844 ( .A1(i_data_bus[500]), .A2(n8123), .B1(
        i_data_bus[468]), .B2(n8124), .ZN(n8093) );
  AOI22D1BWP30P140LVT U11845 ( .A1(i_data_bus[404]), .A2(n8122), .B1(
        i_data_bus[436]), .B2(n8125), .ZN(n8092) );
  ND2D1BWP30P140LVT U11846 ( .A1(n8093), .A2(n8092), .ZN(N2601) );
  AOI22D1BWP30P140LVT U11847 ( .A1(i_data_bus[400]), .A2(n8122), .B1(
        i_data_bus[464]), .B2(n8124), .ZN(n8095) );
  AOI22D1BWP30P140LVT U11848 ( .A1(i_data_bus[496]), .A2(n8123), .B1(
        i_data_bus[432]), .B2(n8125), .ZN(n8094) );
  ND2D1BWP30P140LVT U11849 ( .A1(n8095), .A2(n8094), .ZN(N2597) );
  AOI22D1BWP30P140LVT U11850 ( .A1(i_data_bus[463]), .A2(n8124), .B1(
        i_data_bus[495]), .B2(n8123), .ZN(n8097) );
  AOI22D1BWP30P140LVT U11851 ( .A1(i_data_bus[399]), .A2(n8122), .B1(
        i_data_bus[431]), .B2(n8125), .ZN(n8096) );
  ND2D1BWP30P140LVT U11852 ( .A1(n8097), .A2(n8096), .ZN(N2596) );
  AOI22D1BWP30P140LVT U11853 ( .A1(i_data_bus[395]), .A2(n8122), .B1(
        i_data_bus[491]), .B2(n8123), .ZN(n8099) );
  AOI22D1BWP30P140LVT U11854 ( .A1(i_data_bus[459]), .A2(n8124), .B1(
        i_data_bus[427]), .B2(n8125), .ZN(n8098) );
  ND2D1BWP30P140LVT U11855 ( .A1(n8099), .A2(n8098), .ZN(N2592) );
  AOI22D1BWP30P140LVT U11856 ( .A1(i_data_bus[456]), .A2(n8124), .B1(
        i_data_bus[392]), .B2(n8122), .ZN(n8101) );
  AOI22D1BWP30P140LVT U11857 ( .A1(i_data_bus[488]), .A2(n8123), .B1(
        i_data_bus[424]), .B2(n8125), .ZN(n8100) );
  ND2D1BWP30P140LVT U11858 ( .A1(n8101), .A2(n8100), .ZN(N2589) );
  AOI22D1BWP30P140LVT U11859 ( .A1(i_data_bus[388]), .A2(n8122), .B1(
        i_data_bus[484]), .B2(n8123), .ZN(n8103) );
  AOI22D1BWP30P140LVT U11860 ( .A1(i_data_bus[452]), .A2(n8124), .B1(
        i_data_bus[420]), .B2(n8125), .ZN(n8102) );
  ND2D1BWP30P140LVT U11861 ( .A1(n8103), .A2(n8102), .ZN(N2585) );
  AOI22D1BWP30P140LVT U11862 ( .A1(i_data_bus[386]), .A2(n8122), .B1(
        i_data_bus[450]), .B2(n8124), .ZN(n8105) );
  AOI22D1BWP30P140LVT U11863 ( .A1(i_data_bus[482]), .A2(n8123), .B1(
        i_data_bus[418]), .B2(n8125), .ZN(n8104) );
  ND2D1BWP30P140LVT U11864 ( .A1(n8105), .A2(n8104), .ZN(N2583) );
  AOI22D1BWP30P140LVT U11865 ( .A1(i_data_bus[508]), .A2(n8123), .B1(
        i_data_bus[412]), .B2(n8122), .ZN(n8107) );
  AOI22D1BWP30P140LVT U11866 ( .A1(i_data_bus[444]), .A2(n8125), .B1(
        i_data_bus[476]), .B2(n8124), .ZN(n8106) );
  ND2D1BWP30P140LVT U11867 ( .A1(n8107), .A2(n8106), .ZN(N2609) );
  AOI22D1BWP30P140LVT U11868 ( .A1(i_data_bus[409]), .A2(n8122), .B1(
        i_data_bus[505]), .B2(n8123), .ZN(n8109) );
  AOI22D1BWP30P140LVT U11869 ( .A1(i_data_bus[441]), .A2(n8125), .B1(
        i_data_bus[473]), .B2(n8124), .ZN(n8108) );
  ND2D1BWP30P140LVT U11870 ( .A1(n8109), .A2(n8108), .ZN(N2606) );
  AOI22D1BWP30P140LVT U11871 ( .A1(i_data_bus[504]), .A2(n8123), .B1(
        i_data_bus[408]), .B2(n8122), .ZN(n8111) );
  AOI22D1BWP30P140LVT U11872 ( .A1(i_data_bus[440]), .A2(n8125), .B1(
        i_data_bus[472]), .B2(n8124), .ZN(n8110) );
  ND2D1BWP30P140LVT U11873 ( .A1(n8111), .A2(n8110), .ZN(N2605) );
  AOI22D1BWP30P140LVT U11874 ( .A1(i_data_bus[439]), .A2(n8125), .B1(
        i_data_bus[503]), .B2(n8123), .ZN(n8113) );
  AOI22D1BWP30P140LVT U11875 ( .A1(i_data_bus[407]), .A2(n8122), .B1(
        i_data_bus[471]), .B2(n8124), .ZN(n8112) );
  ND2D1BWP30P140LVT U11876 ( .A1(n8113), .A2(n8112), .ZN(N2604) );
  AOI22D1BWP30P140LVT U11877 ( .A1(i_data_bus[438]), .A2(n8125), .B1(
        i_data_bus[406]), .B2(n8122), .ZN(n8115) );
  AOI22D1BWP30P140LVT U11878 ( .A1(i_data_bus[502]), .A2(n8123), .B1(
        i_data_bus[470]), .B2(n8124), .ZN(n8114) );
  ND2D1BWP30P140LVT U11879 ( .A1(n8115), .A2(n8114), .ZN(N2603) );
  AOI22D1BWP30P140LVT U11880 ( .A1(i_data_bus[428]), .A2(n8125), .B1(
        i_data_bus[492]), .B2(n8123), .ZN(n8117) );
  AOI22D1BWP30P140LVT U11881 ( .A1(i_data_bus[396]), .A2(n8122), .B1(
        i_data_bus[460]), .B2(n8124), .ZN(n8116) );
  ND2D1BWP30P140LVT U11882 ( .A1(n8117), .A2(n8116), .ZN(N2593) );
  AOI22D1BWP30P140LVT U11883 ( .A1(i_data_bus[426]), .A2(n8125), .B1(
        i_data_bus[490]), .B2(n8123), .ZN(n8119) );
  AOI22D1BWP30P140LVT U11884 ( .A1(i_data_bus[394]), .A2(n8122), .B1(
        i_data_bus[458]), .B2(n8124), .ZN(n8118) );
  ND2D1BWP30P140LVT U11885 ( .A1(n8119), .A2(n8118), .ZN(N2591) );
  AOI22D1BWP30P140LVT U11886 ( .A1(i_data_bus[390]), .A2(n8122), .B1(
        i_data_bus[486]), .B2(n8123), .ZN(n8121) );
  AOI22D1BWP30P140LVT U11887 ( .A1(i_data_bus[422]), .A2(n8125), .B1(
        i_data_bus[454]), .B2(n8124), .ZN(n8120) );
  ND2D1BWP30P140LVT U11888 ( .A1(n8121), .A2(n8120), .ZN(N2587) );
  AOI22D1BWP30P140LVT U11889 ( .A1(i_data_bus[485]), .A2(n8123), .B1(
        i_data_bus[389]), .B2(n8122), .ZN(n8127) );
  AOI22D1BWP30P140LVT U11890 ( .A1(i_data_bus[421]), .A2(n8125), .B1(
        i_data_bus[453]), .B2(n8124), .ZN(n8126) );
  ND2D1BWP30P140LVT U11891 ( .A1(n8127), .A2(n8126), .ZN(N2586) );
  AOI22D1BWP30P140LVT U11892 ( .A1(i_data_bus[1010]), .A2(n8230), .B1(
        i_data_bus[978]), .B2(n8232), .ZN(n8129) );
  AOI22D1BWP30P140LVT U11893 ( .A1(i_data_bus[914]), .A2(n8233), .B1(
        i_data_bus[946]), .B2(n8231), .ZN(n8128) );
  ND2D1BWP30P140LVT U11894 ( .A1(n8129), .A2(n8128), .ZN(N8399) );
  AOI22D1BWP30P140LVT U11895 ( .A1(i_data_bus[950]), .A2(n8231), .B1(
        i_data_bus[982]), .B2(n8232), .ZN(n8131) );
  AOI22D1BWP30P140LVT U11896 ( .A1(i_data_bus[918]), .A2(n8233), .B1(
        i_data_bus[1014]), .B2(n8230), .ZN(n8130) );
  ND2D1BWP30P140LVT U11897 ( .A1(n8131), .A2(n8130), .ZN(N8403) );
  AOI22D1BWP30P140LVT U11898 ( .A1(i_data_bus[930]), .A2(n8231), .B1(
        i_data_bus[962]), .B2(n8232), .ZN(n8133) );
  AOI22D1BWP30P140LVT U11899 ( .A1(i_data_bus[898]), .A2(n8233), .B1(
        i_data_bus[994]), .B2(n8230), .ZN(n8132) );
  ND2D1BWP30P140LVT U11900 ( .A1(n8133), .A2(n8132), .ZN(N8383) );
  AOI22D1BWP30P140LVT U11901 ( .A1(i_data_bus[1021]), .A2(n8230), .B1(
        i_data_bus[989]), .B2(n8232), .ZN(n8135) );
  AOI22D1BWP30P140LVT U11902 ( .A1(i_data_bus[957]), .A2(n8231), .B1(
        i_data_bus[925]), .B2(n8233), .ZN(n8134) );
  ND2D1BWP30P140LVT U11903 ( .A1(n8135), .A2(n8134), .ZN(N8410) );
  AOI22D1BWP30P140LVT U11904 ( .A1(i_data_bus[913]), .A2(n8233), .B1(
        i_data_bus[977]), .B2(n8232), .ZN(n8137) );
  AOI22D1BWP30P140LVT U11905 ( .A1(i_data_bus[945]), .A2(n8231), .B1(
        i_data_bus[1009]), .B2(n8230), .ZN(n8136) );
  ND2D1BWP30P140LVT U11906 ( .A1(n8137), .A2(n8136), .ZN(N8398) );
  AOI22D1BWP30P140LVT U11907 ( .A1(i_data_bus[480]), .A2(n8194), .B1(
        i_data_bus[384]), .B2(n6224), .ZN(n8139) );
  AOI22D1BWP30P140LVT U11908 ( .A1(i_data_bus[416]), .A2(n8196), .B1(
        i_data_bus[448]), .B2(n8195), .ZN(n8138) );
  ND2D1BWP30P140LVT U11909 ( .A1(n8139), .A2(n8138), .ZN(N3943) );
  AOI22D1BWP30P140LVT U11910 ( .A1(i_data_bus[933]), .A2(n8256), .B1(
        i_data_bus[965]), .B2(n8257), .ZN(n8141) );
  AOI22D1BWP30P140LVT U11911 ( .A1(i_data_bus[901]), .A2(n8258), .B1(
        i_data_bus[997]), .B2(n8255), .ZN(n8140) );
  ND2D1BWP30P140LVT U11912 ( .A1(n8141), .A2(n8140), .ZN(N11110) );
  AOI22D1BWP30P140LVT U11913 ( .A1(i_data_bus[934]), .A2(n8256), .B1(
        i_data_bus[966]), .B2(n8257), .ZN(n8143) );
  AOI22D1BWP30P140LVT U11914 ( .A1(i_data_bus[902]), .A2(n8258), .B1(
        i_data_bus[998]), .B2(n8255), .ZN(n8142) );
  ND2D1BWP30P140LVT U11915 ( .A1(n8143), .A2(n8142), .ZN(N11111) );
  AOI22D1BWP30P140LVT U11916 ( .A1(i_data_bus[930]), .A2(n8256), .B1(
        i_data_bus[962]), .B2(n8257), .ZN(n8145) );
  AOI22D1BWP30P140LVT U11917 ( .A1(i_data_bus[898]), .A2(n8258), .B1(
        i_data_bus[994]), .B2(n8255), .ZN(n8144) );
  ND2D1BWP30P140LVT U11918 ( .A1(n8145), .A2(n8144), .ZN(N11107) );
  AOI22D1BWP30P140LVT U11919 ( .A1(i_data_bus[899]), .A2(n8258), .B1(
        i_data_bus[963]), .B2(n8257), .ZN(n8147) );
  AOI22D1BWP30P140LVT U11920 ( .A1(i_data_bus[995]), .A2(n8255), .B1(
        i_data_bus[931]), .B2(n8256), .ZN(n8146) );
  ND2D1BWP30P140LVT U11921 ( .A1(n8147), .A2(n8146), .ZN(N11108) );
  AOI22D1BWP30P140LVT U11922 ( .A1(i_data_bus[909]), .A2(n8258), .B1(
        i_data_bus[973]), .B2(n8257), .ZN(n8149) );
  AOI22D1BWP30P140LVT U11923 ( .A1(i_data_bus[1005]), .A2(n8255), .B1(
        i_data_bus[941]), .B2(n8256), .ZN(n8148) );
  ND2D1BWP30P140LVT U11924 ( .A1(n8149), .A2(n8148), .ZN(N11118) );
  AOI22D1BWP30P140LVT U11925 ( .A1(i_data_bus[918]), .A2(n8258), .B1(
        i_data_bus[982]), .B2(n8257), .ZN(n8151) );
  AOI22D1BWP30P140LVT U11926 ( .A1(i_data_bus[1014]), .A2(n8255), .B1(
        i_data_bus[950]), .B2(n8256), .ZN(n8150) );
  ND2D1BWP30P140LVT U11927 ( .A1(n8151), .A2(n8150), .ZN(N11127) );
  AOI22D1BWP30P140LVT U11928 ( .A1(i_data_bus[914]), .A2(n8258), .B1(
        i_data_bus[978]), .B2(n8257), .ZN(n8153) );
  AOI22D1BWP30P140LVT U11929 ( .A1(i_data_bus[1010]), .A2(n8255), .B1(
        i_data_bus[946]), .B2(n8256), .ZN(n8152) );
  ND2D1BWP30P140LVT U11930 ( .A1(n8153), .A2(n8152), .ZN(N11123) );
  AOI22D1BWP30P140LVT U11931 ( .A1(i_data_bus[922]), .A2(n8258), .B1(
        i_data_bus[986]), .B2(n8257), .ZN(n8155) );
  AOI22D1BWP30P140LVT U11932 ( .A1(i_data_bus[954]), .A2(n8256), .B1(
        i_data_bus[1018]), .B2(n8255), .ZN(n8154) );
  ND2D1BWP30P140LVT U11933 ( .A1(n8155), .A2(n8154), .ZN(N11131) );
  AOI22D1BWP30P140LVT U11934 ( .A1(i_data_bus[896]), .A2(n8258), .B1(
        i_data_bus[960]), .B2(n8257), .ZN(n8157) );
  AOI22D1BWP30P140LVT U11935 ( .A1(i_data_bus[928]), .A2(n8256), .B1(
        i_data_bus[992]), .B2(n8255), .ZN(n8156) );
  ND2D1BWP30P140LVT U11936 ( .A1(n8157), .A2(n8156), .ZN(N11105) );
  AOI22D1BWP30P140LVT U11937 ( .A1(i_data_bus[912]), .A2(n8258), .B1(
        i_data_bus[976]), .B2(n8257), .ZN(n8159) );
  AOI22D1BWP30P140LVT U11938 ( .A1(i_data_bus[944]), .A2(n8256), .B1(
        i_data_bus[1008]), .B2(n8255), .ZN(n8158) );
  ND2D1BWP30P140LVT U11939 ( .A1(n8159), .A2(n8158), .ZN(N11121) );
  AOI22D1BWP30P140LVT U11940 ( .A1(i_data_bus[921]), .A2(n8258), .B1(
        i_data_bus[985]), .B2(n8257), .ZN(n8161) );
  AOI22D1BWP30P140LVT U11941 ( .A1(i_data_bus[953]), .A2(n8256), .B1(
        i_data_bus[1017]), .B2(n8255), .ZN(n8160) );
  ND2D1BWP30P140LVT U11942 ( .A1(n8161), .A2(n8160), .ZN(N11130) );
  AOI22D1BWP30P140LVT U11943 ( .A1(i_data_bus[1022]), .A2(n8255), .B1(
        i_data_bus[990]), .B2(n8257), .ZN(n8163) );
  AOI22D1BWP30P140LVT U11944 ( .A1(i_data_bus[958]), .A2(n8256), .B1(
        i_data_bus[926]), .B2(n8258), .ZN(n8162) );
  ND2D1BWP30P140LVT U11945 ( .A1(n8163), .A2(n8162), .ZN(N11135) );
  AOI22D1BWP30P140LVT U11946 ( .A1(i_data_bus[1006]), .A2(n8339), .B1(
        i_data_bus[974]), .B2(n8341), .ZN(n8165) );
  AOI22D1BWP30P140LVT U11947 ( .A1(i_data_bus[910]), .A2(n8342), .B1(
        i_data_bus[942]), .B2(n8340), .ZN(n8164) );
  ND2D1BWP30P140LVT U11948 ( .A1(n8165), .A2(n8164), .ZN(N10269) );
  AOI22D1BWP30P140LVT U11949 ( .A1(i_data_bus[954]), .A2(n8351), .B1(
        i_data_bus[986]), .B2(n8353), .ZN(n8167) );
  AOI22D1BWP30P140LVT U11950 ( .A1(i_data_bus[922]), .A2(n8354), .B1(
        i_data_bus[1018]), .B2(n8352), .ZN(n8166) );
  ND2D1BWP30P140LVT U11951 ( .A1(n8167), .A2(n8166), .ZN(N4833) );
  AOI22D1BWP30P140LVT U11952 ( .A1(i_data_bus[1006]), .A2(n8352), .B1(
        i_data_bus[974]), .B2(n8353), .ZN(n8169) );
  AOI22D1BWP30P140LVT U11953 ( .A1(i_data_bus[910]), .A2(n8354), .B1(
        i_data_bus[942]), .B2(n8351), .ZN(n8168) );
  ND2D1BWP30P140LVT U11954 ( .A1(n8169), .A2(n8168), .ZN(N4821) );
  AOI22D1BWP30P140LVT U11955 ( .A1(i_data_bus[921]), .A2(n8354), .B1(
        i_data_bus[985]), .B2(n8353), .ZN(n8171) );
  AOI22D1BWP30P140LVT U11956 ( .A1(i_data_bus[953]), .A2(n8351), .B1(
        i_data_bus[1017]), .B2(n8352), .ZN(n8170) );
  ND2D1BWP30P140LVT U11957 ( .A1(n8171), .A2(n8170), .ZN(N4832) );
  AOI22D1BWP30P140LVT U11958 ( .A1(i_data_bus[915]), .A2(n8354), .B1(
        i_data_bus[979]), .B2(n8353), .ZN(n8173) );
  AOI22D1BWP30P140LVT U11959 ( .A1(i_data_bus[947]), .A2(n8351), .B1(
        i_data_bus[1011]), .B2(n8352), .ZN(n8172) );
  ND2D1BWP30P140LVT U11960 ( .A1(n8173), .A2(n8172), .ZN(N4826) );
  AOI22D1BWP30P140LVT U11961 ( .A1(i_data_bus[901]), .A2(n8354), .B1(
        i_data_bus[965]), .B2(n8353), .ZN(n8175) );
  AOI22D1BWP30P140LVT U11962 ( .A1(i_data_bus[933]), .A2(n8351), .B1(
        i_data_bus[997]), .B2(n8352), .ZN(n8174) );
  ND2D1BWP30P140LVT U11963 ( .A1(n8175), .A2(n8174), .ZN(N4812) );
  AOI22D1BWP30P140LVT U11964 ( .A1(i_data_bus[1023]), .A2(n8339), .B1(
        i_data_bus[991]), .B2(n8341), .ZN(n8177) );
  AOI22D1BWP30P140LVT U11965 ( .A1(i_data_bus[959]), .A2(n8340), .B1(
        i_data_bus[927]), .B2(n8342), .ZN(n8176) );
  ND2D1BWP30P140LVT U11966 ( .A1(n8177), .A2(n8176), .ZN(N10286) );
  AOI22D1BWP30P140LVT U11967 ( .A1(i_data_bus[1008]), .A2(n8339), .B1(
        i_data_bus[976]), .B2(n8341), .ZN(n8179) );
  AOI22D1BWP30P140LVT U11968 ( .A1(i_data_bus[944]), .A2(n8340), .B1(
        i_data_bus[912]), .B2(n8342), .ZN(n8178) );
  ND2D1BWP30P140LVT U11969 ( .A1(n8179), .A2(n8178), .ZN(N10271) );
  AOI22D1BWP30P140LVT U11970 ( .A1(i_data_bus[959]), .A2(n8351), .B1(
        i_data_bus[991]), .B2(n8353), .ZN(n8181) );
  AOI22D1BWP30P140LVT U11971 ( .A1(i_data_bus[1023]), .A2(n8352), .B1(
        i_data_bus[927]), .B2(n8354), .ZN(n8180) );
  ND2D1BWP30P140LVT U11972 ( .A1(n8181), .A2(n8180), .ZN(N4838) );
  AOI22D1BWP30P140LVT U11973 ( .A1(i_data_bus[1012]), .A2(n8352), .B1(
        i_data_bus[980]), .B2(n8353), .ZN(n8183) );
  AOI22D1BWP30P140LVT U11974 ( .A1(i_data_bus[948]), .A2(n8351), .B1(
        i_data_bus[916]), .B2(n8354), .ZN(n8182) );
  ND2D1BWP30P140LVT U11975 ( .A1(n8183), .A2(n8182), .ZN(N4827) );
  AOI22D1BWP30P140LVT U11976 ( .A1(i_data_bus[944]), .A2(n8351), .B1(
        i_data_bus[976]), .B2(n8353), .ZN(n8185) );
  AOI22D1BWP30P140LVT U11977 ( .A1(i_data_bus[1008]), .A2(n8352), .B1(
        i_data_bus[912]), .B2(n8354), .ZN(n8184) );
  ND2D1BWP30P140LVT U11978 ( .A1(n8185), .A2(n8184), .ZN(N4823) );
  AOI22D1BWP30P140LVT U11979 ( .A1(i_data_bus[996]), .A2(n8352), .B1(
        i_data_bus[964]), .B2(n8353), .ZN(n8187) );
  AOI22D1BWP30P140LVT U11980 ( .A1(i_data_bus[932]), .A2(n8351), .B1(
        i_data_bus[900]), .B2(n8354), .ZN(n8186) );
  ND2D1BWP30P140LVT U11981 ( .A1(n8187), .A2(n8186), .ZN(N4811) );
  AOI22D1BWP30P140LVT U11982 ( .A1(n8194), .A2(i_data_bus[489]), .B1(n6224), 
        .B2(i_data_bus[393]), .ZN(n8189) );
  AOI22D1BWP30P140LVT U11983 ( .A1(n8196), .A2(i_data_bus[425]), .B1(n8195), 
        .B2(i_data_bus[457]), .ZN(n8188) );
  ND2D1BWP30P140LVT U11984 ( .A1(n8189), .A2(n8188), .ZN(N3952) );
  AOI22D1BWP30P140LVT U11985 ( .A1(n8194), .A2(i_data_bus[484]), .B1(n6224), 
        .B2(i_data_bus[388]), .ZN(n8191) );
  AOI22D1BWP30P140LVT U11986 ( .A1(n8196), .A2(i_data_bus[420]), .B1(n8195), 
        .B2(i_data_bus[452]), .ZN(n8190) );
  ND2D1BWP30P140LVT U11987 ( .A1(n8191), .A2(n8190), .ZN(N3947) );
  AOI22D1BWP30P140LVT U11988 ( .A1(n8194), .A2(i_data_bus[483]), .B1(n6224), 
        .B2(i_data_bus[387]), .ZN(n8193) );
  AOI22D1BWP30P140LVT U11989 ( .A1(n8196), .A2(i_data_bus[419]), .B1(n8195), 
        .B2(i_data_bus[451]), .ZN(n8192) );
  ND2D1BWP30P140LVT U11990 ( .A1(n8193), .A2(n8192), .ZN(N3946) );
  AOI22D1BWP30P140LVT U11991 ( .A1(n8194), .A2(i_data_bus[481]), .B1(n6224), 
        .B2(i_data_bus[385]), .ZN(n8198) );
  AOI22D1BWP30P140LVT U11992 ( .A1(n8196), .A2(i_data_bus[417]), .B1(n8195), 
        .B2(i_data_bus[449]), .ZN(n8197) );
  ND2D1BWP30P140LVT U11993 ( .A1(n8198), .A2(n8197), .ZN(N3944) );
  AOI22D1BWP30P140LVT U11994 ( .A1(i_data_bus[898]), .A2(n8206), .B1(
        i_data_bus[994]), .B2(n8205), .ZN(n8200) );
  AOI22D1BWP30P140LVT U11995 ( .A1(i_data_bus[930]), .A2(n8208), .B1(
        i_data_bus[962]), .B2(n8207), .ZN(n8199) );
  ND2D1BWP30P140LVT U11996 ( .A1(n8200), .A2(n8199), .ZN(N5659) );
  AOI22D1BWP30P140LVT U11997 ( .A1(i_data_bus[921]), .A2(n8206), .B1(
        i_data_bus[953]), .B2(n8208), .ZN(n8202) );
  AOI22D1BWP30P140LVT U11998 ( .A1(i_data_bus[1017]), .A2(n8205), .B1(
        i_data_bus[985]), .B2(n8207), .ZN(n8201) );
  ND2D1BWP30P140LVT U11999 ( .A1(n8202), .A2(n8201), .ZN(N5682) );
  AOI22D1BWP30P140LVT U12000 ( .A1(i_data_bus[957]), .A2(n8208), .B1(
        i_data_bus[1021]), .B2(n8205), .ZN(n8204) );
  AOI22D1BWP30P140LVT U12001 ( .A1(i_data_bus[925]), .A2(n8206), .B1(
        i_data_bus[989]), .B2(n8207), .ZN(n8203) );
  ND2D1BWP30P140LVT U12002 ( .A1(n8204), .A2(n8203), .ZN(N5686) );
  AOI22D1BWP30P140LVT U12003 ( .A1(i_data_bus[896]), .A2(n8206), .B1(
        i_data_bus[992]), .B2(n8205), .ZN(n8210) );
  AOI22D1BWP30P140LVT U12004 ( .A1(i_data_bus[928]), .A2(n8208), .B1(
        i_data_bus[960]), .B2(n8207), .ZN(n8209) );
  ND2D1BWP30P140LVT U12005 ( .A1(n8210), .A2(n8209), .ZN(N5657) );
  AOI22D1BWP30P140LVT U12006 ( .A1(i_data_bus[959]), .A2(n8231), .B1(
        i_data_bus[927]), .B2(n8233), .ZN(n8212) );
  AOI22D1BWP30P140LVT U12007 ( .A1(i_data_bus[1023]), .A2(n8230), .B1(
        i_data_bus[991]), .B2(n8232), .ZN(n8211) );
  ND2D1BWP30P140LVT U12008 ( .A1(n8212), .A2(n8211), .ZN(N8412) );
  AOI22D1BWP30P140LVT U12009 ( .A1(i_data_bus[921]), .A2(n8233), .B1(
        i_data_bus[953]), .B2(n8231), .ZN(n8214) );
  AOI22D1BWP30P140LVT U12010 ( .A1(i_data_bus[1017]), .A2(n8230), .B1(
        i_data_bus[985]), .B2(n8232), .ZN(n8213) );
  ND2D1BWP30P140LVT U12011 ( .A1(n8214), .A2(n8213), .ZN(N8406) );
  AOI22D1BWP30P140LVT U12012 ( .A1(i_data_bus[919]), .A2(n8233), .B1(
        i_data_bus[1015]), .B2(n8230), .ZN(n8216) );
  AOI22D1BWP30P140LVT U12013 ( .A1(i_data_bus[951]), .A2(n8231), .B1(
        i_data_bus[983]), .B2(n8232), .ZN(n8215) );
  ND2D1BWP30P140LVT U12014 ( .A1(n8216), .A2(n8215), .ZN(N8404) );
  AOI22D1BWP30P140LVT U12015 ( .A1(i_data_bus[944]), .A2(n8231), .B1(
        i_data_bus[912]), .B2(n8233), .ZN(n8218) );
  AOI22D1BWP30P140LVT U12016 ( .A1(i_data_bus[1008]), .A2(n8230), .B1(
        i_data_bus[976]), .B2(n8232), .ZN(n8217) );
  ND2D1BWP30P140LVT U12017 ( .A1(n8218), .A2(n8217), .ZN(N8397) );
  AOI22D1BWP30P140LVT U12018 ( .A1(i_data_bus[910]), .A2(n8233), .B1(
        i_data_bus[942]), .B2(n8231), .ZN(n8220) );
  AOI22D1BWP30P140LVT U12019 ( .A1(i_data_bus[1006]), .A2(n8230), .B1(
        i_data_bus[974]), .B2(n8232), .ZN(n8219) );
  ND2D1BWP30P140LVT U12020 ( .A1(n8220), .A2(n8219), .ZN(N8395) );
  AOI22D1BWP30P140LVT U12021 ( .A1(i_data_bus[902]), .A2(n8233), .B1(
        i_data_bus[998]), .B2(n8230), .ZN(n8222) );
  AOI22D1BWP30P140LVT U12022 ( .A1(i_data_bus[934]), .A2(n8231), .B1(
        i_data_bus[966]), .B2(n8232), .ZN(n8221) );
  ND2D1BWP30P140LVT U12023 ( .A1(n8222), .A2(n8221), .ZN(N8387) );
  AOI22D1BWP30P140LVT U12024 ( .A1(i_data_bus[899]), .A2(n8233), .B1(
        i_data_bus[995]), .B2(n8230), .ZN(n8224) );
  AOI22D1BWP30P140LVT U12025 ( .A1(i_data_bus[931]), .A2(n8231), .B1(
        i_data_bus[963]), .B2(n8232), .ZN(n8223) );
  ND2D1BWP30P140LVT U12026 ( .A1(n8224), .A2(n8223), .ZN(N8384) );
  INR4D1BWP30P140LVT U12027 ( .A1(i_cmd[49]), .B1(i_cmd[33]), .B2(n10667), 
        .B3(n11138), .ZN(n10218) );
  NR4D1BWP30P140LVT U12028 ( .A1(i_cmd[41]), .A2(n10670), .A3(n11140), .A4(
        n8225), .ZN(n10220) );
  AOI22D1BWP30P140LVT U12029 ( .A1(i_data_bus[209]), .A2(n10218), .B1(
        i_data_bus[241]), .B2(n10220), .ZN(n8227) );
  NR4D1BWP30P140LVT U12030 ( .A1(i_cmd[57]), .A2(n11141), .A3(n10664), .A4(
        n8225), .ZN(n10219) );
  NR3D0P7BWP30P140LVT U12031 ( .A1(i_cmd[49]), .A2(i_cmd[41]), .A3(i_cmd[57]), 
        .ZN(n11137) );
  AOI22D1BWP30P140LVT U12032 ( .A1(i_data_bus[177]), .A2(n10219), .B1(
        i_data_bus[145]), .B2(n6213), .ZN(n8226) );
  ND2D1BWP30P140LVT U12033 ( .A1(n8227), .A2(n8226), .ZN(N2422) );
  AOI22D1BWP30P140LVT U12034 ( .A1(i_data_bus[947]), .A2(n8231), .B1(
        i_data_bus[1011]), .B2(n8230), .ZN(n8229) );
  AOI22D1BWP30P140LVT U12035 ( .A1(i_data_bus[915]), .A2(n8233), .B1(
        i_data_bus[979]), .B2(n8232), .ZN(n8228) );
  ND2D1BWP30P140LVT U12036 ( .A1(n8229), .A2(n8228), .ZN(N8400) );
  AOI22D1BWP30P140LVT U12037 ( .A1(i_data_bus[928]), .A2(n8231), .B1(
        i_data_bus[992]), .B2(n8230), .ZN(n8235) );
  AOI22D1BWP30P140LVT U12038 ( .A1(i_data_bus[896]), .A2(n8233), .B1(
        i_data_bus[960]), .B2(n8232), .ZN(n8234) );
  ND2D1BWP30P140LVT U12039 ( .A1(n8235), .A2(n8234), .ZN(N8381) );
  AOI22D1BWP30P140LVT U12040 ( .A1(i_data_bus[996]), .A2(n8255), .B1(
        i_data_bus[900]), .B2(n8258), .ZN(n8237) );
  AOI22D1BWP30P140LVT U12041 ( .A1(i_data_bus[932]), .A2(n8256), .B1(
        i_data_bus[964]), .B2(n8257), .ZN(n8236) );
  ND2D1BWP30P140LVT U12042 ( .A1(n8237), .A2(n8236), .ZN(N11109) );
  AOI22D1BWP30P140LVT U12043 ( .A1(i_data_bus[906]), .A2(n8258), .B1(
        i_data_bus[1002]), .B2(n8255), .ZN(n8239) );
  AOI22D1BWP30P140LVT U12044 ( .A1(i_data_bus[938]), .A2(n8256), .B1(
        i_data_bus[970]), .B2(n8257), .ZN(n8238) );
  ND2D1BWP30P140LVT U12045 ( .A1(n8239), .A2(n8238), .ZN(N11115) );
  AOI22D1BWP30P140LVT U12046 ( .A1(i_data_bus[957]), .A2(n8256), .B1(
        i_data_bus[925]), .B2(n8258), .ZN(n8241) );
  AOI22D1BWP30P140LVT U12047 ( .A1(i_data_bus[1021]), .A2(n8255), .B1(
        i_data_bus[989]), .B2(n8257), .ZN(n8240) );
  ND2D1BWP30P140LVT U12048 ( .A1(n8241), .A2(n8240), .ZN(N11134) );
  INR4D1BWP30P140LVT U12049 ( .A1(i_cmd[52]), .B1(i_cmd[36]), .B2(n10667), 
        .B3(n11044), .ZN(n10223) );
  NR4D1BWP30P140LVT U12050 ( .A1(i_cmd[44]), .A2(n10670), .A3(n8242), .A4(
        n8243), .ZN(n10226) );
  AOI22D1BWP30P140LVT U12051 ( .A1(i_data_bus[223]), .A2(n10223), .B1(
        i_data_bus[255]), .B2(n10226), .ZN(n8246) );
  NR4D1BWP30P140LVT U12052 ( .A1(i_cmd[60]), .A2(n8244), .A3(n10664), .A4(
        n8243), .ZN(n10225) );
  NR3D0P7BWP30P140LVT U12053 ( .A1(i_cmd[52]), .A2(i_cmd[44]), .A3(i_cmd[60]), 
        .ZN(n11040) );
  AOI22D1BWP30P140LVT U12054 ( .A1(i_data_bus[191]), .A2(n10225), .B1(
        i_data_bus[159]), .B2(n10224), .ZN(n8245) );
  ND2D1BWP30P140LVT U12055 ( .A1(n8246), .A2(n8245), .ZN(N6266) );
  AOI22D1BWP30P140LVT U12056 ( .A1(i_data_bus[177]), .A2(n10225), .B1(
        i_data_bus[241]), .B2(n10226), .ZN(n8248) );
  AOI22D1BWP30P140LVT U12057 ( .A1(i_data_bus[209]), .A2(n10223), .B1(
        i_data_bus[145]), .B2(n10224), .ZN(n8247) );
  ND2D1BWP30P140LVT U12058 ( .A1(n8248), .A2(n8247), .ZN(N6252) );
  AOI22D1BWP30P140LVT U12059 ( .A1(i_data_bus[173]), .A2(n10225), .B1(
        i_data_bus[237]), .B2(n10226), .ZN(n8250) );
  AOI22D1BWP30P140LVT U12060 ( .A1(i_data_bus[205]), .A2(n10223), .B1(
        i_data_bus[141]), .B2(n10224), .ZN(n8249) );
  ND2D1BWP30P140LVT U12061 ( .A1(n8250), .A2(n8249), .ZN(N6248) );
  AOI22D1BWP30P140LVT U12062 ( .A1(i_data_bus[164]), .A2(n10225), .B1(
        i_data_bus[228]), .B2(n10226), .ZN(n8252) );
  AOI22D1BWP30P140LVT U12063 ( .A1(i_data_bus[196]), .A2(n10223), .B1(
        i_data_bus[132]), .B2(n10224), .ZN(n8251) );
  ND2D1BWP30P140LVT U12064 ( .A1(n8252), .A2(n8251), .ZN(N6239) );
  AOI22D1BWP30P140LVT U12065 ( .A1(i_data_bus[162]), .A2(n10225), .B1(
        i_data_bus[226]), .B2(n10226), .ZN(n8254) );
  AOI22D1BWP30P140LVT U12066 ( .A1(i_data_bus[194]), .A2(n10223), .B1(
        i_data_bus[130]), .B2(n10224), .ZN(n8253) );
  ND2D1BWP30P140LVT U12067 ( .A1(n8254), .A2(n8253), .ZN(N6237) );
  AOI22D1BWP30P140LVT U12068 ( .A1(i_data_bus[940]), .A2(n8256), .B1(
        i_data_bus[1004]), .B2(n8255), .ZN(n8260) );
  AOI22D1BWP30P140LVT U12069 ( .A1(i_data_bus[908]), .A2(n8258), .B1(
        i_data_bus[972]), .B2(n8257), .ZN(n8259) );
  ND2D1BWP30P140LVT U12070 ( .A1(n8260), .A2(n8259), .ZN(N11117) );
  AOI22D1BWP30P140LVT U12071 ( .A1(n8720), .A2(i_data_bus[931]), .B1(n8721), 
        .B2(i_data_bus[963]), .ZN(n8262) );
  AOI22D1BWP30P140LVT U12072 ( .A1(n8722), .A2(i_data_bus[899]), .B1(n8719), 
        .B2(i_data_bus[995]), .ZN(n8261) );
  ND2D1BWP30P140LVT U12073 ( .A1(n8262), .A2(n8261), .ZN(N2936) );
  AOI22D1BWP30P140LVT U12074 ( .A1(n8722), .A2(i_data_bus[900]), .B1(n8721), 
        .B2(i_data_bus[964]), .ZN(n8264) );
  AOI22D1BWP30P140LVT U12075 ( .A1(n8720), .A2(i_data_bus[932]), .B1(n8719), 
        .B2(i_data_bus[996]), .ZN(n8263) );
  ND2D1BWP30P140LVT U12076 ( .A1(n8264), .A2(n8263), .ZN(N2937) );
  AOI22D1BWP30P140LVT U12077 ( .A1(n8722), .A2(i_data_bus[912]), .B1(n8721), 
        .B2(i_data_bus[976]), .ZN(n8266) );
  AOI22D1BWP30P140LVT U12078 ( .A1(n8720), .A2(i_data_bus[944]), .B1(n8719), 
        .B2(i_data_bus[1008]), .ZN(n8265) );
  ND2D1BWP30P140LVT U12079 ( .A1(n8266), .A2(n8265), .ZN(N2949) );
  AOI22D1BWP30P140LVT U12080 ( .A1(n8722), .A2(i_data_bus[927]), .B1(n8721), 
        .B2(i_data_bus[991]), .ZN(n8268) );
  AOI22D1BWP30P140LVT U12081 ( .A1(n8720), .A2(i_data_bus[959]), .B1(n8719), 
        .B2(i_data_bus[1023]), .ZN(n8267) );
  ND2D1BWP30P140LVT U12082 ( .A1(n8268), .A2(n8267), .ZN(N2964) );
  AOI22D1BWP30P140LVT U12083 ( .A1(n8722), .A2(i_data_bus[926]), .B1(n8721), 
        .B2(i_data_bus[990]), .ZN(n8270) );
  AOI22D1BWP30P140LVT U12084 ( .A1(n8720), .A2(i_data_bus[958]), .B1(n8719), 
        .B2(i_data_bus[1022]), .ZN(n8269) );
  ND2D1BWP30P140LVT U12085 ( .A1(n8270), .A2(n8269), .ZN(N2963) );
  AOI22D1BWP30P140LVT U12086 ( .A1(n8722), .A2(i_data_bus[925]), .B1(n8721), 
        .B2(i_data_bus[989]), .ZN(n8272) );
  AOI22D1BWP30P140LVT U12087 ( .A1(n8720), .A2(i_data_bus[957]), .B1(n8719), 
        .B2(i_data_bus[1021]), .ZN(n8271) );
  ND2D1BWP30P140LVT U12088 ( .A1(n8272), .A2(n8271), .ZN(N2962) );
  AOI22D1BWP30P140LVT U12089 ( .A1(n8720), .A2(i_data_bus[950]), .B1(n8721), 
        .B2(i_data_bus[982]), .ZN(n8274) );
  AOI22D1BWP30P140LVT U12090 ( .A1(n8722), .A2(i_data_bus[918]), .B1(n8719), 
        .B2(i_data_bus[1014]), .ZN(n8273) );
  ND2D1BWP30P140LVT U12091 ( .A1(n8274), .A2(n8273), .ZN(N2955) );
  AOI22D1BWP30P140LVT U12092 ( .A1(n8722), .A2(i_data_bus[916]), .B1(n8721), 
        .B2(i_data_bus[980]), .ZN(n8276) );
  AOI22D1BWP30P140LVT U12093 ( .A1(n8720), .A2(i_data_bus[948]), .B1(n8719), 
        .B2(i_data_bus[1012]), .ZN(n8275) );
  ND2D1BWP30P140LVT U12094 ( .A1(n8276), .A2(n8275), .ZN(N2953) );
  AOI22D1BWP30P140LVT U12095 ( .A1(n8720), .A2(i_data_bus[946]), .B1(n8721), 
        .B2(i_data_bus[978]), .ZN(n8278) );
  AOI22D1BWP30P140LVT U12096 ( .A1(n8722), .A2(i_data_bus[914]), .B1(n8719), 
        .B2(i_data_bus[1010]), .ZN(n8277) );
  ND2D1BWP30P140LVT U12097 ( .A1(n8278), .A2(n8277), .ZN(N2951) );
  INR4D1BWP30P140LVT U12098 ( .A1(i_cmd[50]), .B1(i_cmd[34]), .B2(n10667), 
        .B3(n11107), .ZN(n10033) );
  NR4D1BWP30P140LVT U12099 ( .A1(i_cmd[42]), .A2(n10670), .A3(n11109), .A4(
        n8279), .ZN(n10035) );
  AOI22D1BWP30P140LVT U12100 ( .A1(i_data_bus[223]), .A2(n10033), .B1(
        i_data_bus[255]), .B2(n10035), .ZN(n8281) );
  NR4D1BWP30P140LVT U12101 ( .A1(i_cmd[58]), .A2(n11110), .A3(n10664), .A4(
        n8279), .ZN(n10034) );
  NR3D0P7BWP30P140LVT U12102 ( .A1(i_cmd[42]), .A2(i_cmd[58]), .A3(i_cmd[50]), 
        .ZN(n11106) );
  AOI22D1BWP30P140LVT U12103 ( .A1(i_data_bus[191]), .A2(n10034), .B1(
        i_data_bus[159]), .B2(n10026), .ZN(n8280) );
  ND2D1BWP30P140LVT U12104 ( .A1(n8281), .A2(n8280), .ZN(N3542) );
  AOI22D1BWP30P140LVT U12105 ( .A1(i_data_bus[177]), .A2(n10034), .B1(
        i_data_bus[241]), .B2(n10035), .ZN(n8283) );
  AOI22D1BWP30P140LVT U12106 ( .A1(i_data_bus[209]), .A2(n10033), .B1(
        i_data_bus[145]), .B2(n10026), .ZN(n8282) );
  ND2D1BWP30P140LVT U12107 ( .A1(n8283), .A2(n8282), .ZN(N3528) );
  AOI22D1BWP30P140LVT U12108 ( .A1(i_data_bus[164]), .A2(n10034), .B1(
        i_data_bus[228]), .B2(n10035), .ZN(n8285) );
  AOI22D1BWP30P140LVT U12109 ( .A1(i_data_bus[196]), .A2(n10033), .B1(
        i_data_bus[132]), .B2(n10026), .ZN(n8284) );
  ND2D1BWP30P140LVT U12110 ( .A1(n8285), .A2(n8284), .ZN(N3515) );
  AOI22D1BWP30P140LVT U12111 ( .A1(i_data_bus[604]), .A2(n10252), .B1(
        i_data_bus[636]), .B2(n10254), .ZN(n8287) );
  AOI22D1BWP30P140LVT U12112 ( .A1(i_data_bus[572]), .A2(n10253), .B1(
        i_data_bus[540]), .B2(n10245), .ZN(n8286) );
  ND2D1BWP30P140LVT U12113 ( .A1(n8287), .A2(n8286), .ZN(N9635) );
  AOI22D1BWP30P140LVT U12114 ( .A1(i_data_bus[567]), .A2(n10253), .B1(
        i_data_bus[631]), .B2(n10254), .ZN(n8289) );
  AOI22D1BWP30P140LVT U12115 ( .A1(i_data_bus[535]), .A2(n10245), .B1(
        i_data_bus[599]), .B2(n10252), .ZN(n8288) );
  ND2D1BWP30P140LVT U12116 ( .A1(n8289), .A2(n8288), .ZN(N9630) );
  AOI22D1BWP30P140LVT U12117 ( .A1(i_data_bus[531]), .A2(n10245), .B1(
        i_data_bus[627]), .B2(n10254), .ZN(n8291) );
  AOI22D1BWP30P140LVT U12118 ( .A1(i_data_bus[563]), .A2(n10253), .B1(
        i_data_bus[595]), .B2(n10252), .ZN(n8290) );
  ND2D1BWP30P140LVT U12119 ( .A1(n8291), .A2(n8290), .ZN(N9626) );
  AOI22D1BWP30P140LVT U12120 ( .A1(i_data_bus[561]), .A2(n10253), .B1(
        i_data_bus[625]), .B2(n10254), .ZN(n8293) );
  AOI22D1BWP30P140LVT U12121 ( .A1(i_data_bus[529]), .A2(n10245), .B1(
        i_data_bus[593]), .B2(n10252), .ZN(n8292) );
  ND2D1BWP30P140LVT U12122 ( .A1(n8293), .A2(n8292), .ZN(N9624) );
  AOI22D1BWP30P140LVT U12123 ( .A1(i_data_bus[919]), .A2(n8342), .B1(
        i_data_bus[1015]), .B2(n8339), .ZN(n8295) );
  AOI22D1BWP30P140LVT U12124 ( .A1(i_data_bus[951]), .A2(n8340), .B1(
        i_data_bus[983]), .B2(n8341), .ZN(n8294) );
  ND2D1BWP30P140LVT U12125 ( .A1(n8295), .A2(n8294), .ZN(N10278) );
  AOI22D1BWP30P140LVT U12126 ( .A1(i_data_bus[996]), .A2(n8339), .B1(
        i_data_bus[900]), .B2(n8342), .ZN(n8297) );
  AOI22D1BWP30P140LVT U12127 ( .A1(i_data_bus[932]), .A2(n8340), .B1(
        i_data_bus[964]), .B2(n8341), .ZN(n8296) );
  ND2D1BWP30P140LVT U12128 ( .A1(n8297), .A2(n8296), .ZN(N10259) );
  AOI22D1BWP30P140LVT U12129 ( .A1(i_data_bus[899]), .A2(n8354), .B1(
        i_data_bus[931]), .B2(n8351), .ZN(n8299) );
  AOI22D1BWP30P140LVT U12130 ( .A1(i_data_bus[995]), .A2(n8352), .B1(
        i_data_bus[963]), .B2(n8353), .ZN(n8298) );
  ND2D1BWP30P140LVT U12131 ( .A1(n8299), .A2(n8298), .ZN(N4810) );
  AOI22D1BWP30P140LVT U12132 ( .A1(i_data_bus[898]), .A2(n8342), .B1(
        i_data_bus[994]), .B2(n8339), .ZN(n8301) );
  AOI22D1BWP30P140LVT U12133 ( .A1(i_data_bus[930]), .A2(n8340), .B1(
        i_data_bus[962]), .B2(n8341), .ZN(n8300) );
  ND2D1BWP30P140LVT U12134 ( .A1(n8301), .A2(n8300), .ZN(N10257) );
  AOI22D1BWP30P140LVT U12135 ( .A1(i_data_bus[957]), .A2(n8351), .B1(
        i_data_bus[925]), .B2(n8354), .ZN(n8303) );
  AOI22D1BWP30P140LVT U12136 ( .A1(i_data_bus[1021]), .A2(n8352), .B1(
        i_data_bus[989]), .B2(n8353), .ZN(n8302) );
  ND2D1BWP30P140LVT U12137 ( .A1(n8303), .A2(n8302), .ZN(N4836) );
  AOI22D1BWP30P140LVT U12138 ( .A1(i_data_bus[911]), .A2(n8354), .B1(
        i_data_bus[1007]), .B2(n8352), .ZN(n8305) );
  AOI22D1BWP30P140LVT U12139 ( .A1(i_data_bus[943]), .A2(n8351), .B1(
        i_data_bus[975]), .B2(n8353), .ZN(n8304) );
  ND2D1BWP30P140LVT U12140 ( .A1(n8305), .A2(n8304), .ZN(N4822) );
  AOI22D1BWP30P140LVT U12141 ( .A1(i_data_bus[1003]), .A2(n8352), .B1(
        i_data_bus[907]), .B2(n8354), .ZN(n8307) );
  AOI22D1BWP30P140LVT U12142 ( .A1(i_data_bus[939]), .A2(n8351), .B1(
        i_data_bus[971]), .B2(n8353), .ZN(n8306) );
  ND2D1BWP30P140LVT U12143 ( .A1(n8307), .A2(n8306), .ZN(N4818) );
  AOI22D1BWP30P140LVT U12144 ( .A1(i_data_bus[902]), .A2(n8354), .B1(
        i_data_bus[998]), .B2(n8352), .ZN(n8309) );
  AOI22D1BWP30P140LVT U12145 ( .A1(i_data_bus[934]), .A2(n8351), .B1(
        i_data_bus[966]), .B2(n8353), .ZN(n8308) );
  ND2D1BWP30P140LVT U12146 ( .A1(n8309), .A2(n8308), .ZN(N4813) );
  AOI22D1BWP30P140LVT U12147 ( .A1(i_data_bus[948]), .A2(n8340), .B1(
        i_data_bus[916]), .B2(n8342), .ZN(n8311) );
  AOI22D1BWP30P140LVT U12148 ( .A1(i_data_bus[1012]), .A2(n8339), .B1(
        i_data_bus[980]), .B2(n8341), .ZN(n8310) );
  ND2D1BWP30P140LVT U12149 ( .A1(n8311), .A2(n8310), .ZN(N10275) );
  AOI22D1BWP30P140LVT U12150 ( .A1(i_data_bus[911]), .A2(n8342), .B1(
        i_data_bus[1007]), .B2(n8339), .ZN(n8313) );
  AOI22D1BWP30P140LVT U12151 ( .A1(i_data_bus[943]), .A2(n8340), .B1(
        i_data_bus[975]), .B2(n8341), .ZN(n8312) );
  ND2D1BWP30P140LVT U12152 ( .A1(n8313), .A2(n8312), .ZN(N10270) );
  AOI22D1BWP30P140LVT U12153 ( .A1(i_data_bus[899]), .A2(n8342), .B1(
        i_data_bus[995]), .B2(n8339), .ZN(n8315) );
  AOI22D1BWP30P140LVT U12154 ( .A1(i_data_bus[931]), .A2(n8340), .B1(
        i_data_bus[963]), .B2(n8341), .ZN(n8314) );
  ND2D1BWP30P140LVT U12155 ( .A1(n8315), .A2(n8314), .ZN(N10258) );
  AOI22D1BWP30P140LVT U12156 ( .A1(i_data_bus[1022]), .A2(n8339), .B1(
        i_data_bus[926]), .B2(n8342), .ZN(n8317) );
  AOI22D1BWP30P140LVT U12157 ( .A1(i_data_bus[958]), .A2(n8340), .B1(
        i_data_bus[990]), .B2(n8341), .ZN(n8316) );
  ND2D1BWP30P140LVT U12158 ( .A1(n8317), .A2(n8316), .ZN(N10285) );
  INR4D1BWP30P140LVT U12159 ( .A1(i_cmd[54]), .B1(i_cmd[38]), .B2(n10667), 
        .B3(n8318), .ZN(n10039) );
  NR4D1BWP30P140LVT U12160 ( .A1(i_cmd[46]), .A2(n10670), .A3(n8319), .A4(
        n8320), .ZN(n10038) );
  AOI22D1BWP30P140LVT U12161 ( .A1(i_data_bus[196]), .A2(n10039), .B1(
        i_data_bus[228]), .B2(n10038), .ZN(n8324) );
  NR4D1BWP30P140LVT U12162 ( .A1(i_cmd[62]), .A2(n8321), .A3(n10664), .A4(
        n8320), .ZN(n10040) );
  AOI22D1BWP30P140LVT U12163 ( .A1(i_data_bus[164]), .A2(n10040), .B1(
        i_data_bus[132]), .B2(n9318), .ZN(n8323) );
  ND2D1BWP30P140LVT U12164 ( .A1(n8324), .A2(n8323), .ZN(N8963) );
  AOI22D1BWP30P140LVT U12165 ( .A1(i_data_bus[957]), .A2(n8340), .B1(
        i_data_bus[1021]), .B2(n8339), .ZN(n8326) );
  AOI22D1BWP30P140LVT U12166 ( .A1(i_data_bus[925]), .A2(n8342), .B1(
        i_data_bus[989]), .B2(n8341), .ZN(n8325) );
  ND2D1BWP30P140LVT U12167 ( .A1(n8326), .A2(n8325), .ZN(N10284) );
  AOI22D1BWP30P140LVT U12168 ( .A1(i_data_bus[954]), .A2(n8340), .B1(
        i_data_bus[1018]), .B2(n8339), .ZN(n8328) );
  AOI22D1BWP30P140LVT U12169 ( .A1(i_data_bus[922]), .A2(n8342), .B1(
        i_data_bus[986]), .B2(n8341), .ZN(n8327) );
  ND2D1BWP30P140LVT U12170 ( .A1(n8328), .A2(n8327), .ZN(N10281) );
  AOI22D1BWP30P140LVT U12171 ( .A1(i_data_bus[1014]), .A2(n8339), .B1(
        i_data_bus[950]), .B2(n8340), .ZN(n8330) );
  AOI22D1BWP30P140LVT U12172 ( .A1(i_data_bus[918]), .A2(n8342), .B1(
        i_data_bus[982]), .B2(n8341), .ZN(n8329) );
  ND2D1BWP30P140LVT U12173 ( .A1(n8330), .A2(n8329), .ZN(N10277) );
  AOI22D1BWP30P140LVT U12174 ( .A1(i_data_bus[953]), .A2(n8340), .B1(
        i_data_bus[1017]), .B2(n8339), .ZN(n8332) );
  AOI22D1BWP30P140LVT U12175 ( .A1(i_data_bus[921]), .A2(n8342), .B1(
        i_data_bus[985]), .B2(n8341), .ZN(n8331) );
  ND2D1BWP30P140LVT U12176 ( .A1(n8332), .A2(n8331), .ZN(N10280) );
  AOI22D1BWP30P140LVT U12177 ( .A1(i_data_bus[938]), .A2(n8340), .B1(
        i_data_bus[1002]), .B2(n8339), .ZN(n8334) );
  AOI22D1BWP30P140LVT U12178 ( .A1(i_data_bus[906]), .A2(n8342), .B1(
        i_data_bus[970]), .B2(n8341), .ZN(n8333) );
  ND2D1BWP30P140LVT U12179 ( .A1(n8334), .A2(n8333), .ZN(N10265) );
  AOI22D1BWP30P140LVT U12180 ( .A1(i_data_bus[955]), .A2(n8340), .B1(
        i_data_bus[1019]), .B2(n8339), .ZN(n8336) );
  AOI22D1BWP30P140LVT U12181 ( .A1(i_data_bus[923]), .A2(n8342), .B1(
        i_data_bus[987]), .B2(n8341), .ZN(n8335) );
  ND2D1BWP30P140LVT U12182 ( .A1(n8336), .A2(n8335), .ZN(N10282) );
  AOI22D1BWP30P140LVT U12183 ( .A1(i_data_bus[928]), .A2(n8340), .B1(
        i_data_bus[992]), .B2(n8339), .ZN(n8338) );
  AOI22D1BWP30P140LVT U12184 ( .A1(i_data_bus[896]), .A2(n8342), .B1(
        i_data_bus[960]), .B2(n8341), .ZN(n8337) );
  ND2D1BWP30P140LVT U12185 ( .A1(n8338), .A2(n8337), .ZN(N10255) );
  AOI22D1BWP30P140LVT U12186 ( .A1(i_data_bus[947]), .A2(n8340), .B1(
        i_data_bus[1011]), .B2(n8339), .ZN(n8344) );
  AOI22D1BWP30P140LVT U12187 ( .A1(i_data_bus[915]), .A2(n8342), .B1(
        i_data_bus[979]), .B2(n8341), .ZN(n8343) );
  ND2D1BWP30P140LVT U12188 ( .A1(n8344), .A2(n8343), .ZN(N10274) );
  AOI22D1BWP30P140LVT U12189 ( .A1(i_data_bus[1005]), .A2(n8352), .B1(
        i_data_bus[941]), .B2(n8351), .ZN(n8346) );
  AOI22D1BWP30P140LVT U12190 ( .A1(i_data_bus[909]), .A2(n8354), .B1(
        i_data_bus[973]), .B2(n8353), .ZN(n8345) );
  ND2D1BWP30P140LVT U12191 ( .A1(n8346), .A2(n8345), .ZN(N4820) );
  AOI22D1BWP30P140LVT U12192 ( .A1(i_data_bus[930]), .A2(n8351), .B1(
        i_data_bus[994]), .B2(n8352), .ZN(n8348) );
  AOI22D1BWP30P140LVT U12193 ( .A1(i_data_bus[898]), .A2(n8354), .B1(
        i_data_bus[962]), .B2(n8353), .ZN(n8347) );
  ND2D1BWP30P140LVT U12194 ( .A1(n8348), .A2(n8347), .ZN(N4809) );
  AOI22D1BWP30P140LVT U12195 ( .A1(i_data_bus[1014]), .A2(n8352), .B1(
        i_data_bus[950]), .B2(n8351), .ZN(n8350) );
  AOI22D1BWP30P140LVT U12196 ( .A1(i_data_bus[918]), .A2(n8354), .B1(
        i_data_bus[982]), .B2(n8353), .ZN(n8349) );
  ND2D1BWP30P140LVT U12197 ( .A1(n8350), .A2(n8349), .ZN(N4829) );
  AOI22D1BWP30P140LVT U12198 ( .A1(i_data_bus[1010]), .A2(n8352), .B1(
        i_data_bus[946]), .B2(n8351), .ZN(n8356) );
  AOI22D1BWP30P140LVT U12199 ( .A1(i_data_bus[914]), .A2(n8354), .B1(
        i_data_bus[978]), .B2(n8353), .ZN(n8355) );
  ND2D1BWP30P140LVT U12200 ( .A1(n8356), .A2(n8355), .ZN(N4825) );
  AOI22D1BWP30P140LVT U12201 ( .A1(i_data_bus[562]), .A2(n10002), .B1(
        i_data_bus[626]), .B2(n10003), .ZN(n8358) );
  AOI22D1BWP30P140LVT U12202 ( .A1(i_data_bus[530]), .A2(n6222), .B1(
        i_data_bus[594]), .B2(n10001), .ZN(n8357) );
  ND2D1BWP30P140LVT U12203 ( .A1(n8358), .A2(n8357), .ZN(N4177) );
  AOI22D1BWP30P140LVT U12204 ( .A1(i_data_bus[556]), .A2(n10002), .B1(
        i_data_bus[620]), .B2(n10003), .ZN(n8360) );
  AOI22D1BWP30P140LVT U12205 ( .A1(i_data_bus[524]), .A2(n6222), .B1(
        i_data_bus[588]), .B2(n10001), .ZN(n8359) );
  ND2D1BWP30P140LVT U12206 ( .A1(n8360), .A2(n8359), .ZN(N4171) );
  AOI22D1BWP30P140LVT U12207 ( .A1(i_data_bus[553]), .A2(n10002), .B1(
        i_data_bus[617]), .B2(n10003), .ZN(n8362) );
  AOI22D1BWP30P140LVT U12208 ( .A1(i_data_bus[521]), .A2(n6222), .B1(
        i_data_bus[585]), .B2(n10001), .ZN(n8361) );
  ND2D1BWP30P140LVT U12209 ( .A1(n8362), .A2(n8361), .ZN(N4168) );
  AOI22D1BWP30P140LVT U12210 ( .A1(i_data_bus[548]), .A2(n10002), .B1(
        i_data_bus[612]), .B2(n10003), .ZN(n8364) );
  AOI22D1BWP30P140LVT U12211 ( .A1(i_data_bus[516]), .A2(n6222), .B1(
        i_data_bus[580]), .B2(n10001), .ZN(n8363) );
  ND2D1BWP30P140LVT U12212 ( .A1(n8364), .A2(n8363), .ZN(N4163) );
  INR4D1BWP30P140LVT U12213 ( .A1(i_cmd[53]), .B1(i_cmd[37]), .B2(n10667), 
        .B3(n11008), .ZN(n10132) );
  NR4D1BWP30P140LVT U12214 ( .A1(i_cmd[45]), .A2(n10670), .A3(n8365), .A4(
        n8366), .ZN(n10131) );
  AOI22D1BWP30P140LVT U12215 ( .A1(i_data_bus[223]), .A2(n10132), .B1(
        i_data_bus[255]), .B2(n10131), .ZN(n8369) );
  NR4D1BWP30P140LVT U12216 ( .A1(i_cmd[61]), .A2(n8367), .A3(n10664), .A4(
        n8366), .ZN(n10133) );
  NR3D0P7BWP30P140LVT U12217 ( .A1(i_cmd[53]), .A2(i_cmd[45]), .A3(i_cmd[61]), 
        .ZN(n11004) );
  AOI22D1BWP30P140LVT U12218 ( .A1(i_data_bus[191]), .A2(n10133), .B1(
        i_data_bus[159]), .B2(n10134), .ZN(n8368) );
  ND2D1BWP30P140LVT U12219 ( .A1(n8369), .A2(n8368), .ZN(N7884) );
  AOI22D1BWP30P140LVT U12220 ( .A1(i_data_bus[196]), .A2(n10132), .B1(
        i_data_bus[228]), .B2(n10131), .ZN(n8371) );
  AOI22D1BWP30P140LVT U12221 ( .A1(i_data_bus[164]), .A2(n10133), .B1(
        i_data_bus[132]), .B2(n10134), .ZN(n8370) );
  ND2D1BWP30P140LVT U12222 ( .A1(n8371), .A2(n8370), .ZN(N7857) );
  AOI22D1BWP30P140LVT U12223 ( .A1(i_data_bus[173]), .A2(n10133), .B1(
        i_data_bus[237]), .B2(n10131), .ZN(n8373) );
  AOI22D1BWP30P140LVT U12224 ( .A1(i_data_bus[205]), .A2(n10132), .B1(
        i_data_bus[141]), .B2(n10134), .ZN(n8372) );
  ND2D1BWP30P140LVT U12225 ( .A1(n8373), .A2(n8372), .ZN(N7866) );
  AOI22D1BWP30P140LVT U12226 ( .A1(i_data_bus[389]), .A2(n10387), .B1(
        i_data_bus[453]), .B2(n10388), .ZN(n8379) );
  AOI22D1BWP30P140LVT U12227 ( .A1(i_data_bus[485]), .A2(n10385), .B1(
        i_data_bus[421]), .B2(n10386), .ZN(n8378) );
  ND2D1BWP30P140LVT U12228 ( .A1(n8379), .A2(n8378), .ZN(N10758) );
  AOI22D1BWP30P140LVT U12229 ( .A1(i_data_bus[414]), .A2(n10387), .B1(
        i_data_bus[478]), .B2(n10388), .ZN(n8381) );
  AOI22D1BWP30P140LVT U12230 ( .A1(i_data_bus[446]), .A2(n10386), .B1(
        i_data_bus[510]), .B2(n10385), .ZN(n8380) );
  ND2D1BWP30P140LVT U12231 ( .A1(n8381), .A2(n8380), .ZN(N10783) );
  AOI22D1BWP30P140LVT U12232 ( .A1(i_data_bus[412]), .A2(n10387), .B1(
        i_data_bus[476]), .B2(n10388), .ZN(n8383) );
  AOI22D1BWP30P140LVT U12233 ( .A1(i_data_bus[444]), .A2(n10386), .B1(
        i_data_bus[508]), .B2(n10385), .ZN(n8382) );
  ND2D1BWP30P140LVT U12234 ( .A1(n8383), .A2(n8382), .ZN(N10781) );
  AOI22D1BWP30P140LVT U12235 ( .A1(i_data_bus[409]), .A2(n10387), .B1(
        i_data_bus[473]), .B2(n10388), .ZN(n8385) );
  AOI22D1BWP30P140LVT U12236 ( .A1(i_data_bus[441]), .A2(n10386), .B1(
        i_data_bus[505]), .B2(n10385), .ZN(n8384) );
  ND2D1BWP30P140LVT U12237 ( .A1(n8385), .A2(n8384), .ZN(N10778) );
  AOI22D1BWP30P140LVT U12238 ( .A1(i_data_bus[408]), .A2(n10387), .B1(
        i_data_bus[472]), .B2(n10388), .ZN(n8387) );
  AOI22D1BWP30P140LVT U12239 ( .A1(i_data_bus[440]), .A2(n10386), .B1(
        i_data_bus[504]), .B2(n10385), .ZN(n8386) );
  ND2D1BWP30P140LVT U12240 ( .A1(n8387), .A2(n8386), .ZN(N10777) );
  AOI22D1BWP30P140LVT U12241 ( .A1(i_data_bus[404]), .A2(n10387), .B1(
        i_data_bus[468]), .B2(n10388), .ZN(n8389) );
  AOI22D1BWP30P140LVT U12242 ( .A1(i_data_bus[436]), .A2(n10386), .B1(
        i_data_bus[500]), .B2(n10385), .ZN(n8388) );
  ND2D1BWP30P140LVT U12243 ( .A1(n8389), .A2(n8388), .ZN(N10773) );
  AOI22D1BWP30P140LVT U12244 ( .A1(i_data_bus[396]), .A2(n10387), .B1(
        i_data_bus[460]), .B2(n10388), .ZN(n8391) );
  AOI22D1BWP30P140LVT U12245 ( .A1(i_data_bus[428]), .A2(n10386), .B1(
        i_data_bus[492]), .B2(n10385), .ZN(n8390) );
  ND2D1BWP30P140LVT U12246 ( .A1(n8391), .A2(n8390), .ZN(N10765) );
  AOI22D1BWP30P140LVT U12247 ( .A1(i_data_bus[407]), .A2(n10387), .B1(
        i_data_bus[439]), .B2(n10386), .ZN(n8393) );
  AOI22D1BWP30P140LVT U12248 ( .A1(i_data_bus[471]), .A2(n10388), .B1(
        i_data_bus[503]), .B2(n10385), .ZN(n8392) );
  ND2D1BWP30P140LVT U12249 ( .A1(n8393), .A2(n8392), .ZN(N10776) );
  AOI22D1BWP30P140LVT U12250 ( .A1(i_data_bus[401]), .A2(n10387), .B1(
        i_data_bus[433]), .B2(n10386), .ZN(n8395) );
  AOI22D1BWP30P140LVT U12251 ( .A1(i_data_bus[465]), .A2(n10388), .B1(
        i_data_bus[497]), .B2(n10385), .ZN(n8394) );
  ND2D1BWP30P140LVT U12252 ( .A1(n8395), .A2(n8394), .ZN(N10770) );
  AOI22D1BWP30P140LVT U12253 ( .A1(i_data_bus[399]), .A2(n10387), .B1(
        i_data_bus[431]), .B2(n10386), .ZN(n8397) );
  AOI22D1BWP30P140LVT U12254 ( .A1(i_data_bus[463]), .A2(n10388), .B1(
        i_data_bus[495]), .B2(n10385), .ZN(n8396) );
  ND2D1BWP30P140LVT U12255 ( .A1(n8397), .A2(n8396), .ZN(N10768) );
  AOI22D1BWP30P140LVT U12256 ( .A1(i_data_bus[386]), .A2(n10387), .B1(
        i_data_bus[418]), .B2(n10386), .ZN(n8399) );
  AOI22D1BWP30P140LVT U12257 ( .A1(i_data_bus[450]), .A2(n10388), .B1(
        i_data_bus[482]), .B2(n10385), .ZN(n8398) );
  ND2D1BWP30P140LVT U12258 ( .A1(n8399), .A2(n8398), .ZN(N10755) );
  AOI22D1BWP30P140LVT U12259 ( .A1(i_data_bus[398]), .A2(n10387), .B1(
        i_data_bus[494]), .B2(n10385), .ZN(n8401) );
  AOI22D1BWP30P140LVT U12260 ( .A1(i_data_bus[430]), .A2(n10386), .B1(
        i_data_bus[462]), .B2(n10388), .ZN(n8400) );
  ND2D1BWP30P140LVT U12261 ( .A1(n8401), .A2(n8400), .ZN(N10767) );
  AOI22D1BWP30P140LVT U12262 ( .A1(i_data_bus[391]), .A2(n10387), .B1(
        i_data_bus[487]), .B2(n10385), .ZN(n8403) );
  AOI22D1BWP30P140LVT U12263 ( .A1(i_data_bus[423]), .A2(n10386), .B1(
        i_data_bus[455]), .B2(n10388), .ZN(n8402) );
  ND2D1BWP30P140LVT U12264 ( .A1(n8403), .A2(n8402), .ZN(N10760) );
  AOI22D1BWP30P140LVT U12265 ( .A1(i_data_bus[413]), .A2(n10387), .B1(
        i_data_bus[509]), .B2(n10385), .ZN(n8405) );
  AOI22D1BWP30P140LVT U12266 ( .A1(i_data_bus[477]), .A2(n10388), .B1(
        i_data_bus[445]), .B2(n10386), .ZN(n8404) );
  ND2D1BWP30P140LVT U12267 ( .A1(n8405), .A2(n8404), .ZN(N10782) );
  AOI22D1BWP30P140LVT U12268 ( .A1(i_data_bus[400]), .A2(n10387), .B1(
        i_data_bus[496]), .B2(n10385), .ZN(n8407) );
  AOI22D1BWP30P140LVT U12269 ( .A1(i_data_bus[464]), .A2(n10388), .B1(
        i_data_bus[432]), .B2(n10386), .ZN(n8406) );
  ND2D1BWP30P140LVT U12270 ( .A1(n8407), .A2(n8406), .ZN(N10769) );
  AOI22D1BWP30P140LVT U12271 ( .A1(i_data_bus[395]), .A2(n10387), .B1(
        i_data_bus[491]), .B2(n10385), .ZN(n8409) );
  AOI22D1BWP30P140LVT U12272 ( .A1(i_data_bus[459]), .A2(n10388), .B1(
        i_data_bus[427]), .B2(n10386), .ZN(n8408) );
  ND2D1BWP30P140LVT U12273 ( .A1(n8409), .A2(n8408), .ZN(N10764) );
  AOI22D1BWP30P140LVT U12274 ( .A1(i_data_bus[388]), .A2(n10387), .B1(
        i_data_bus[484]), .B2(n10385), .ZN(n8411) );
  AOI22D1BWP30P140LVT U12275 ( .A1(i_data_bus[452]), .A2(n10388), .B1(
        i_data_bus[420]), .B2(n10386), .ZN(n8410) );
  ND2D1BWP30P140LVT U12276 ( .A1(n8411), .A2(n8410), .ZN(N10757) );
  AOI22D1BWP30P140LVT U12277 ( .A1(i_data_bus[600]), .A2(n10013), .B1(
        i_data_bus[632]), .B2(n10011), .ZN(n8413) );
  AOI22D1BWP30P140LVT U12278 ( .A1(i_data_bus[568]), .A2(n10012), .B1(
        i_data_bus[536]), .B2(n10006), .ZN(n8412) );
  ND2D1BWP30P140LVT U12279 ( .A1(n8413), .A2(n8412), .ZN(N2693) );
  AOI22D1BWP30P140LVT U12280 ( .A1(i_data_bus[547]), .A2(n10012), .B1(
        i_data_bus[611]), .B2(n10011), .ZN(n8415) );
  AOI22D1BWP30P140LVT U12281 ( .A1(i_data_bus[579]), .A2(n10013), .B1(
        i_data_bus[515]), .B2(n10006), .ZN(n8414) );
  ND2D1BWP30P140LVT U12282 ( .A1(n8415), .A2(n8414), .ZN(N2672) );
  AOI22D1BWP30P140LVT U12283 ( .A1(i_data_bus[553]), .A2(n10012), .B1(
        i_data_bus[617]), .B2(n10011), .ZN(n8417) );
  AOI22D1BWP30P140LVT U12284 ( .A1(i_data_bus[521]), .A2(n10006), .B1(
        i_data_bus[585]), .B2(n10013), .ZN(n8416) );
  ND2D1BWP30P140LVT U12285 ( .A1(n8417), .A2(n8416), .ZN(N2678) );
  AOI22D1BWP30P140LVT U12286 ( .A1(i_data_bus[403]), .A2(n10407), .B1(
        i_data_bus[499]), .B2(n10406), .ZN(n8423) );
  AOI22D1BWP30P140LVT U12287 ( .A1(i_data_bus[467]), .A2(n10408), .B1(
        i_data_bus[435]), .B2(n10405), .ZN(n8422) );
  ND2D1BWP30P140LVT U12288 ( .A1(n8423), .A2(n8422), .ZN(N9410) );
  AOI22D1BWP30P140LVT U12289 ( .A1(i_data_bus[407]), .A2(n10407), .B1(
        i_data_bus[439]), .B2(n10405), .ZN(n8425) );
  AOI22D1BWP30P140LVT U12290 ( .A1(i_data_bus[471]), .A2(n10408), .B1(
        i_data_bus[503]), .B2(n10406), .ZN(n8424) );
  ND2D1BWP30P140LVT U12291 ( .A1(n8425), .A2(n8424), .ZN(N9414) );
  AOI22D1BWP30P140LVT U12292 ( .A1(i_data_bus[399]), .A2(n10407), .B1(
        i_data_bus[431]), .B2(n10405), .ZN(n8427) );
  AOI22D1BWP30P140LVT U12293 ( .A1(i_data_bus[463]), .A2(n10408), .B1(
        i_data_bus[495]), .B2(n10406), .ZN(n8426) );
  ND2D1BWP30P140LVT U12294 ( .A1(n8427), .A2(n8426), .ZN(N9406) );
  AOI22D1BWP30P140LVT U12295 ( .A1(i_data_bus[395]), .A2(n10407), .B1(
        i_data_bus[427]), .B2(n10405), .ZN(n8429) );
  AOI22D1BWP30P140LVT U12296 ( .A1(i_data_bus[459]), .A2(n10408), .B1(
        i_data_bus[491]), .B2(n10406), .ZN(n8428) );
  ND2D1BWP30P140LVT U12297 ( .A1(n8429), .A2(n8428), .ZN(N9402) );
  AOI22D1BWP30P140LVT U12298 ( .A1(i_data_bus[391]), .A2(n10407), .B1(
        i_data_bus[423]), .B2(n10405), .ZN(n8431) );
  AOI22D1BWP30P140LVT U12299 ( .A1(i_data_bus[455]), .A2(n10408), .B1(
        i_data_bus[487]), .B2(n10406), .ZN(n8430) );
  ND2D1BWP30P140LVT U12300 ( .A1(n8431), .A2(n8430), .ZN(N9398) );
  AOI22D1BWP30P140LVT U12301 ( .A1(i_data_bus[413]), .A2(n10407), .B1(
        i_data_bus[445]), .B2(n10405), .ZN(n8433) );
  AOI22D1BWP30P140LVT U12302 ( .A1(i_data_bus[509]), .A2(n10406), .B1(
        i_data_bus[477]), .B2(n10408), .ZN(n8432) );
  ND2D1BWP30P140LVT U12303 ( .A1(n8433), .A2(n8432), .ZN(N9420) );
  AOI22D1BWP30P140LVT U12304 ( .A1(i_data_bus[404]), .A2(n10407), .B1(
        i_data_bus[436]), .B2(n10405), .ZN(n8435) );
  AOI22D1BWP30P140LVT U12305 ( .A1(i_data_bus[500]), .A2(n10406), .B1(
        i_data_bus[468]), .B2(n10408), .ZN(n8434) );
  ND2D1BWP30P140LVT U12306 ( .A1(n8435), .A2(n8434), .ZN(N9411) );
  AOI22D1BWP30P140LVT U12307 ( .A1(i_data_bus[401]), .A2(n10407), .B1(
        i_data_bus[465]), .B2(n10408), .ZN(n8437) );
  AOI22D1BWP30P140LVT U12308 ( .A1(i_data_bus[433]), .A2(n10405), .B1(
        i_data_bus[497]), .B2(n10406), .ZN(n8436) );
  ND2D1BWP30P140LVT U12309 ( .A1(n8437), .A2(n8436), .ZN(N9408) );
  AOI22D1BWP30P140LVT U12310 ( .A1(i_data_bus[400]), .A2(n10407), .B1(
        i_data_bus[464]), .B2(n10408), .ZN(n8439) );
  AOI22D1BWP30P140LVT U12311 ( .A1(i_data_bus[496]), .A2(n10406), .B1(
        i_data_bus[432]), .B2(n10405), .ZN(n8438) );
  ND2D1BWP30P140LVT U12312 ( .A1(n8439), .A2(n8438), .ZN(N9407) );
  AOI22D1BWP30P140LVT U12313 ( .A1(i_data_bus[414]), .A2(n10429), .B1(
        i_data_bus[478]), .B2(n10430), .ZN(n8449) );
  AOI22D1BWP30P140LVT U12314 ( .A1(i_data_bus[446]), .A2(n10427), .B1(
        i_data_bus[510]), .B2(n10428), .ZN(n8448) );
  ND2D1BWP30P140LVT U12315 ( .A1(n8449), .A2(n8448), .ZN(N6697) );
  AOI22D1BWP30P140LVT U12316 ( .A1(i_data_bus[394]), .A2(n10429), .B1(
        i_data_bus[458]), .B2(n10430), .ZN(n8451) );
  AOI22D1BWP30P140LVT U12317 ( .A1(i_data_bus[426]), .A2(n10427), .B1(
        i_data_bus[490]), .B2(n10428), .ZN(n8450) );
  ND2D1BWP30P140LVT U12318 ( .A1(n8451), .A2(n8450), .ZN(N6677) );
  AOI22D1BWP30P140LVT U12319 ( .A1(i_data_bus[404]), .A2(n10429), .B1(
        i_data_bus[436]), .B2(n10427), .ZN(n8453) );
  AOI22D1BWP30P140LVT U12320 ( .A1(i_data_bus[500]), .A2(n10428), .B1(
        i_data_bus[468]), .B2(n10430), .ZN(n8452) );
  ND2D1BWP30P140LVT U12321 ( .A1(n8453), .A2(n8452), .ZN(N6687) );
  AOI22D1BWP30P140LVT U12322 ( .A1(i_data_bus[398]), .A2(n10429), .B1(
        i_data_bus[494]), .B2(n10428), .ZN(n8455) );
  AOI22D1BWP30P140LVT U12323 ( .A1(i_data_bus[430]), .A2(n10427), .B1(
        i_data_bus[462]), .B2(n10430), .ZN(n8454) );
  ND2D1BWP30P140LVT U12324 ( .A1(n8455), .A2(n8454), .ZN(N6681) );
  AOI22D1BWP30P140LVT U12325 ( .A1(i_data_bus[407]), .A2(n10429), .B1(
        i_data_bus[439]), .B2(n10427), .ZN(n8457) );
  AOI22D1BWP30P140LVT U12326 ( .A1(i_data_bus[471]), .A2(n10430), .B1(
        i_data_bus[503]), .B2(n10428), .ZN(n8456) );
  ND2D1BWP30P140LVT U12327 ( .A1(n8457), .A2(n8456), .ZN(N6690) );
  AOI22D1BWP30P140LVT U12328 ( .A1(i_data_bus[403]), .A2(n10429), .B1(
        i_data_bus[435]), .B2(n10427), .ZN(n8459) );
  AOI22D1BWP30P140LVT U12329 ( .A1(i_data_bus[467]), .A2(n10430), .B1(
        i_data_bus[499]), .B2(n10428), .ZN(n8458) );
  ND2D1BWP30P140LVT U12330 ( .A1(n8459), .A2(n8458), .ZN(N6686) );
  AOI22D1BWP30P140LVT U12331 ( .A1(i_data_bus[401]), .A2(n10429), .B1(
        i_data_bus[497]), .B2(n10428), .ZN(n8461) );
  AOI22D1BWP30P140LVT U12332 ( .A1(i_data_bus[465]), .A2(n10430), .B1(
        i_data_bus[433]), .B2(n10427), .ZN(n8460) );
  ND2D1BWP30P140LVT U12333 ( .A1(n8461), .A2(n8460), .ZN(N6684) );
  AOI22D1BWP30P140LVT U12334 ( .A1(i_data_bus[397]), .A2(n10429), .B1(
        i_data_bus[493]), .B2(n10428), .ZN(n8463) );
  AOI22D1BWP30P140LVT U12335 ( .A1(i_data_bus[461]), .A2(n10430), .B1(
        i_data_bus[429]), .B2(n10427), .ZN(n8462) );
  ND2D1BWP30P140LVT U12336 ( .A1(n8463), .A2(n8462), .ZN(N6680) );
  AOI22D1BWP30P140LVT U12337 ( .A1(i_data_bus[395]), .A2(n10429), .B1(
        i_data_bus[491]), .B2(n10428), .ZN(n8465) );
  AOI22D1BWP30P140LVT U12338 ( .A1(i_data_bus[459]), .A2(n10430), .B1(
        i_data_bus[427]), .B2(n10427), .ZN(n8464) );
  ND2D1BWP30P140LVT U12339 ( .A1(n8465), .A2(n8464), .ZN(N6678) );
  AOI22D1BWP30P140LVT U12340 ( .A1(i_data_bus[571]), .A2(n10271), .B1(
        i_data_bus[635]), .B2(n10270), .ZN(n8467) );
  AOI22D1BWP30P140LVT U12341 ( .A1(i_data_bus[603]), .A2(n10269), .B1(
        i_data_bus[539]), .B2(n10272), .ZN(n8466) );
  ND2D1BWP30P140LVT U12342 ( .A1(n8467), .A2(n8466), .ZN(N8144) );
  AOI22D1BWP30P140LVT U12343 ( .A1(i_data_bus[600]), .A2(n10269), .B1(
        i_data_bus[632]), .B2(n10270), .ZN(n8469) );
  AOI22D1BWP30P140LVT U12344 ( .A1(i_data_bus[568]), .A2(n10271), .B1(
        i_data_bus[536]), .B2(n10272), .ZN(n8468) );
  ND2D1BWP30P140LVT U12345 ( .A1(n8469), .A2(n8468), .ZN(N8141) );
  AOI22D1BWP30P140LVT U12346 ( .A1(i_data_bus[540]), .A2(n10272), .B1(
        i_data_bus[636]), .B2(n10270), .ZN(n8471) );
  AOI22D1BWP30P140LVT U12347 ( .A1(i_data_bus[572]), .A2(n10271), .B1(
        i_data_bus[604]), .B2(n10269), .ZN(n8470) );
  ND2D1BWP30P140LVT U12348 ( .A1(n8471), .A2(n8470), .ZN(N8145) );
  INR4D1BWP30P140LVT U12349 ( .A1(i_cmd[86]), .B1(i_cmd[70]), .B2(n10395), 
        .B3(n10957), .ZN(n10275) );
  NR4D1BWP30P140LVT U12350 ( .A1(i_cmd[78]), .A2(n10392), .A3(n10959), .A4(
        n8472), .ZN(n10277) );
  AOI22D1BWP30P140LVT U12351 ( .A1(i_data_bus[349]), .A2(n10275), .B1(
        i_data_bus[381]), .B2(n10277), .ZN(n8474) );
  NR4D1BWP30P140LVT U12352 ( .A1(i_cmd[94]), .A2(n10960), .A3(n10391), .A4(
        n8472), .ZN(n10276) );
  NR3D0P7BWP30P140LVT U12353 ( .A1(i_cmd[78]), .A2(i_cmd[94]), .A3(i_cmd[86]), 
        .ZN(n10956) );
  AOI22D1BWP30P140LVT U12354 ( .A1(i_data_bus[317]), .A2(n10276), .B1(
        i_data_bus[285]), .B2(n6227), .ZN(n8473) );
  ND2D1BWP30P140LVT U12355 ( .A1(n8474), .A2(n8473), .ZN(N9204) );
  AOI22D1BWP30P140LVT U12356 ( .A1(i_data_bus[335]), .A2(n10275), .B1(
        i_data_bus[367]), .B2(n10277), .ZN(n8476) );
  AOI22D1BWP30P140LVT U12357 ( .A1(i_data_bus[303]), .A2(n10276), .B1(
        i_data_bus[271]), .B2(n6227), .ZN(n8475) );
  ND2D1BWP30P140LVT U12358 ( .A1(n8476), .A2(n8475), .ZN(N9190) );
  AOI22D1BWP30P140LVT U12359 ( .A1(i_data_bus[322]), .A2(n10275), .B1(
        i_data_bus[354]), .B2(n10277), .ZN(n8478) );
  AOI22D1BWP30P140LVT U12360 ( .A1(i_data_bus[290]), .A2(n10276), .B1(
        i_data_bus[258]), .B2(n6227), .ZN(n8477) );
  ND2D1BWP30P140LVT U12361 ( .A1(n8478), .A2(n8477), .ZN(N9177) );
  INR4D1BWP30P140LVT U12362 ( .A1(i_cmd[87]), .B1(i_cmd[71]), .B2(n10395), 
        .B3(n10928), .ZN(n9879) );
  NR4D1BWP30P140LVT U12363 ( .A1(i_cmd[79]), .A2(n10392), .A3(n10930), .A4(
        n8479), .ZN(n9877) );
  AOI22D1BWP30P140LVT U12364 ( .A1(i_data_bus[321]), .A2(n9879), .B1(
        i_data_bus[353]), .B2(n9877), .ZN(n8481) );
  NR4D1BWP30P140LVT U12365 ( .A1(i_cmd[95]), .A2(n10931), .A3(n10391), .A4(
        n8479), .ZN(n9878) );
  NR3D0P7BWP30P140LVT U12366 ( .A1(i_cmd[87]), .A2(i_cmd[79]), .A3(i_cmd[95]), 
        .ZN(n10927) );
  AOI22D1BWP30P140LVT U12367 ( .A1(i_data_bus[289]), .A2(n9878), .B1(
        i_data_bus[257]), .B2(n6217), .ZN(n8480) );
  ND2D1BWP30P140LVT U12368 ( .A1(n8481), .A2(n8480), .ZN(N10666) );
  AOI22D1BWP30P140LVT U12369 ( .A1(i_data_bus[319]), .A2(n9878), .B1(
        i_data_bus[383]), .B2(n9877), .ZN(n8483) );
  AOI22D1BWP30P140LVT U12370 ( .A1(i_data_bus[351]), .A2(n9879), .B1(
        i_data_bus[287]), .B2(n6217), .ZN(n8482) );
  ND2D1BWP30P140LVT U12371 ( .A1(n8483), .A2(n8482), .ZN(N10696) );
  AOI22D1BWP30P140LVT U12372 ( .A1(i_data_bus[290]), .A2(n9878), .B1(
        i_data_bus[354]), .B2(n9877), .ZN(n8485) );
  AOI22D1BWP30P140LVT U12373 ( .A1(i_data_bus[322]), .A2(n9879), .B1(
        i_data_bus[258]), .B2(n6217), .ZN(n8484) );
  ND2D1BWP30P140LVT U12374 ( .A1(n8485), .A2(n8484), .ZN(N10667) );
  INR4D1BWP30P140LVT U12375 ( .A1(i_cmd[22]), .B1(i_cmd[6]), .B2(n10632), .B3(
        n10967), .ZN(n9790) );
  NR4D1BWP30P140LVT U12376 ( .A1(i_cmd[30]), .A2(n10634), .A3(n8486), .A4(
        n8487), .ZN(n9791) );
  AOI22D1BWP30P140LVT U12377 ( .A1(i_data_bus[74]), .A2(n9790), .B1(
        i_data_bus[42]), .B2(n9791), .ZN(n8490) );
  NR4D1BWP30P140LVT U12378 ( .A1(i_cmd[14]), .A2(n8488), .A3(n10630), .A4(
        n8487), .ZN(n9792) );
  NR3D0P7BWP30P140LVT U12379 ( .A1(i_cmd[22]), .A2(i_cmd[30]), .A3(i_cmd[14]), 
        .ZN(n10963) );
  AOI22D1BWP30P140LVT U12380 ( .A1(i_data_bus[106]), .A2(n9792), .B1(
        i_data_bus[10]), .B2(n6223), .ZN(n8489) );
  ND2D1BWP30P140LVT U12381 ( .A1(n8490), .A2(n8489), .ZN(N8753) );
  INR4D1BWP30P140LVT U12382 ( .A1(i_cmd[21]), .B1(i_cmd[5]), .B2(n10632), .B3(
        n11013), .ZN(n10115) );
  NR4D1BWP30P140LVT U12383 ( .A1(i_cmd[29]), .A2(n10634), .A3(n8491), .A4(
        n8492), .ZN(n10118) );
  AOI22D1BWP30P140LVT U12384 ( .A1(i_data_bus[76]), .A2(n10115), .B1(
        i_data_bus[44]), .B2(n10118), .ZN(n8495) );
  NR4D1BWP30P140LVT U12385 ( .A1(i_cmd[13]), .A2(n8493), .A3(n10630), .A4(
        n8492), .ZN(n10117) );
  NR3D0P7BWP30P140LVT U12386 ( .A1(i_cmd[21]), .A2(i_cmd[29]), .A3(i_cmd[13]), 
        .ZN(n11009) );
  AOI22D1BWP30P140LVT U12387 ( .A1(i_data_bus[108]), .A2(n10117), .B1(
        i_data_bus[12]), .B2(n10116), .ZN(n8494) );
  ND2D1BWP30P140LVT U12388 ( .A1(n8495), .A2(n8494), .ZN(N7777) );
  INR4D1BWP30P140LVT U12389 ( .A1(i_cmd[83]), .B1(i_cmd[67]), .B2(n10395), 
        .B3(n11083), .ZN(n9755) );
  NR4D1BWP30P140LVT U12390 ( .A1(i_cmd[91]), .A2(n10391), .A3(n11085), .A4(
        n8496), .ZN(n9758) );
  AOI22D1BWP30P140LVT U12391 ( .A1(i_data_bus[340]), .A2(n9755), .B1(
        i_data_bus[308]), .B2(n9758), .ZN(n8498) );
  NR4D1BWP30P140LVT U12392 ( .A1(i_cmd[75]), .A2(n11086), .A3(n10392), .A4(
        n8496), .ZN(n9757) );
  NR3D0P7BWP30P140LVT U12393 ( .A1(i_cmd[83]), .A2(i_cmd[91]), .A3(i_cmd[75]), 
        .ZN(n11082) );
  AOI22D1BWP30P140LVT U12394 ( .A1(i_data_bus[372]), .A2(n9757), .B1(
        i_data_bus[276]), .B2(n9756), .ZN(n8497) );
  ND2D1BWP30P140LVT U12395 ( .A1(n8498), .A2(n8497), .ZN(N5237) );
  AOI22D1BWP30P140LVT U12396 ( .A1(i_data_bus[118]), .A2(n10117), .B1(
        i_data_bus[54]), .B2(n10118), .ZN(n8500) );
  AOI22D1BWP30P140LVT U12397 ( .A1(i_data_bus[86]), .A2(n10115), .B1(
        i_data_bus[22]), .B2(n10116), .ZN(n8499) );
  ND2D1BWP30P140LVT U12398 ( .A1(n8500), .A2(n8499), .ZN(N7787) );
  INR4D1BWP30P140LVT U12399 ( .A1(i_cmd[18]), .B1(i_cmd[2]), .B2(n10632), .B3(
        n8501), .ZN(n9914) );
  NR4D1BWP30P140LVT U12400 ( .A1(i_cmd[10]), .A2(n10630), .A3(n8502), .A4(
        n8503), .ZN(n9915) );
  AOI22D1BWP30P140LVT U12401 ( .A1(i_data_bus[87]), .A2(n9914), .B1(
        i_data_bus[119]), .B2(n9915), .ZN(n8507) );
  NR4D1BWP30P140LVT U12402 ( .A1(i_cmd[26]), .A2(n8504), .A3(n10634), .A4(
        n8503), .ZN(n9916) );
  AOI22D1BWP30P140LVT U12403 ( .A1(i_data_bus[55]), .A2(n9916), .B1(
        i_data_bus[23]), .B2(n6218), .ZN(n8506) );
  ND2D1BWP30P140LVT U12404 ( .A1(n8507), .A2(n8506), .ZN(N3318) );
  AOI22D1BWP30P140LVT U12405 ( .A1(i_data_bus[118]), .A2(n9792), .B1(
        i_data_bus[54]), .B2(n9791), .ZN(n8509) );
  AOI22D1BWP30P140LVT U12406 ( .A1(i_data_bus[86]), .A2(n9790), .B1(
        i_data_bus[22]), .B2(n6223), .ZN(n8508) );
  ND2D1BWP30P140LVT U12407 ( .A1(n8509), .A2(n8508), .ZN(N8765) );
  AOI22D1BWP30P140LVT U12408 ( .A1(i_data_bus[378]), .A2(n9757), .B1(
        i_data_bus[314]), .B2(n9758), .ZN(n8511) );
  AOI22D1BWP30P140LVT U12409 ( .A1(i_data_bus[346]), .A2(n9755), .B1(
        i_data_bus[282]), .B2(n9756), .ZN(n8510) );
  ND2D1BWP30P140LVT U12410 ( .A1(n8511), .A2(n8510), .ZN(N5243) );
  AOI22D1BWP30P140LVT U12411 ( .A1(i_data_bus[61]), .A2(n9916), .B1(
        i_data_bus[125]), .B2(n9915), .ZN(n8513) );
  AOI22D1BWP30P140LVT U12412 ( .A1(i_data_bus[93]), .A2(n9914), .B1(
        i_data_bus[29]), .B2(n6218), .ZN(n8512) );
  ND2D1BWP30P140LVT U12413 ( .A1(n8513), .A2(n8512), .ZN(N3324) );
  AOI22D1BWP30P140LVT U12414 ( .A1(i_data_bus[60]), .A2(n9916), .B1(
        i_data_bus[124]), .B2(n9915), .ZN(n8515) );
  AOI22D1BWP30P140LVT U12415 ( .A1(i_data_bus[92]), .A2(n9914), .B1(
        i_data_bus[28]), .B2(n6218), .ZN(n8514) );
  ND2D1BWP30P140LVT U12416 ( .A1(n8515), .A2(n8514), .ZN(N3323) );
  AOI22D1BWP30P140LVT U12417 ( .A1(i_data_bus[205]), .A2(n10218), .B1(
        i_data_bus[141]), .B2(n6213), .ZN(n8517) );
  AOI22D1BWP30P140LVT U12418 ( .A1(i_data_bus[173]), .A2(n10219), .B1(
        i_data_bus[237]), .B2(n10220), .ZN(n8516) );
  ND2D1BWP30P140LVT U12419 ( .A1(n8517), .A2(n8516), .ZN(N2418) );
  AOI22D1BWP30P140LVT U12420 ( .A1(i_data_bus[230]), .A2(n10131), .B1(
        i_data_bus[198]), .B2(n10132), .ZN(n8519) );
  AOI22D1BWP30P140LVT U12421 ( .A1(i_data_bus[166]), .A2(n10133), .B1(
        i_data_bus[134]), .B2(n10134), .ZN(n8518) );
  ND2D1BWP30P140LVT U12422 ( .A1(n8519), .A2(n8518), .ZN(N7859) );
  AOI22D1BWP30P140LVT U12423 ( .A1(i_data_bus[160]), .A2(n10225), .B1(
        i_data_bus[192]), .B2(n10223), .ZN(n8521) );
  AOI22D1BWP30P140LVT U12424 ( .A1(i_data_bus[224]), .A2(n10226), .B1(
        i_data_bus[128]), .B2(n10224), .ZN(n8520) );
  ND2D1BWP30P140LVT U12425 ( .A1(n8521), .A2(n8520), .ZN(N6235) );
  INR4D1BWP30P140LVT U12426 ( .A1(i_cmd[85]), .B1(i_cmd[69]), .B2(n10395), 
        .B3(n10998), .ZN(n9844) );
  NR4D1BWP30P140LVT U12427 ( .A1(i_cmd[93]), .A2(n10391), .A3(n11000), .A4(
        n8522), .ZN(n9843) );
  AOI22D1BWP30P140LVT U12428 ( .A1(i_data_bus[328]), .A2(n9844), .B1(
        i_data_bus[296]), .B2(n9843), .ZN(n8524) );
  NR4D1BWP30P140LVT U12429 ( .A1(i_cmd[77]), .A2(n11001), .A3(n10392), .A4(
        n8522), .ZN(n9845) );
  NR3D0P7BWP30P140LVT U12430 ( .A1(i_cmd[85]), .A2(i_cmd[93]), .A3(i_cmd[77]), 
        .ZN(n10997) );
  AOI22D1BWP30P140LVT U12431 ( .A1(i_data_bus[360]), .A2(n9845), .B1(
        i_data_bus[264]), .B2(n9846), .ZN(n8523) );
  ND2D1BWP30P140LVT U12432 ( .A1(n8524), .A2(n8523), .ZN(N7949) );
  INR4D1BWP30P140LVT U12433 ( .A1(i_cmd[81]), .B1(i_cmd[65]), .B2(n10395), 
        .B3(n11136), .ZN(n9774) );
  NR4D1BWP30P140LVT U12434 ( .A1(i_cmd[73]), .A2(n10392), .A3(n8525), .A4(
        n8526), .ZN(n9773) );
  AOI22D1BWP30P140LVT U12435 ( .A1(i_data_bus[351]), .A2(n9774), .B1(
        i_data_bus[383]), .B2(n9773), .ZN(n8529) );
  NR4D1BWP30P140LVT U12436 ( .A1(i_cmd[89]), .A2(n8527), .A3(n10391), .A4(
        n8526), .ZN(n9775) );
  NR3D0P7BWP30P140LVT U12437 ( .A1(i_cmd[81]), .A2(i_cmd[73]), .A3(i_cmd[89]), 
        .ZN(n11132) );
  ND2D1BWP30P140LVT U12438 ( .A1(n11132), .A2(i_cmd[65]), .ZN(n11134) );
  AOI22D1BWP30P140LVT U12439 ( .A1(i_data_bus[319]), .A2(n9775), .B1(
        i_data_bus[287]), .B2(n6216), .ZN(n8528) );
  ND2D1BWP30P140LVT U12440 ( .A1(n8529), .A2(n8528), .ZN(N2524) );
  AOI22D1BWP30P140LVT U12441 ( .A1(i_data_bus[349]), .A2(n9774), .B1(
        i_data_bus[381]), .B2(n9773), .ZN(n8531) );
  AOI22D1BWP30P140LVT U12442 ( .A1(i_data_bus[317]), .A2(n9775), .B1(
        i_data_bus[285]), .B2(n6216), .ZN(n8530) );
  ND2D1BWP30P140LVT U12443 ( .A1(n8531), .A2(n8530), .ZN(N2522) );
  AOI22D1BWP30P140LVT U12444 ( .A1(i_data_bus[369]), .A2(n9845), .B1(
        i_data_bus[305]), .B2(n9843), .ZN(n8533) );
  AOI22D1BWP30P140LVT U12445 ( .A1(i_data_bus[337]), .A2(n9844), .B1(
        i_data_bus[273]), .B2(n9846), .ZN(n8532) );
  ND2D1BWP30P140LVT U12446 ( .A1(n8533), .A2(n8532), .ZN(N7958) );
  INR4D1BWP30P140LVT U12447 ( .A1(i_cmd[51]), .B1(i_cmd[35]), .B2(n10667), 
        .B3(n11090), .ZN(n9521) );
  NR4D1BWP30P140LVT U12448 ( .A1(i_cmd[59]), .A2(n10664), .A3(n11092), .A4(
        n8534), .ZN(n9519) );
  AOI22D1BWP30P140LVT U12449 ( .A1(i_data_bus[199]), .A2(n9521), .B1(
        i_data_bus[167]), .B2(n9519), .ZN(n8536) );
  NR4D1BWP30P140LVT U12450 ( .A1(i_cmd[43]), .A2(n11093), .A3(n10670), .A4(
        n8534), .ZN(n9520) );
  NR3D0P7BWP30P140LVT U12451 ( .A1(i_cmd[51]), .A2(i_cmd[59]), .A3(i_cmd[43]), 
        .ZN(n11089) );
  AOI22D1BWP30P140LVT U12452 ( .A1(i_data_bus[231]), .A2(n9520), .B1(
        i_data_bus[135]), .B2(n9522), .ZN(n8535) );
  ND2D1BWP30P140LVT U12453 ( .A1(n8536), .A2(n8535), .ZN(N5136) );
  NR4D1BWP30P140LVT U12454 ( .A1(i_cmd[27]), .A2(n8537), .A3(n10634), .A4(
        n8538), .ZN(n10087) );
  NR4D1BWP30P140LVT U12455 ( .A1(i_cmd[11]), .A2(n10630), .A3(n8539), .A4(
        n8538), .ZN(n10085) );
  AOI22D1BWP30P140LVT U12456 ( .A1(i_data_bus[41]), .A2(n10087), .B1(
        i_data_bus[105]), .B2(n10085), .ZN(n8543) );
  INR4D1BWP30P140LVT U12457 ( .A1(i_cmd[19]), .B1(i_cmd[3]), .B2(n10632), .B3(
        n8540), .ZN(n10086) );
  AOI22D1BWP30P140LVT U12458 ( .A1(i_data_bus[73]), .A2(n10086), .B1(
        i_data_bus[9]), .B2(n10088), .ZN(n8542) );
  ND2D1BWP30P140LVT U12459 ( .A1(n8543), .A2(n8542), .ZN(N5050) );
  AOI22D1BWP30P140LVT U12460 ( .A1(i_data_bus[249]), .A2(n9520), .B1(
        i_data_bus[185]), .B2(n9519), .ZN(n8545) );
  AOI22D1BWP30P140LVT U12461 ( .A1(i_data_bus[217]), .A2(n9521), .B1(
        i_data_bus[153]), .B2(n9522), .ZN(n8544) );
  ND2D1BWP30P140LVT U12462 ( .A1(n8545), .A2(n8544), .ZN(N5154) );
  AOI22D1BWP30P140LVT U12463 ( .A1(i_data_bus[244]), .A2(n9520), .B1(
        i_data_bus[180]), .B2(n9519), .ZN(n8547) );
  AOI22D1BWP30P140LVT U12464 ( .A1(i_data_bus[212]), .A2(n9521), .B1(
        i_data_bus[148]), .B2(n9522), .ZN(n8546) );
  ND2D1BWP30P140LVT U12465 ( .A1(n8547), .A2(n8546), .ZN(N5149) );
  AOI22D1BWP30P140LVT U12466 ( .A1(i_data_bus[229]), .A2(n9520), .B1(
        i_data_bus[165]), .B2(n9519), .ZN(n8549) );
  AOI22D1BWP30P140LVT U12467 ( .A1(i_data_bus[197]), .A2(n9521), .B1(
        i_data_bus[133]), .B2(n9522), .ZN(n8548) );
  ND2D1BWP30P140LVT U12468 ( .A1(n8549), .A2(n8548), .ZN(N5134) );
  AOI22D1BWP30P140LVT U12469 ( .A1(i_data_bus[222]), .A2(n9521), .B1(
        i_data_bus[254]), .B2(n9520), .ZN(n8551) );
  AOI22D1BWP30P140LVT U12470 ( .A1(i_data_bus[190]), .A2(n9519), .B1(
        i_data_bus[158]), .B2(n9522), .ZN(n8550) );
  ND2D1BWP30P140LVT U12471 ( .A1(n8551), .A2(n8550), .ZN(N5159) );
  AOI22D1BWP30P140LVT U12472 ( .A1(i_data_bus[373]), .A2(n9773), .B1(
        i_data_bus[341]), .B2(n9774), .ZN(n8553) );
  AOI22D1BWP30P140LVT U12473 ( .A1(i_data_bus[309]), .A2(n9775), .B1(
        i_data_bus[277]), .B2(n6216), .ZN(n8552) );
  ND2D1BWP30P140LVT U12474 ( .A1(n8553), .A2(n8552), .ZN(N2514) );
  AOI22D1BWP30P140LVT U12475 ( .A1(i_data_bus[224]), .A2(n10038), .B1(
        i_data_bus[192]), .B2(n10039), .ZN(n8555) );
  AOI22D1BWP30P140LVT U12476 ( .A1(i_data_bus[160]), .A2(n10040), .B1(
        i_data_bus[128]), .B2(n9318), .ZN(n8554) );
  ND2D1BWP30P140LVT U12477 ( .A1(n8555), .A2(n8554), .ZN(N8959) );
  AOI22D1BWP30P140LVT U12478 ( .A1(i_data_bus[162]), .A2(n10040), .B1(
        i_data_bus[194]), .B2(n10039), .ZN(n8557) );
  AOI22D1BWP30P140LVT U12479 ( .A1(i_data_bus[226]), .A2(n10038), .B1(
        i_data_bus[130]), .B2(n9318), .ZN(n8556) );
  ND2D1BWP30P140LVT U12480 ( .A1(n8557), .A2(n8556), .ZN(N8961) );
  AOI22D1BWP30P140LVT U12481 ( .A1(i_data_bus[161]), .A2(n10040), .B1(
        i_data_bus[193]), .B2(n10039), .ZN(n8559) );
  AOI22D1BWP30P140LVT U12482 ( .A1(i_data_bus[225]), .A2(n10038), .B1(
        i_data_bus[129]), .B2(n9318), .ZN(n8558) );
  ND2D1BWP30P140LVT U12483 ( .A1(n8559), .A2(n8558), .ZN(N8960) );
  AOI22D1BWP30P140LVT U12484 ( .A1(i_data_bus[312]), .A2(n9775), .B1(
        i_data_bus[344]), .B2(n9774), .ZN(n8561) );
  AOI22D1BWP30P140LVT U12485 ( .A1(i_data_bus[376]), .A2(n9773), .B1(
        i_data_bus[280]), .B2(n6216), .ZN(n8560) );
  ND2D1BWP30P140LVT U12486 ( .A1(n8561), .A2(n8560), .ZN(N2517) );
  AOI22D1BWP30P140LVT U12487 ( .A1(i_data_bus[301]), .A2(n9775), .B1(
        i_data_bus[333]), .B2(n9774), .ZN(n8563) );
  AOI22D1BWP30P140LVT U12488 ( .A1(i_data_bus[365]), .A2(n9773), .B1(
        i_data_bus[269]), .B2(n6216), .ZN(n8562) );
  ND2D1BWP30P140LVT U12489 ( .A1(n8563), .A2(n8562), .ZN(N2506) );
  AOI22D1BWP30P140LVT U12490 ( .A1(i_data_bus[297]), .A2(n9775), .B1(
        i_data_bus[329]), .B2(n9774), .ZN(n8565) );
  AOI22D1BWP30P140LVT U12491 ( .A1(i_data_bus[361]), .A2(n9773), .B1(
        i_data_bus[265]), .B2(n6216), .ZN(n8564) );
  ND2D1BWP30P140LVT U12492 ( .A1(n8565), .A2(n8564), .ZN(N2502) );
  NR4D1BWP30P140LVT U12493 ( .A1(i_cmd[90]), .A2(n8566), .A3(n10391), .A4(
        n8567), .ZN(n9732) );
  NR4D1BWP30P140LVT U12494 ( .A1(i_cmd[74]), .A2(n10392), .A3(n8568), .A4(
        n8567), .ZN(n9730) );
  AOI22D1BWP30P140LVT U12495 ( .A1(i_data_bus[319]), .A2(n9732), .B1(
        i_data_bus[383]), .B2(n9730), .ZN(n8572) );
  INR4D1BWP30P140LVT U12496 ( .A1(i_cmd[82]), .B1(i_cmd[66]), .B2(n10395), 
        .B3(n8569), .ZN(n9731) );
  AOI22D1BWP30P140LVT U12497 ( .A1(i_data_bus[351]), .A2(n9731), .B1(
        i_data_bus[287]), .B2(n6219), .ZN(n8571) );
  ND2D1BWP30P140LVT U12498 ( .A1(n8572), .A2(n8571), .ZN(N3758) );
  AOI22D1BWP30P140LVT U12499 ( .A1(i_data_bus[214]), .A2(n10223), .B1(
        i_data_bus[150]), .B2(n10224), .ZN(n8574) );
  AOI22D1BWP30P140LVT U12500 ( .A1(i_data_bus[182]), .A2(n10225), .B1(
        i_data_bus[246]), .B2(n10226), .ZN(n8573) );
  ND2D1BWP30P140LVT U12501 ( .A1(n8574), .A2(n8573), .ZN(N6257) );
  AOI22D1BWP30P140LVT U12502 ( .A1(i_data_bus[139]), .A2(n10224), .B1(
        i_data_bus[203]), .B2(n10223), .ZN(n8576) );
  AOI22D1BWP30P140LVT U12503 ( .A1(i_data_bus[171]), .A2(n10225), .B1(
        i_data_bus[235]), .B2(n10226), .ZN(n8575) );
  ND2D1BWP30P140LVT U12504 ( .A1(n8576), .A2(n8575), .ZN(N6246) );
  AOI22D1BWP30P140LVT U12505 ( .A1(i_data_bus[169]), .A2(n10225), .B1(
        i_data_bus[201]), .B2(n10223), .ZN(n8578) );
  AOI22D1BWP30P140LVT U12506 ( .A1(i_data_bus[137]), .A2(n10224), .B1(
        i_data_bus[233]), .B2(n10226), .ZN(n8577) );
  ND2D1BWP30P140LVT U12507 ( .A1(n8578), .A2(n8577), .ZN(N6244) );
  NR3D0P7BWP30P140LVT U12508 ( .A1(inner_first_stage_valid_reg[6]), .A2(
        inner_first_stage_valid_reg[7]), .A3(n11173), .ZN(n8579) );
  NR3D0P7BWP30P140LVT U12509 ( .A1(inner_first_stage_valid_reg[1]), .A2(
        inner_first_stage_valid_reg[5]), .A3(inner_first_stage_valid_reg[3]), 
        .ZN(n8584) );
  INR3D0BWP30P140LVT U12510 ( .A1(n8584), .B1(inner_first_stage_valid_reg[2]), 
        .B2(inner_first_stage_valid_reg[0]), .ZN(n8588) );
  INR4D1BWP30P140LVT U12511 ( .A1(inner_first_stage_valid_reg[3]), .B1(
        inner_first_stage_valid_reg[1]), .B2(inner_first_stage_valid_reg[5]), 
        .B3(n8583), .ZN(n11342) );
  INVD1BWP30P140LVT U12512 ( .I(inner_first_stage_valid_reg[6]), .ZN(n8582) );
  OR2D1BWP30P140LVT U12513 ( .A1(inner_first_stage_valid_reg[7]), .A2(n11173), 
        .Z(n8581) );
  INR4D1BWP30P140LVT U12514 ( .A1(n8588), .B1(n8582), .B2(
        inner_first_stage_valid_reg[4]), .B3(n8581), .ZN(n11341) );
  NR4D0BWP30P140LVT U12515 ( .A1(n11340), .A2(n11339), .A3(n11342), .A4(n11341), .ZN(n8590) );
  INR3D2BWP30P140LVT U12516 ( .A1(inner_first_stage_valid_reg[5]), .B1(
        inner_first_stage_valid_reg[1]), .B2(n8586), .ZN(n11351) );
  NR3D0P7BWP30P140LVT U12517 ( .A1(inner_first_stage_valid_reg[6]), .A2(
        inner_first_stage_valid_reg[4]), .A3(n11173), .ZN(n8587) );
  ND3D1BWP30P140LVT U12518 ( .A1(inner_first_stage_valid_reg[0]), .A2(n8584), 
        .A3(n8587), .ZN(n8585) );
  INR3D2BWP30P140LVT U12519 ( .A1(inner_first_stage_valid_reg[1]), .B1(
        inner_first_stage_valid_reg[5]), .B2(n8586), .ZN(n11344) );
  NR4D0BWP30P140LVT U12520 ( .A1(n11351), .A2(n11345), .A3(n11344), .A4(n11343), .ZN(n8589) );
  AOI22D1BWP30P140LVT U12521 ( .A1(i_data_bus[579]), .A2(n10183), .B1(
        i_data_bus[611]), .B2(n10185), .ZN(n8592) );
  AOI22D1BWP30P140LVT U12522 ( .A1(i_data_bus[547]), .A2(n10184), .B1(
        i_data_bus[515]), .B2(n10182), .ZN(n8591) );
  ND2D1BWP30P140LVT U12523 ( .A1(n8592), .A2(n8591), .ZN(N6886) );
  AOI22D1BWP30P140LVT U12524 ( .A1(i_data_bus[188]), .A2(n10219), .B1(
        i_data_bus[220]), .B2(n10218), .ZN(n8594) );
  AOI22D1BWP30P140LVT U12525 ( .A1(i_data_bus[252]), .A2(n10220), .B1(
        i_data_bus[156]), .B2(n6213), .ZN(n8593) );
  ND2D1BWP30P140LVT U12526 ( .A1(n8594), .A2(n8593), .ZN(N2433) );
  AOI22D1BWP30P140LVT U12527 ( .A1(i_data_bus[179]), .A2(n10219), .B1(
        i_data_bus[211]), .B2(n10218), .ZN(n8596) );
  AOI22D1BWP30P140LVT U12528 ( .A1(i_data_bus[243]), .A2(n10220), .B1(
        i_data_bus[147]), .B2(n6213), .ZN(n8595) );
  ND2D1BWP30P140LVT U12529 ( .A1(n8596), .A2(n8595), .ZN(N2424) );
  AOI22D1BWP30P140LVT U12530 ( .A1(i_data_bus[164]), .A2(n10219), .B1(
        i_data_bus[196]), .B2(n10218), .ZN(n8598) );
  AOI22D1BWP30P140LVT U12531 ( .A1(i_data_bus[228]), .A2(n10220), .B1(
        i_data_bus[132]), .B2(n6213), .ZN(n8597) );
  ND2D1BWP30P140LVT U12532 ( .A1(n8598), .A2(n8597), .ZN(N2409) );
  AOI22D1BWP30P140LVT U12533 ( .A1(i_data_bus[252]), .A2(n9520), .B1(
        i_data_bus[220]), .B2(n9521), .ZN(n8600) );
  AOI22D1BWP30P140LVT U12534 ( .A1(i_data_bus[188]), .A2(n9519), .B1(
        i_data_bus[156]), .B2(n9522), .ZN(n8599) );
  ND2D1BWP30P140LVT U12535 ( .A1(n8600), .A2(n8599), .ZN(N5157) );
  AOI22D1BWP30P140LVT U12536 ( .A1(i_data_bus[225]), .A2(n9520), .B1(
        i_data_bus[193]), .B2(n9521), .ZN(n8602) );
  AOI22D1BWP30P140LVT U12537 ( .A1(i_data_bus[161]), .A2(n9519), .B1(
        i_data_bus[129]), .B2(n9522), .ZN(n8601) );
  ND2D1BWP30P140LVT U12538 ( .A1(n8602), .A2(n8601), .ZN(N5130) );
  AOI22D1BWP30P140LVT U12539 ( .A1(i_data_bus[224]), .A2(n9520), .B1(
        i_data_bus[192]), .B2(n9521), .ZN(n8604) );
  AOI22D1BWP30P140LVT U12540 ( .A1(i_data_bus[160]), .A2(n9519), .B1(
        i_data_bus[128]), .B2(n9522), .ZN(n8603) );
  ND2D1BWP30P140LVT U12541 ( .A1(n8604), .A2(n8603), .ZN(N5129) );
  AOI22D1BWP30P140LVT U12542 ( .A1(i_data_bus[164]), .A2(n9519), .B1(
        i_data_bus[196]), .B2(n9521), .ZN(n8606) );
  AOI22D1BWP30P140LVT U12543 ( .A1(i_data_bus[228]), .A2(n9520), .B1(
        i_data_bus[132]), .B2(n9522), .ZN(n8605) );
  ND2D1BWP30P140LVT U12544 ( .A1(n8606), .A2(n8605), .ZN(N5133) );
  NR4D1BWP30P140LVT U12545 ( .A1(i_cmd[25]), .A2(n10634), .A3(n11147), .A4(
        n8607), .ZN(n9977) );
  INR4D1BWP30P140LVT U12546 ( .A1(i_cmd[17]), .B1(i_cmd[1]), .B2(n10632), .B3(
        n11145), .ZN(n9976) );
  AOI22D1BWP30P140LVT U12547 ( .A1(i_data_bus[36]), .A2(n9977), .B1(
        i_data_bus[68]), .B2(n9976), .ZN(n8609) );
  NR4D1BWP30P140LVT U12548 ( .A1(i_cmd[9]), .A2(n11148), .A3(n10630), .A4(
        n8607), .ZN(n9978) );
  NR3D0P7BWP30P140LVT U12549 ( .A1(i_cmd[17]), .A2(i_cmd[25]), .A3(i_cmd[9]), 
        .ZN(n11144) );
  AOI22D1BWP30P140LVT U12550 ( .A1(i_data_bus[100]), .A2(n9978), .B1(
        i_data_bus[4]), .B2(n9969), .ZN(n8608) );
  ND2D1BWP30P140LVT U12551 ( .A1(n8609), .A2(n8608), .ZN(N2321) );
  AOI22D1BWP30P140LVT U12552 ( .A1(i_data_bus[225]), .A2(n10220), .B1(
        i_data_bus[193]), .B2(n10218), .ZN(n8611) );
  AOI22D1BWP30P140LVT U12553 ( .A1(i_data_bus[161]), .A2(n10219), .B1(
        i_data_bus[129]), .B2(n6213), .ZN(n8610) );
  ND2D1BWP30P140LVT U12554 ( .A1(n8611), .A2(n8610), .ZN(N2406) );
  AOI22D1BWP30P140LVT U12555 ( .A1(i_data_bus[572]), .A2(n10184), .B1(
        i_data_bus[636]), .B2(n10185), .ZN(n8613) );
  AOI22D1BWP30P140LVT U12556 ( .A1(i_data_bus[604]), .A2(n10183), .B1(
        i_data_bus[540]), .B2(n10182), .ZN(n8612) );
  ND2D1BWP30P140LVT U12557 ( .A1(n8613), .A2(n8612), .ZN(N6911) );
  AOI22D1BWP30P140LVT U12558 ( .A1(i_data_bus[551]), .A2(n10184), .B1(
        i_data_bus[615]), .B2(n10185), .ZN(n8615) );
  AOI22D1BWP30P140LVT U12559 ( .A1(i_data_bus[583]), .A2(n10183), .B1(
        i_data_bus[519]), .B2(n10182), .ZN(n8614) );
  ND2D1BWP30P140LVT U12560 ( .A1(n8615), .A2(n8614), .ZN(N6890) );
  AOI22D1BWP30P140LVT U12561 ( .A1(i_data_bus[36]), .A2(n10087), .B1(
        i_data_bus[68]), .B2(n10086), .ZN(n8617) );
  AOI22D1BWP30P140LVT U12562 ( .A1(i_data_bus[100]), .A2(n10085), .B1(
        i_data_bus[4]), .B2(n10088), .ZN(n8616) );
  ND2D1BWP30P140LVT U12563 ( .A1(n8617), .A2(n8616), .ZN(N5045) );
  AOI22D1BWP30P140LVT U12564 ( .A1(i_data_bus[35]), .A2(n10087), .B1(
        i_data_bus[67]), .B2(n10086), .ZN(n8619) );
  AOI22D1BWP30P140LVT U12565 ( .A1(i_data_bus[99]), .A2(n10085), .B1(
        i_data_bus[3]), .B2(n10088), .ZN(n8618) );
  ND2D1BWP30P140LVT U12566 ( .A1(n8619), .A2(n8618), .ZN(N5044) );
  AOI22D1BWP30P140LVT U12567 ( .A1(i_data_bus[604]), .A2(n9936), .B1(
        i_data_bus[636]), .B2(n9933), .ZN(n8621) );
  AOI22D1BWP30P140LVT U12568 ( .A1(i_data_bus[572]), .A2(n9935), .B1(
        i_data_bus[540]), .B2(n9934), .ZN(n8620) );
  ND2D1BWP30P140LVT U12569 ( .A1(n8621), .A2(n8620), .ZN(N5421) );
  AOI22D1BWP30P140LVT U12570 ( .A1(i_data_bus[579]), .A2(n9936), .B1(
        i_data_bus[611]), .B2(n9933), .ZN(n8623) );
  AOI22D1BWP30P140LVT U12571 ( .A1(i_data_bus[547]), .A2(n9935), .B1(
        i_data_bus[515]), .B2(n9934), .ZN(n8622) );
  ND2D1BWP30P140LVT U12572 ( .A1(n8623), .A2(n8622), .ZN(N5396) );
  AOI22D1BWP30P140LVT U12573 ( .A1(i_data_bus[189]), .A2(n10219), .B1(
        i_data_bus[221]), .B2(n10218), .ZN(n8625) );
  AOI22D1BWP30P140LVT U12574 ( .A1(i_data_bus[157]), .A2(n6213), .B1(
        i_data_bus[253]), .B2(n10220), .ZN(n8624) );
  ND2D1BWP30P140LVT U12575 ( .A1(n8625), .A2(n8624), .ZN(N2434) );
  AOI22D1BWP30P140LVT U12576 ( .A1(i_data_bus[175]), .A2(n10219), .B1(
        i_data_bus[207]), .B2(n10218), .ZN(n8627) );
  AOI22D1BWP30P140LVT U12577 ( .A1(i_data_bus[143]), .A2(n6213), .B1(
        i_data_bus[239]), .B2(n10220), .ZN(n8626) );
  ND2D1BWP30P140LVT U12578 ( .A1(n8627), .A2(n8626), .ZN(N2420) );
  AOI22D1BWP30P140LVT U12579 ( .A1(i_data_bus[137]), .A2(n6213), .B1(
        i_data_bus[201]), .B2(n10218), .ZN(n8629) );
  AOI22D1BWP30P140LVT U12580 ( .A1(i_data_bus[169]), .A2(n10219), .B1(
        i_data_bus[233]), .B2(n10220), .ZN(n8628) );
  ND2D1BWP30P140LVT U12581 ( .A1(n8629), .A2(n8628), .ZN(N2414) );
  AOI22D1BWP30P140LVT U12582 ( .A1(i_data_bus[536]), .A2(n10182), .B1(
        i_data_bus[632]), .B2(n10185), .ZN(n8631) );
  AOI22D1BWP30P140LVT U12583 ( .A1(i_data_bus[568]), .A2(n10184), .B1(
        i_data_bus[600]), .B2(n10183), .ZN(n8630) );
  ND2D1BWP30P140LVT U12584 ( .A1(n8631), .A2(n8630), .ZN(N6907) );
  AOI22D1BWP30P140LVT U12585 ( .A1(i_data_bus[562]), .A2(n10184), .B1(
        i_data_bus[626]), .B2(n10185), .ZN(n8633) );
  AOI22D1BWP30P140LVT U12586 ( .A1(i_data_bus[530]), .A2(n10182), .B1(
        i_data_bus[594]), .B2(n10183), .ZN(n8632) );
  ND2D1BWP30P140LVT U12587 ( .A1(n8633), .A2(n8632), .ZN(N6901) );
  AOI22D1BWP30P140LVT U12588 ( .A1(i_data_bus[556]), .A2(n10184), .B1(
        i_data_bus[620]), .B2(n10185), .ZN(n8635) );
  AOI22D1BWP30P140LVT U12589 ( .A1(i_data_bus[524]), .A2(n10182), .B1(
        i_data_bus[588]), .B2(n10183), .ZN(n8634) );
  ND2D1BWP30P140LVT U12590 ( .A1(n8635), .A2(n8634), .ZN(N6895) );
  AOI22D1BWP30P140LVT U12591 ( .A1(i_data_bus[550]), .A2(n10184), .B1(
        i_data_bus[614]), .B2(n10185), .ZN(n8637) );
  AOI22D1BWP30P140LVT U12592 ( .A1(i_data_bus[518]), .A2(n10182), .B1(
        i_data_bus[582]), .B2(n10183), .ZN(n8636) );
  ND2D1BWP30P140LVT U12593 ( .A1(n8637), .A2(n8636), .ZN(N6889) );
  AOI22D1BWP30P140LVT U12594 ( .A1(i_data_bus[516]), .A2(n10182), .B1(
        i_data_bus[612]), .B2(n10185), .ZN(n8639) );
  AOI22D1BWP30P140LVT U12595 ( .A1(i_data_bus[548]), .A2(n10184), .B1(
        i_data_bus[580]), .B2(n10183), .ZN(n8638) );
  ND2D1BWP30P140LVT U12596 ( .A1(n8639), .A2(n8638), .ZN(N6887) );
  AOI22D1BWP30P140LVT U12597 ( .A1(i_data_bus[539]), .A2(n9934), .B1(
        i_data_bus[635]), .B2(n9933), .ZN(n8641) );
  AOI22D1BWP30P140LVT U12598 ( .A1(i_data_bus[571]), .A2(n9935), .B1(
        i_data_bus[603]), .B2(n9936), .ZN(n8640) );
  ND2D1BWP30P140LVT U12599 ( .A1(n8641), .A2(n8640), .ZN(N5420) );
  AOI22D1BWP30P140LVT U12600 ( .A1(i_data_bus[536]), .A2(n9934), .B1(
        i_data_bus[632]), .B2(n9933), .ZN(n8643) );
  AOI22D1BWP30P140LVT U12601 ( .A1(i_data_bus[568]), .A2(n9935), .B1(
        i_data_bus[600]), .B2(n9936), .ZN(n8642) );
  ND2D1BWP30P140LVT U12602 ( .A1(n8643), .A2(n8642), .ZN(N5417) );
  AOI22D1BWP30P140LVT U12603 ( .A1(i_data_bus[567]), .A2(n9935), .B1(
        i_data_bus[631]), .B2(n9933), .ZN(n8645) );
  AOI22D1BWP30P140LVT U12604 ( .A1(i_data_bus[535]), .A2(n9934), .B1(
        i_data_bus[599]), .B2(n9936), .ZN(n8644) );
  ND2D1BWP30P140LVT U12605 ( .A1(n8645), .A2(n8644), .ZN(N5416) );
  AOI22D1BWP30P140LVT U12606 ( .A1(i_data_bus[562]), .A2(n9935), .B1(
        i_data_bus[626]), .B2(n9933), .ZN(n8647) );
  AOI22D1BWP30P140LVT U12607 ( .A1(i_data_bus[530]), .A2(n9934), .B1(
        i_data_bus[594]), .B2(n9936), .ZN(n8646) );
  ND2D1BWP30P140LVT U12608 ( .A1(n8647), .A2(n8646), .ZN(N5411) );
  AOI22D1BWP30P140LVT U12609 ( .A1(i_data_bus[556]), .A2(n9935), .B1(
        i_data_bus[620]), .B2(n9933), .ZN(n8649) );
  AOI22D1BWP30P140LVT U12610 ( .A1(i_data_bus[524]), .A2(n9934), .B1(
        i_data_bus[588]), .B2(n9936), .ZN(n8648) );
  ND2D1BWP30P140LVT U12611 ( .A1(n8649), .A2(n8648), .ZN(N5405) );
  AOI22D1BWP30P140LVT U12612 ( .A1(i_data_bus[518]), .A2(n9934), .B1(
        i_data_bus[614]), .B2(n9933), .ZN(n8651) );
  AOI22D1BWP30P140LVT U12613 ( .A1(i_data_bus[550]), .A2(n9935), .B1(
        i_data_bus[582]), .B2(n9936), .ZN(n8650) );
  ND2D1BWP30P140LVT U12614 ( .A1(n8651), .A2(n8650), .ZN(N5399) );
  AOI22D1BWP30P140LVT U12615 ( .A1(i_data_bus[190]), .A2(n10034), .B1(
        i_data_bus[158]), .B2(n10026), .ZN(n8653) );
  AOI22D1BWP30P140LVT U12616 ( .A1(i_data_bus[222]), .A2(n10033), .B1(
        i_data_bus[254]), .B2(n10035), .ZN(n8652) );
  ND2D1BWP30P140LVT U12617 ( .A1(n8653), .A2(n8652), .ZN(N3541) );
  AOI22D1BWP30P140LVT U12618 ( .A1(i_data_bus[182]), .A2(n10034), .B1(
        i_data_bus[150]), .B2(n10026), .ZN(n8655) );
  AOI22D1BWP30P140LVT U12619 ( .A1(i_data_bus[214]), .A2(n10033), .B1(
        i_data_bus[246]), .B2(n10035), .ZN(n8654) );
  ND2D1BWP30P140LVT U12620 ( .A1(n8655), .A2(n8654), .ZN(N3533) );
  AOI22D1BWP30P140LVT U12621 ( .A1(i_data_bus[205]), .A2(n10033), .B1(
        i_data_bus[141]), .B2(n10026), .ZN(n8657) );
  AOI22D1BWP30P140LVT U12622 ( .A1(i_data_bus[173]), .A2(n10034), .B1(
        i_data_bus[237]), .B2(n10035), .ZN(n8656) );
  ND2D1BWP30P140LVT U12623 ( .A1(n8657), .A2(n8656), .ZN(N3524) );
  AOI22D1BWP30P140LVT U12624 ( .A1(i_data_bus[162]), .A2(n10034), .B1(
        i_data_bus[130]), .B2(n10026), .ZN(n8659) );
  AOI22D1BWP30P140LVT U12625 ( .A1(i_data_bus[194]), .A2(n10033), .B1(
        i_data_bus[226]), .B2(n10035), .ZN(n8658) );
  ND2D1BWP30P140LVT U12626 ( .A1(n8659), .A2(n8658), .ZN(N3513) );
  AOI22D1BWP30P140LVT U12627 ( .A1(i_data_bus[1008]), .A2(n9543), .B1(
        i_data_bus[976]), .B2(n9544), .ZN(n8661) );
  AOI22D1BWP30P140LVT U12628 ( .A1(i_data_bus[944]), .A2(n9545), .B1(
        i_data_bus[912]), .B2(n6226), .ZN(n8660) );
  ND2D1BWP30P140LVT U12629 ( .A1(n8661), .A2(n8660), .ZN(N2099) );
  AOI22D1BWP30P140LVT U12630 ( .A1(i_data_bus[932]), .A2(n9545), .B1(
        i_data_bus[964]), .B2(n9544), .ZN(n8663) );
  AOI22D1BWP30P140LVT U12631 ( .A1(i_data_bus[996]), .A2(n9543), .B1(
        i_data_bus[900]), .B2(n6226), .ZN(n8662) );
  ND2D1BWP30P140LVT U12632 ( .A1(n8663), .A2(n8662), .ZN(N2087) );
  AOI22D1BWP30P140LVT U12633 ( .A1(i_data_bus[571]), .A2(n10253), .B1(
        i_data_bus[603]), .B2(n10252), .ZN(n8665) );
  AOI22D1BWP30P140LVT U12634 ( .A1(i_data_bus[539]), .A2(n10245), .B1(
        i_data_bus[635]), .B2(n10254), .ZN(n8664) );
  ND2D1BWP30P140LVT U12635 ( .A1(n8665), .A2(n8664), .ZN(N9634) );
  AOI22D1BWP30P140LVT U12636 ( .A1(i_data_bus[568]), .A2(n10253), .B1(
        i_data_bus[600]), .B2(n10252), .ZN(n8667) );
  AOI22D1BWP30P140LVT U12637 ( .A1(i_data_bus[536]), .A2(n10245), .B1(
        i_data_bus[632]), .B2(n10254), .ZN(n8666) );
  ND2D1BWP30P140LVT U12638 ( .A1(n8667), .A2(n8666), .ZN(N9631) );
  AOI22D1BWP30P140LVT U12639 ( .A1(i_data_bus[551]), .A2(n10253), .B1(
        i_data_bus[519]), .B2(n10245), .ZN(n8669) );
  AOI22D1BWP30P140LVT U12640 ( .A1(i_data_bus[583]), .A2(n10252), .B1(
        i_data_bus[615]), .B2(n10254), .ZN(n8668) );
  ND2D1BWP30P140LVT U12641 ( .A1(n8669), .A2(n8668), .ZN(N9614) );
  AOI22D1BWP30P140LVT U12642 ( .A1(i_data_bus[995]), .A2(n9543), .B1(
        i_data_bus[963]), .B2(n9544), .ZN(n8671) );
  AOI22D1BWP30P140LVT U12643 ( .A1(i_data_bus[899]), .A2(n6226), .B1(
        i_data_bus[931]), .B2(n9545), .ZN(n8670) );
  ND2D1BWP30P140LVT U12644 ( .A1(n8671), .A2(n8670), .ZN(N2086) );
  AOI22D1BWP30P140LVT U12645 ( .A1(i_data_bus[1014]), .A2(n9543), .B1(
        i_data_bus[982]), .B2(n9544), .ZN(n8673) );
  AOI22D1BWP30P140LVT U12646 ( .A1(i_data_bus[918]), .A2(n6226), .B1(
        i_data_bus[950]), .B2(n9545), .ZN(n8672) );
  ND2D1BWP30P140LVT U12647 ( .A1(n8673), .A2(n8672), .ZN(N2105) );
  AOI22D1BWP30P140LVT U12648 ( .A1(i_data_bus[901]), .A2(n6226), .B1(
        i_data_bus[965]), .B2(n9544), .ZN(n8675) );
  AOI22D1BWP30P140LVT U12649 ( .A1(i_data_bus[933]), .A2(n9545), .B1(
        i_data_bus[997]), .B2(n9543), .ZN(n8674) );
  ND2D1BWP30P140LVT U12650 ( .A1(n8675), .A2(n8674), .ZN(N2088) );
  AOI22D1BWP30P140LVT U12651 ( .A1(i_data_bus[921]), .A2(n6226), .B1(
        i_data_bus[985]), .B2(n9544), .ZN(n8677) );
  AOI22D1BWP30P140LVT U12652 ( .A1(i_data_bus[953]), .A2(n9545), .B1(
        i_data_bus[1017]), .B2(n9543), .ZN(n8676) );
  ND2D1BWP30P140LVT U12653 ( .A1(n8677), .A2(n8676), .ZN(N2108) );
  AOI22D1BWP30P140LVT U12654 ( .A1(i_data_bus[920]), .A2(n6226), .B1(
        i_data_bus[984]), .B2(n9544), .ZN(n8679) );
  AOI22D1BWP30P140LVT U12655 ( .A1(i_data_bus[952]), .A2(n9545), .B1(
        i_data_bus[1016]), .B2(n9543), .ZN(n8678) );
  ND2D1BWP30P140LVT U12656 ( .A1(n8679), .A2(n8678), .ZN(N2107) );
  AOI22D1BWP30P140LVT U12657 ( .A1(i_data_bus[919]), .A2(n6226), .B1(
        i_data_bus[983]), .B2(n9544), .ZN(n8681) );
  AOI22D1BWP30P140LVT U12658 ( .A1(i_data_bus[951]), .A2(n9545), .B1(
        i_data_bus[1015]), .B2(n9543), .ZN(n8680) );
  ND2D1BWP30P140LVT U12659 ( .A1(n8681), .A2(n8680), .ZN(N2106) );
  AOI22D1BWP30P140LVT U12660 ( .A1(i_data_bus[913]), .A2(n6226), .B1(
        i_data_bus[977]), .B2(n9544), .ZN(n8683) );
  AOI22D1BWP30P140LVT U12661 ( .A1(i_data_bus[945]), .A2(n9545), .B1(
        i_data_bus[1009]), .B2(n9543), .ZN(n8682) );
  ND2D1BWP30P140LVT U12662 ( .A1(n8683), .A2(n8682), .ZN(N2100) );
  AOI22D1BWP30P140LVT U12663 ( .A1(i_data_bus[905]), .A2(n6226), .B1(
        i_data_bus[969]), .B2(n9544), .ZN(n8685) );
  AOI22D1BWP30P140LVT U12664 ( .A1(i_data_bus[937]), .A2(n9545), .B1(
        i_data_bus[1001]), .B2(n9543), .ZN(n8684) );
  ND2D1BWP30P140LVT U12665 ( .A1(n8685), .A2(n8684), .ZN(N2092) );
  AOI22D1BWP30P140LVT U12666 ( .A1(i_data_bus[376]), .A2(n9877), .B1(
        i_data_bus[344]), .B2(n9879), .ZN(n8687) );
  AOI22D1BWP30P140LVT U12667 ( .A1(i_data_bus[312]), .A2(n9878), .B1(
        i_data_bus[280]), .B2(n6217), .ZN(n8686) );
  ND2D1BWP30P140LVT U12668 ( .A1(n8687), .A2(n8686), .ZN(N10689) );
  AOI22D1BWP30P140LVT U12669 ( .A1(i_data_bus[361]), .A2(n9877), .B1(
        i_data_bus[329]), .B2(n9879), .ZN(n8689) );
  AOI22D1BWP30P140LVT U12670 ( .A1(i_data_bus[297]), .A2(n9878), .B1(
        i_data_bus[265]), .B2(n6217), .ZN(n8688) );
  ND2D1BWP30P140LVT U12671 ( .A1(n8689), .A2(n8688), .ZN(N10674) );
  AOI22D1BWP30P140LVT U12672 ( .A1(i_data_bus[289]), .A2(n9843), .B1(
        i_data_bus[321]), .B2(n9844), .ZN(n8691) );
  AOI22D1BWP30P140LVT U12673 ( .A1(i_data_bus[353]), .A2(n9845), .B1(
        i_data_bus[257]), .B2(n9846), .ZN(n8690) );
  ND2D1BWP30P140LVT U12674 ( .A1(n8691), .A2(n8690), .ZN(N7942) );
  NR4D1BWP30P140LVT U12675 ( .A1(i_cmd[76]), .A2(n8692), .A3(n10392), .A4(
        n11037), .ZN(n10051) );
  INR4D1BWP30P140LVT U12676 ( .A1(i_cmd[84]), .B1(i_cmd[68]), .B2(n10395), 
        .B3(n11034), .ZN(n10054) );
  AOI22D1BWP30P140LVT U12677 ( .A1(i_data_bus[361]), .A2(n10051), .B1(
        i_data_bus[329]), .B2(n10054), .ZN(n8694) );
  NR4D1BWP30P140LVT U12678 ( .A1(i_cmd[92]), .A2(n8692), .A3(n10391), .A4(
        n11036), .ZN(n10053) );
  NR3D0P7BWP30P140LVT U12679 ( .A1(i_cmd[84]), .A2(i_cmd[92]), .A3(i_cmd[76]), 
        .ZN(n11033) );
  AOI22D1BWP30P140LVT U12680 ( .A1(i_data_bus[297]), .A2(n10053), .B1(
        i_data_bus[265]), .B2(n10052), .ZN(n8693) );
  ND2D1BWP30P140LVT U12681 ( .A1(n8694), .A2(n8693), .ZN(N6460) );
  AOI22D1BWP30P140LVT U12682 ( .A1(i_data_bus[373]), .A2(n10051), .B1(
        i_data_bus[341]), .B2(n10054), .ZN(n8696) );
  AOI22D1BWP30P140LVT U12683 ( .A1(i_data_bus[309]), .A2(n10053), .B1(
        i_data_bus[277]), .B2(n10052), .ZN(n8695) );
  ND2D1BWP30P140LVT U12684 ( .A1(n8696), .A2(n8695), .ZN(N6472) );
  AOI22D1BWP30P140LVT U12685 ( .A1(n8722), .A2(i_data_bus[897]), .B1(n8719), 
        .B2(i_data_bus[993]), .ZN(n8698) );
  AOI22D1BWP30P140LVT U12686 ( .A1(n8720), .A2(i_data_bus[929]), .B1(n8721), 
        .B2(i_data_bus[961]), .ZN(n8697) );
  ND2D1BWP30P140LVT U12687 ( .A1(n8698), .A2(n8697), .ZN(N2934) );
  AOI22D1BWP30P140LVT U12688 ( .A1(n8722), .A2(i_data_bus[902]), .B1(n8719), 
        .B2(i_data_bus[998]), .ZN(n8700) );
  AOI22D1BWP30P140LVT U12689 ( .A1(n8720), .A2(i_data_bus[934]), .B1(n8721), 
        .B2(i_data_bus[966]), .ZN(n8699) );
  ND2D1BWP30P140LVT U12690 ( .A1(n8700), .A2(n8699), .ZN(N2939) );
  AOI22D1BWP30P140LVT U12691 ( .A1(n8720), .A2(i_data_bus[937]), .B1(n8719), 
        .B2(i_data_bus[1001]), .ZN(n8702) );
  AOI22D1BWP30P140LVT U12692 ( .A1(n8722), .A2(i_data_bus[905]), .B1(n8721), 
        .B2(i_data_bus[969]), .ZN(n8701) );
  ND2D1BWP30P140LVT U12693 ( .A1(n8702), .A2(n8701), .ZN(N2942) );
  AOI22D1BWP30P140LVT U12694 ( .A1(n8722), .A2(i_data_bus[903]), .B1(n8719), 
        .B2(i_data_bus[999]), .ZN(n8704) );
  AOI22D1BWP30P140LVT U12695 ( .A1(n8720), .A2(i_data_bus[935]), .B1(n8721), 
        .B2(i_data_bus[967]), .ZN(n8703) );
  ND2D1BWP30P140LVT U12696 ( .A1(n8704), .A2(n8703), .ZN(N2940) );
  AOI22D1BWP30P140LVT U12697 ( .A1(n8722), .A2(i_data_bus[907]), .B1(n8719), 
        .B2(i_data_bus[1003]), .ZN(n8706) );
  AOI22D1BWP30P140LVT U12698 ( .A1(n8720), .A2(i_data_bus[939]), .B1(n8721), 
        .B2(i_data_bus[971]), .ZN(n8705) );
  ND2D1BWP30P140LVT U12699 ( .A1(n8706), .A2(n8705), .ZN(N2944) );
  AOI22D1BWP30P140LVT U12700 ( .A1(n8720), .A2(i_data_bus[941]), .B1(n8719), 
        .B2(i_data_bus[1005]), .ZN(n8708) );
  AOI22D1BWP30P140LVT U12701 ( .A1(n8722), .A2(i_data_bus[909]), .B1(n8721), 
        .B2(i_data_bus[973]), .ZN(n8707) );
  ND2D1BWP30P140LVT U12702 ( .A1(n8708), .A2(n8707), .ZN(N2946) );
  AOI22D1BWP30P140LVT U12703 ( .A1(n8720), .A2(i_data_bus[940]), .B1(n8719), 
        .B2(i_data_bus[1004]), .ZN(n8710) );
  AOI22D1BWP30P140LVT U12704 ( .A1(n8722), .A2(i_data_bus[908]), .B1(n8721), 
        .B2(i_data_bus[972]), .ZN(n8709) );
  ND2D1BWP30P140LVT U12705 ( .A1(n8710), .A2(n8709), .ZN(N2945) );
  AOI22D1BWP30P140LVT U12706 ( .A1(n8722), .A2(i_data_bus[911]), .B1(n8719), 
        .B2(i_data_bus[1007]), .ZN(n8712) );
  AOI22D1BWP30P140LVT U12707 ( .A1(n8720), .A2(i_data_bus[943]), .B1(n8721), 
        .B2(i_data_bus[975]), .ZN(n8711) );
  ND2D1BWP30P140LVT U12708 ( .A1(n8712), .A2(n8711), .ZN(N2948) );
  AOI22D1BWP30P140LVT U12709 ( .A1(n8720), .A2(i_data_bus[955]), .B1(n8719), 
        .B2(i_data_bus[1019]), .ZN(n8714) );
  AOI22D1BWP30P140LVT U12710 ( .A1(n8722), .A2(i_data_bus[923]), .B1(n8721), 
        .B2(i_data_bus[987]), .ZN(n8713) );
  ND2D1BWP30P140LVT U12711 ( .A1(n8714), .A2(n8713), .ZN(N2960) );
  AOI22D1BWP30P140LVT U12712 ( .A1(n8722), .A2(i_data_bus[917]), .B1(n8719), 
        .B2(i_data_bus[1013]), .ZN(n8716) );
  AOI22D1BWP30P140LVT U12713 ( .A1(n8720), .A2(i_data_bus[949]), .B1(n8721), 
        .B2(i_data_bus[981]), .ZN(n8715) );
  ND2D1BWP30P140LVT U12714 ( .A1(n8716), .A2(n8715), .ZN(N2954) );
  AOI22D1BWP30P140LVT U12715 ( .A1(n8720), .A2(i_data_bus[947]), .B1(n8719), 
        .B2(i_data_bus[1011]), .ZN(n8718) );
  AOI22D1BWP30P140LVT U12716 ( .A1(n8722), .A2(i_data_bus[915]), .B1(n8721), 
        .B2(i_data_bus[979]), .ZN(n8717) );
  ND2D1BWP30P140LVT U12717 ( .A1(n8718), .A2(n8717), .ZN(N2952) );
  AOI22D1BWP30P140LVT U12718 ( .A1(n8720), .A2(i_data_bus[945]), .B1(n8719), 
        .B2(i_data_bus[1009]), .ZN(n8724) );
  AOI22D1BWP30P140LVT U12719 ( .A1(n8722), .A2(i_data_bus[913]), .B1(n8721), 
        .B2(i_data_bus[977]), .ZN(n8723) );
  ND2D1BWP30P140LVT U12720 ( .A1(n8724), .A2(n8723), .ZN(N2950) );
  AOI22D1BWP30P140LVT U12721 ( .A1(i_data_bus[376]), .A2(n9845), .B1(
        i_data_bus[344]), .B2(n9844), .ZN(n8726) );
  AOI22D1BWP30P140LVT U12722 ( .A1(i_data_bus[312]), .A2(n9843), .B1(
        i_data_bus[280]), .B2(n9846), .ZN(n8725) );
  ND2D1BWP30P140LVT U12723 ( .A1(n8726), .A2(n8725), .ZN(N7965) );
  AOI22D1BWP30P140LVT U12724 ( .A1(i_data_bus[143]), .A2(n9318), .B1(
        i_data_bus[207]), .B2(n10039), .ZN(n8728) );
  AOI22D1BWP30P140LVT U12725 ( .A1(i_data_bus[175]), .A2(n10040), .B1(
        i_data_bus[239]), .B2(n10038), .ZN(n8727) );
  ND2D1BWP30P140LVT U12726 ( .A1(n8728), .A2(n8727), .ZN(N8974) );
  AOI22D1BWP30P140LVT U12727 ( .A1(i_data_bus[189]), .A2(n10040), .B1(
        i_data_bus[221]), .B2(n10039), .ZN(n8730) );
  AOI22D1BWP30P140LVT U12728 ( .A1(i_data_bus[157]), .A2(n9318), .B1(
        i_data_bus[253]), .B2(n10038), .ZN(n8729) );
  ND2D1BWP30P140LVT U12729 ( .A1(n8730), .A2(n8729), .ZN(N8988) );
  AOI22D1BWP30P140LVT U12730 ( .A1(i_data_bus[147]), .A2(n9318), .B1(
        i_data_bus[211]), .B2(n10039), .ZN(n8732) );
  AOI22D1BWP30P140LVT U12731 ( .A1(i_data_bus[179]), .A2(n10040), .B1(
        i_data_bus[243]), .B2(n10038), .ZN(n8731) );
  ND2D1BWP30P140LVT U12732 ( .A1(n8732), .A2(n8731), .ZN(N8978) );
  AOI22D1BWP30P140LVT U12733 ( .A1(i_data_bus[177]), .A2(n10040), .B1(
        i_data_bus[145]), .B2(n9318), .ZN(n8734) );
  AOI22D1BWP30P140LVT U12734 ( .A1(i_data_bus[209]), .A2(n10039), .B1(
        i_data_bus[241]), .B2(n10038), .ZN(n8733) );
  ND2D1BWP30P140LVT U12735 ( .A1(n8734), .A2(n8733), .ZN(N8976) );
  AOI22D1BWP30P140LVT U12736 ( .A1(i_data_bus[176]), .A2(n10040), .B1(
        i_data_bus[208]), .B2(n10039), .ZN(n8736) );
  AOI22D1BWP30P140LVT U12737 ( .A1(i_data_bus[144]), .A2(n9318), .B1(
        i_data_bus[240]), .B2(n10038), .ZN(n8735) );
  ND2D1BWP30P140LVT U12738 ( .A1(n8736), .A2(n8735), .ZN(N8975) );
  AOI22D1BWP30P140LVT U12739 ( .A1(i_data_bus[140]), .A2(n9318), .B1(
        i_data_bus[204]), .B2(n10039), .ZN(n8738) );
  AOI22D1BWP30P140LVT U12740 ( .A1(i_data_bus[172]), .A2(n10040), .B1(
        i_data_bus[236]), .B2(n10038), .ZN(n8737) );
  ND2D1BWP30P140LVT U12741 ( .A1(n8738), .A2(n8737), .ZN(N8971) );
  AOI22D1BWP30P140LVT U12742 ( .A1(i_data_bus[139]), .A2(n9318), .B1(
        i_data_bus[203]), .B2(n10039), .ZN(n8740) );
  AOI22D1BWP30P140LVT U12743 ( .A1(i_data_bus[171]), .A2(n10040), .B1(
        i_data_bus[235]), .B2(n10038), .ZN(n8739) );
  ND2D1BWP30P140LVT U12744 ( .A1(n8740), .A2(n8739), .ZN(N8970) );
  AOI22D1BWP30P140LVT U12745 ( .A1(i_data_bus[604]), .A2(n10001), .B1(
        i_data_bus[540]), .B2(n6222), .ZN(n8742) );
  AOI22D1BWP30P140LVT U12746 ( .A1(i_data_bus[572]), .A2(n10002), .B1(
        i_data_bus[636]), .B2(n10003), .ZN(n8741) );
  ND2D1BWP30P140LVT U12747 ( .A1(n8742), .A2(n8741), .ZN(N4187) );
  AOI22D1BWP30P140LVT U12748 ( .A1(i_data_bus[603]), .A2(n10001), .B1(
        i_data_bus[539]), .B2(n6222), .ZN(n8744) );
  AOI22D1BWP30P140LVT U12749 ( .A1(i_data_bus[571]), .A2(n10002), .B1(
        i_data_bus[635]), .B2(n10003), .ZN(n8743) );
  ND2D1BWP30P140LVT U12750 ( .A1(n8744), .A2(n8743), .ZN(N4186) );
  AOI22D1BWP30P140LVT U12751 ( .A1(i_data_bus[570]), .A2(n10002), .B1(
        i_data_bus[602]), .B2(n10001), .ZN(n8746) );
  AOI22D1BWP30P140LVT U12752 ( .A1(i_data_bus[538]), .A2(n6222), .B1(
        i_data_bus[634]), .B2(n10003), .ZN(n8745) );
  ND2D1BWP30P140LVT U12753 ( .A1(n8746), .A2(n8745), .ZN(N4185) );
  AOI22D1BWP30P140LVT U12754 ( .A1(i_data_bus[568]), .A2(n10002), .B1(
        i_data_bus[536]), .B2(n6222), .ZN(n8748) );
  AOI22D1BWP30P140LVT U12755 ( .A1(i_data_bus[600]), .A2(n10001), .B1(
        i_data_bus[632]), .B2(n10003), .ZN(n8747) );
  ND2D1BWP30P140LVT U12756 ( .A1(n8748), .A2(n8747), .ZN(N4183) );
  AOI22D1BWP30P140LVT U12757 ( .A1(i_data_bus[561]), .A2(n10002), .B1(
        i_data_bus[593]), .B2(n10001), .ZN(n8750) );
  AOI22D1BWP30P140LVT U12758 ( .A1(i_data_bus[529]), .A2(n6222), .B1(
        i_data_bus[625]), .B2(n10003), .ZN(n8749) );
  ND2D1BWP30P140LVT U12759 ( .A1(n8750), .A2(n8749), .ZN(N4176) );
  AOI22D1BWP30P140LVT U12760 ( .A1(i_data_bus[550]), .A2(n10002), .B1(
        i_data_bus[582]), .B2(n10001), .ZN(n8752) );
  AOI22D1BWP30P140LVT U12761 ( .A1(i_data_bus[518]), .A2(n6222), .B1(
        i_data_bus[614]), .B2(n10003), .ZN(n8751) );
  ND2D1BWP30P140LVT U12762 ( .A1(n8752), .A2(n8751), .ZN(N4165) );
  AOI22D1BWP30P140LVT U12763 ( .A1(i_data_bus[547]), .A2(n10002), .B1(
        i_data_bus[515]), .B2(n6222), .ZN(n8754) );
  AOI22D1BWP30P140LVT U12764 ( .A1(i_data_bus[579]), .A2(n10001), .B1(
        i_data_bus[611]), .B2(n10003), .ZN(n8753) );
  ND2D1BWP30P140LVT U12765 ( .A1(n8754), .A2(n8753), .ZN(N4162) );
  AOI22D1BWP30P140LVT U12766 ( .A1(i_data_bus[376]), .A2(n9730), .B1(
        i_data_bus[344]), .B2(n9731), .ZN(n8756) );
  AOI22D1BWP30P140LVT U12767 ( .A1(i_data_bus[312]), .A2(n9732), .B1(
        i_data_bus[280]), .B2(n6219), .ZN(n8755) );
  ND2D1BWP30P140LVT U12768 ( .A1(n8756), .A2(n8755), .ZN(N3751) );
  AOI22D1BWP30P140LVT U12769 ( .A1(i_data_bus[373]), .A2(n9730), .B1(
        i_data_bus[341]), .B2(n9731), .ZN(n8758) );
  AOI22D1BWP30P140LVT U12770 ( .A1(i_data_bus[309]), .A2(n9732), .B1(
        i_data_bus[277]), .B2(n6219), .ZN(n8757) );
  ND2D1BWP30P140LVT U12771 ( .A1(n8758), .A2(n8757), .ZN(N3748) );
  AOI22D1BWP30P140LVT U12772 ( .A1(i_data_bus[361]), .A2(n9730), .B1(
        i_data_bus[329]), .B2(n9731), .ZN(n8760) );
  AOI22D1BWP30P140LVT U12773 ( .A1(i_data_bus[297]), .A2(n9732), .B1(
        i_data_bus[265]), .B2(n6219), .ZN(n8759) );
  ND2D1BWP30P140LVT U12774 ( .A1(n8760), .A2(n8759), .ZN(N3736) );
  AOI22D1BWP30P140LVT U12775 ( .A1(i_data_bus[243]), .A2(n10035), .B1(
        i_data_bus[211]), .B2(n10033), .ZN(n8762) );
  AOI22D1BWP30P140LVT U12776 ( .A1(i_data_bus[179]), .A2(n10034), .B1(
        i_data_bus[147]), .B2(n10026), .ZN(n8761) );
  ND2D1BWP30P140LVT U12777 ( .A1(n8762), .A2(n8761), .ZN(N3530) );
  AOI22D1BWP30P140LVT U12778 ( .A1(i_data_bus[98]), .A2(n9915), .B1(
        i_data_bus[66]), .B2(n9914), .ZN(n8764) );
  AOI22D1BWP30P140LVT U12779 ( .A1(i_data_bus[34]), .A2(n9916), .B1(
        i_data_bus[2]), .B2(n6218), .ZN(n8763) );
  ND2D1BWP30P140LVT U12780 ( .A1(n8764), .A2(n8763), .ZN(N3297) );
  AOI22D1BWP30P140LVT U12781 ( .A1(i_data_bus[161]), .A2(n10034), .B1(
        i_data_bus[193]), .B2(n10033), .ZN(n8766) );
  AOI22D1BWP30P140LVT U12782 ( .A1(i_data_bus[225]), .A2(n10035), .B1(
        i_data_bus[129]), .B2(n10026), .ZN(n8765) );
  ND2D1BWP30P140LVT U12783 ( .A1(n8766), .A2(n8765), .ZN(N3512) );
  AOI22D1BWP30P140LVT U12784 ( .A1(i_data_bus[187]), .A2(n10034), .B1(
        i_data_bus[219]), .B2(n10033), .ZN(n8768) );
  AOI22D1BWP30P140LVT U12785 ( .A1(i_data_bus[155]), .A2(n10026), .B1(
        i_data_bus[251]), .B2(n10035), .ZN(n8767) );
  ND2D1BWP30P140LVT U12786 ( .A1(n8768), .A2(n8767), .ZN(N3538) );
  AOI22D1BWP30P140LVT U12787 ( .A1(i_data_bus[154]), .A2(n10026), .B1(
        i_data_bus[218]), .B2(n10033), .ZN(n8770) );
  AOI22D1BWP30P140LVT U12788 ( .A1(i_data_bus[186]), .A2(n10034), .B1(
        i_data_bus[250]), .B2(n10035), .ZN(n8769) );
  ND2D1BWP30P140LVT U12789 ( .A1(n8770), .A2(n8769), .ZN(N3537) );
  AOI22D1BWP30P140LVT U12790 ( .A1(i_data_bus[175]), .A2(n10034), .B1(
        i_data_bus[207]), .B2(n10033), .ZN(n8772) );
  AOI22D1BWP30P140LVT U12791 ( .A1(i_data_bus[143]), .A2(n10026), .B1(
        i_data_bus[239]), .B2(n10035), .ZN(n8771) );
  ND2D1BWP30P140LVT U12792 ( .A1(n8772), .A2(n8771), .ZN(N3526) );
  AOI22D1BWP30P140LVT U12793 ( .A1(i_data_bus[189]), .A2(n10034), .B1(
        i_data_bus[221]), .B2(n10033), .ZN(n8774) );
  AOI22D1BWP30P140LVT U12794 ( .A1(i_data_bus[157]), .A2(n10026), .B1(
        i_data_bus[253]), .B2(n10035), .ZN(n8773) );
  ND2D1BWP30P140LVT U12795 ( .A1(n8774), .A2(n8773), .ZN(N3540) );
  AOI22D1BWP30P140LVT U12796 ( .A1(i_data_bus[190]), .A2(n10133), .B1(
        i_data_bus[158]), .B2(n10134), .ZN(n8776) );
  AOI22D1BWP30P140LVT U12797 ( .A1(i_data_bus[222]), .A2(n10132), .B1(
        i_data_bus[254]), .B2(n10131), .ZN(n8775) );
  ND2D1BWP30P140LVT U12798 ( .A1(n8776), .A2(n8775), .ZN(N7883) );
  AOI22D1BWP30P140LVT U12799 ( .A1(i_data_bus[156]), .A2(n10134), .B1(
        i_data_bus[220]), .B2(n10132), .ZN(n8778) );
  AOI22D1BWP30P140LVT U12800 ( .A1(i_data_bus[188]), .A2(n10133), .B1(
        i_data_bus[252]), .B2(n10131), .ZN(n8777) );
  ND2D1BWP30P140LVT U12801 ( .A1(n8778), .A2(n8777), .ZN(N7881) );
  AOI22D1BWP30P140LVT U12802 ( .A1(i_data_bus[182]), .A2(n10133), .B1(
        i_data_bus[150]), .B2(n10134), .ZN(n8780) );
  AOI22D1BWP30P140LVT U12803 ( .A1(i_data_bus[214]), .A2(n10132), .B1(
        i_data_bus[246]), .B2(n10131), .ZN(n8779) );
  ND2D1BWP30P140LVT U12804 ( .A1(n8780), .A2(n8779), .ZN(N7875) );
  AOI22D1BWP30P140LVT U12805 ( .A1(i_data_bus[209]), .A2(n10132), .B1(
        i_data_bus[145]), .B2(n10134), .ZN(n8782) );
  AOI22D1BWP30P140LVT U12806 ( .A1(i_data_bus[177]), .A2(n10133), .B1(
        i_data_bus[241]), .B2(n10131), .ZN(n8781) );
  ND2D1BWP30P140LVT U12807 ( .A1(n8782), .A2(n8781), .ZN(N7870) );
  AOI22D1BWP30P140LVT U12808 ( .A1(i_data_bus[144]), .A2(n10134), .B1(
        i_data_bus[208]), .B2(n10132), .ZN(n8784) );
  AOI22D1BWP30P140LVT U12809 ( .A1(i_data_bus[176]), .A2(n10133), .B1(
        i_data_bus[240]), .B2(n10131), .ZN(n8783) );
  ND2D1BWP30P140LVT U12810 ( .A1(n8784), .A2(n8783), .ZN(N7869) );
  AOI22D1BWP30P140LVT U12811 ( .A1(i_data_bus[137]), .A2(n10134), .B1(
        i_data_bus[201]), .B2(n10132), .ZN(n8786) );
  AOI22D1BWP30P140LVT U12812 ( .A1(i_data_bus[169]), .A2(n10133), .B1(
        i_data_bus[233]), .B2(n10131), .ZN(n8785) );
  ND2D1BWP30P140LVT U12813 ( .A1(n8786), .A2(n8785), .ZN(N7862) );
  AOI22D1BWP30P140LVT U12814 ( .A1(i_data_bus[162]), .A2(n10133), .B1(
        i_data_bus[130]), .B2(n10134), .ZN(n8788) );
  AOI22D1BWP30P140LVT U12815 ( .A1(i_data_bus[194]), .A2(n10132), .B1(
        i_data_bus[226]), .B2(n10131), .ZN(n8787) );
  ND2D1BWP30P140LVT U12816 ( .A1(n8788), .A2(n8787), .ZN(N7855) );
  AOI22D1BWP30P140LVT U12817 ( .A1(i_data_bus[129]), .A2(n10134), .B1(
        i_data_bus[193]), .B2(n10132), .ZN(n8790) );
  AOI22D1BWP30P140LVT U12818 ( .A1(i_data_bus[161]), .A2(n10133), .B1(
        i_data_bus[225]), .B2(n10131), .ZN(n8789) );
  ND2D1BWP30P140LVT U12819 ( .A1(n8790), .A2(n8789), .ZN(N7854) );
  AOI22D1BWP30P140LVT U12820 ( .A1(i_data_bus[139]), .A2(n10134), .B1(
        i_data_bus[203]), .B2(n10132), .ZN(n8792) );
  AOI22D1BWP30P140LVT U12821 ( .A1(i_data_bus[171]), .A2(n10133), .B1(
        i_data_bus[235]), .B2(n10131), .ZN(n8791) );
  ND2D1BWP30P140LVT U12822 ( .A1(n8792), .A2(n8791), .ZN(N7864) );
  AOI22D1BWP30P140LVT U12823 ( .A1(i_data_bus[1022]), .A2(n9663), .B1(
        i_data_bus[990]), .B2(n9662), .ZN(n8794) );
  AOI22D1BWP30P140LVT U12824 ( .A1(i_data_bus[958]), .A2(n9660), .B1(
        i_data_bus[926]), .B2(n9661), .ZN(n8793) );
  ND2D1BWP30P140LVT U12825 ( .A1(n8794), .A2(n8793), .ZN(N7561) );
  AOI22D1BWP30P140LVT U12826 ( .A1(i_data_bus[1012]), .A2(n9663), .B1(
        i_data_bus[980]), .B2(n9662), .ZN(n8796) );
  AOI22D1BWP30P140LVT U12827 ( .A1(i_data_bus[948]), .A2(n9660), .B1(
        i_data_bus[916]), .B2(n9661), .ZN(n8795) );
  ND2D1BWP30P140LVT U12828 ( .A1(n8796), .A2(n8795), .ZN(N7551) );
  AOI22D1BWP30P140LVT U12829 ( .A1(i_data_bus[944]), .A2(n9660), .B1(
        i_data_bus[976]), .B2(n9662), .ZN(n8798) );
  AOI22D1BWP30P140LVT U12830 ( .A1(i_data_bus[1008]), .A2(n9663), .B1(
        i_data_bus[912]), .B2(n9661), .ZN(n8797) );
  ND2D1BWP30P140LVT U12831 ( .A1(n8798), .A2(n8797), .ZN(N7547) );
  AOI22D1BWP30P140LVT U12832 ( .A1(i_data_bus[939]), .A2(n9660), .B1(
        i_data_bus[971]), .B2(n9662), .ZN(n8800) );
  AOI22D1BWP30P140LVT U12833 ( .A1(i_data_bus[1003]), .A2(n9663), .B1(
        i_data_bus[907]), .B2(n9661), .ZN(n8799) );
  ND2D1BWP30P140LVT U12834 ( .A1(n8800), .A2(n8799), .ZN(N7542) );
  AOI22D1BWP30P140LVT U12835 ( .A1(i_data_bus[1017]), .A2(n9663), .B1(
        i_data_bus[985]), .B2(n9662), .ZN(n8802) );
  AOI22D1BWP30P140LVT U12836 ( .A1(i_data_bus[921]), .A2(n9661), .B1(
        i_data_bus[953]), .B2(n9660), .ZN(n8801) );
  ND2D1BWP30P140LVT U12837 ( .A1(n8802), .A2(n8801), .ZN(N7556) );
  AOI22D1BWP30P140LVT U12838 ( .A1(i_data_bus[995]), .A2(n9663), .B1(
        i_data_bus[963]), .B2(n9662), .ZN(n8804) );
  AOI22D1BWP30P140LVT U12839 ( .A1(i_data_bus[899]), .A2(n9661), .B1(
        i_data_bus[931]), .B2(n9660), .ZN(n8803) );
  ND2D1BWP30P140LVT U12840 ( .A1(n8804), .A2(n8803), .ZN(N7534) );
  AOI22D1BWP30P140LVT U12841 ( .A1(i_data_bus[925]), .A2(n9661), .B1(
        i_data_bus[989]), .B2(n9662), .ZN(n8806) );
  AOI22D1BWP30P140LVT U12842 ( .A1(i_data_bus[957]), .A2(n9660), .B1(
        i_data_bus[1021]), .B2(n9663), .ZN(n8805) );
  ND2D1BWP30P140LVT U12843 ( .A1(n8806), .A2(n8805), .ZN(N7560) );
  AOI22D1BWP30P140LVT U12844 ( .A1(i_data_bus[922]), .A2(n9661), .B1(
        i_data_bus[986]), .B2(n9662), .ZN(n8808) );
  AOI22D1BWP30P140LVT U12845 ( .A1(i_data_bus[954]), .A2(n9660), .B1(
        i_data_bus[1018]), .B2(n9663), .ZN(n8807) );
  ND2D1BWP30P140LVT U12846 ( .A1(n8808), .A2(n8807), .ZN(N7557) );
  AOI22D1BWP30P140LVT U12847 ( .A1(i_data_bus[943]), .A2(n9660), .B1(
        i_data_bus[975]), .B2(n9662), .ZN(n8810) );
  AOI22D1BWP30P140LVT U12848 ( .A1(i_data_bus[911]), .A2(n9661), .B1(
        i_data_bus[1007]), .B2(n9663), .ZN(n8809) );
  ND2D1BWP30P140LVT U12849 ( .A1(n8810), .A2(n8809), .ZN(N7546) );
  AOI22D1BWP30P140LVT U12850 ( .A1(i_data_bus[898]), .A2(n9661), .B1(
        i_data_bus[962]), .B2(n9662), .ZN(n8812) );
  AOI22D1BWP30P140LVT U12851 ( .A1(i_data_bus[930]), .A2(n9660), .B1(
        i_data_bus[994]), .B2(n9663), .ZN(n8811) );
  ND2D1BWP30P140LVT U12852 ( .A1(n8812), .A2(n8811), .ZN(N7533) );
  AOI22D1BWP30P140LVT U12853 ( .A1(i_data_bus[896]), .A2(n9661), .B1(
        i_data_bus[960]), .B2(n9662), .ZN(n8814) );
  AOI22D1BWP30P140LVT U12854 ( .A1(i_data_bus[928]), .A2(n9660), .B1(
        i_data_bus[992]), .B2(n9663), .ZN(n8813) );
  ND2D1BWP30P140LVT U12855 ( .A1(n8814), .A2(n8813), .ZN(N7531) );
  AOI22D1BWP30P140LVT U12856 ( .A1(i_data_bus[435]), .A2(n10386), .B1(
        i_data_bus[499]), .B2(n10385), .ZN(n8816) );
  AOI22D1BWP30P140LVT U12857 ( .A1(i_data_bus[403]), .A2(n10387), .B1(
        i_data_bus[467]), .B2(n10388), .ZN(n8815) );
  ND2D1BWP30P140LVT U12858 ( .A1(n8816), .A2(n8815), .ZN(N10772) );
  AOI22D1BWP30P140LVT U12859 ( .A1(i_data_bus[426]), .A2(n10386), .B1(
        i_data_bus[490]), .B2(n10385), .ZN(n8818) );
  AOI22D1BWP30P140LVT U12860 ( .A1(i_data_bus[394]), .A2(n10387), .B1(
        i_data_bus[458]), .B2(n10388), .ZN(n8817) );
  ND2D1BWP30P140LVT U12861 ( .A1(n8818), .A2(n8817), .ZN(N10763) );
  AOI22D1BWP30P140LVT U12862 ( .A1(i_data_bus[422]), .A2(n10386), .B1(
        i_data_bus[486]), .B2(n10385), .ZN(n8820) );
  AOI22D1BWP30P140LVT U12863 ( .A1(i_data_bus[390]), .A2(n10387), .B1(
        i_data_bus[454]), .B2(n10388), .ZN(n8819) );
  ND2D1BWP30P140LVT U12864 ( .A1(n8820), .A2(n8819), .ZN(N10759) );
  AOI22D1BWP30P140LVT U12865 ( .A1(i_data_bus[461]), .A2(n10388), .B1(
        i_data_bus[493]), .B2(n10385), .ZN(n8822) );
  AOI22D1BWP30P140LVT U12866 ( .A1(i_data_bus[397]), .A2(n10387), .B1(
        i_data_bus[429]), .B2(n10386), .ZN(n8821) );
  ND2D1BWP30P140LVT U12867 ( .A1(n8822), .A2(n8821), .ZN(N10766) );
  INVD1BWP30P140LVT U12868 ( .I(inner_first_stage_valid_reg[62]), .ZN(n8828)
         );
  INVD1BWP30P140LVT U12869 ( .I(inner_first_stage_valid_reg[63]), .ZN(n8826)
         );
  INR4D0BWP30P140LVT U12870 ( .A1(n8825), .B1(inner_first_stage_valid_reg[56]), 
        .B2(inner_first_stage_valid_reg[58]), .B3(n8823), .ZN(n8834) );
  INR3D2BWP30P140LVT U12871 ( .A1(inner_first_stage_valid_reg[57]), .B1(
        inner_first_stage_valid_reg[61]), .B2(n8832), .ZN(n12296) );
  NR3D0P7BWP30P140LVT U12872 ( .A1(inner_first_stage_valid_reg[62]), .A2(
        inner_first_stage_valid_reg[63]), .A3(n11173), .ZN(n8830) );
  NR3D0P7BWP30P140LVT U12873 ( .A1(inner_first_stage_valid_reg[59]), .A2(
        inner_first_stage_valid_reg[57]), .A3(inner_first_stage_valid_reg[61]), 
        .ZN(n8829) );
  INR3D0BWP30P140LVT U12874 ( .A1(n8829), .B1(inner_first_stage_valid_reg[56]), 
        .B2(inner_first_stage_valid_reg[58]), .ZN(n8824) );
  NR4D0BWP30P140LVT U12875 ( .A1(n12296), .A2(n12295), .A3(n12297), .A4(n6211), 
        .ZN(n8836) );
  IND3D1BWP30P140LVT U12876 ( .A1(inner_first_stage_valid_reg[60]), .B1(n8830), 
        .B2(n8829), .ZN(n8831) );
  INR3D2BWP30P140LVT U12877 ( .A1(inner_first_stage_valid_reg[56]), .B1(
        inner_first_stage_valid_reg[58]), .B2(n8831), .ZN(n12294) );
  INR3D2BWP30P140LVT U12878 ( .A1(inner_first_stage_valid_reg[58]), .B1(
        inner_first_stage_valid_reg[56]), .B2(n8831), .ZN(n12293) );
  INR3D2BWP30P140LVT U12879 ( .A1(inner_first_stage_valid_reg[61]), .B1(
        inner_first_stage_valid_reg[57]), .B2(n8832), .ZN(n12292) );
  INR4D1BWP30P140LVT U12880 ( .A1(n8834), .B1(inner_first_stage_valid_reg[61]), 
        .B2(inner_first_stage_valid_reg[57]), .B3(n8833), .ZN(n12291) );
  NR4D0BWP30P140LVT U12881 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(n8835) );
  AOI22D1BWP30P140LVT U12882 ( .A1(i_data_bus[516]), .A2(n10006), .B1(
        i_data_bus[580]), .B2(n10013), .ZN(n8838) );
  AOI22D1BWP30P140LVT U12883 ( .A1(i_data_bus[548]), .A2(n10012), .B1(
        i_data_bus[612]), .B2(n10011), .ZN(n8837) );
  ND2D1BWP30P140LVT U12884 ( .A1(n8838), .A2(n8837), .ZN(N2673) );
  AOI22D1BWP30P140LVT U12885 ( .A1(i_data_bus[572]), .A2(n10012), .B1(
        i_data_bus[540]), .B2(n10006), .ZN(n8840) );
  AOI22D1BWP30P140LVT U12886 ( .A1(i_data_bus[604]), .A2(n10013), .B1(
        i_data_bus[636]), .B2(n10011), .ZN(n8839) );
  ND2D1BWP30P140LVT U12887 ( .A1(n8840), .A2(n8839), .ZN(N2697) );
  AOI22D1BWP30P140LVT U12888 ( .A1(i_data_bus[571]), .A2(n10012), .B1(
        i_data_bus[603]), .B2(n10013), .ZN(n8842) );
  AOI22D1BWP30P140LVT U12889 ( .A1(i_data_bus[539]), .A2(n10006), .B1(
        i_data_bus[635]), .B2(n10011), .ZN(n8841) );
  ND2D1BWP30P140LVT U12890 ( .A1(n8842), .A2(n8841), .ZN(N2696) );
  AOI22D1BWP30P140LVT U12891 ( .A1(i_data_bus[535]), .A2(n10006), .B1(
        i_data_bus[599]), .B2(n10013), .ZN(n8844) );
  AOI22D1BWP30P140LVT U12892 ( .A1(i_data_bus[567]), .A2(n10012), .B1(
        i_data_bus[631]), .B2(n10011), .ZN(n8843) );
  ND2D1BWP30P140LVT U12893 ( .A1(n8844), .A2(n8843), .ZN(N2692) );
  AOI22D1BWP30P140LVT U12894 ( .A1(i_data_bus[563]), .A2(n10012), .B1(
        i_data_bus[595]), .B2(n10013), .ZN(n8846) );
  AOI22D1BWP30P140LVT U12895 ( .A1(i_data_bus[531]), .A2(n10006), .B1(
        i_data_bus[627]), .B2(n10011), .ZN(n8845) );
  ND2D1BWP30P140LVT U12896 ( .A1(n8846), .A2(n8845), .ZN(N2688) );
  AOI22D1BWP30P140LVT U12897 ( .A1(i_data_bus[562]), .A2(n10012), .B1(
        i_data_bus[594]), .B2(n10013), .ZN(n8848) );
  AOI22D1BWP30P140LVT U12898 ( .A1(i_data_bus[530]), .A2(n10006), .B1(
        i_data_bus[626]), .B2(n10011), .ZN(n8847) );
  ND2D1BWP30P140LVT U12899 ( .A1(n8848), .A2(n8847), .ZN(N2687) );
  AOI22D1BWP30P140LVT U12900 ( .A1(i_data_bus[529]), .A2(n10006), .B1(
        i_data_bus[593]), .B2(n10013), .ZN(n8850) );
  AOI22D1BWP30P140LVT U12901 ( .A1(i_data_bus[561]), .A2(n10012), .B1(
        i_data_bus[625]), .B2(n10011), .ZN(n8849) );
  ND2D1BWP30P140LVT U12902 ( .A1(n8850), .A2(n8849), .ZN(N2686) );
  AOI22D1BWP30P140LVT U12903 ( .A1(i_data_bus[558]), .A2(n10012), .B1(
        i_data_bus[526]), .B2(n10006), .ZN(n8852) );
  AOI22D1BWP30P140LVT U12904 ( .A1(i_data_bus[590]), .A2(n10013), .B1(
        i_data_bus[622]), .B2(n10011), .ZN(n8851) );
  ND2D1BWP30P140LVT U12905 ( .A1(n8852), .A2(n8851), .ZN(N2683) );
  AOI22D1BWP30P140LVT U12906 ( .A1(i_data_bus[550]), .A2(n10012), .B1(
        i_data_bus[582]), .B2(n10013), .ZN(n8854) );
  AOI22D1BWP30P140LVT U12907 ( .A1(i_data_bus[518]), .A2(n10006), .B1(
        i_data_bus[614]), .B2(n10011), .ZN(n8853) );
  ND2D1BWP30P140LVT U12908 ( .A1(n8854), .A2(n8853), .ZN(N2675) );
  AOI22D1BWP30P140LVT U12909 ( .A1(i_data_bus[34]), .A2(n9791), .B1(
        i_data_bus[66]), .B2(n9790), .ZN(n8856) );
  AOI22D1BWP30P140LVT U12910 ( .A1(i_data_bus[98]), .A2(n9792), .B1(
        i_data_bus[2]), .B2(n6223), .ZN(n8855) );
  ND2D1BWP30P140LVT U12911 ( .A1(n8856), .A2(n8855), .ZN(N8745) );
  AOI22D1BWP30P140LVT U12912 ( .A1(i_data_bus[99]), .A2(n9792), .B1(
        i_data_bus[67]), .B2(n9790), .ZN(n8858) );
  AOI22D1BWP30P140LVT U12913 ( .A1(i_data_bus[35]), .A2(n9791), .B1(
        i_data_bus[3]), .B2(n6223), .ZN(n8857) );
  ND2D1BWP30P140LVT U12914 ( .A1(n8858), .A2(n8857), .ZN(N8746) );
  AOI22D1BWP30P140LVT U12915 ( .A1(i_data_bus[349]), .A2(n9731), .B1(
        i_data_bus[317]), .B2(n9732), .ZN(n8860) );
  AOI22D1BWP30P140LVT U12916 ( .A1(i_data_bus[381]), .A2(n9730), .B1(
        i_data_bus[285]), .B2(n6219), .ZN(n8859) );
  ND2D1BWP30P140LVT U12917 ( .A1(n8860), .A2(n8859), .ZN(N3756) );
  AOI22D1BWP30P140LVT U12918 ( .A1(i_data_bus[335]), .A2(n9755), .B1(
        i_data_bus[367]), .B2(n9757), .ZN(n8862) );
  AOI22D1BWP30P140LVT U12919 ( .A1(i_data_bus[303]), .A2(n9758), .B1(
        i_data_bus[271]), .B2(n9756), .ZN(n8861) );
  ND2D1BWP30P140LVT U12920 ( .A1(n8862), .A2(n8861), .ZN(N5232) );
  AOI22D1BWP30P140LVT U12921 ( .A1(i_data_bus[430]), .A2(n10405), .B1(
        i_data_bus[462]), .B2(n10408), .ZN(n8864) );
  AOI22D1BWP30P140LVT U12922 ( .A1(i_data_bus[398]), .A2(n10407), .B1(
        i_data_bus[494]), .B2(n10406), .ZN(n8863) );
  ND2D1BWP30P140LVT U12923 ( .A1(n8864), .A2(n8863), .ZN(N9405) );
  AOI22D1BWP30P140LVT U12924 ( .A1(i_data_bus[506]), .A2(n10406), .B1(
        i_data_bus[474]), .B2(n10408), .ZN(n8866) );
  AOI22D1BWP30P140LVT U12925 ( .A1(i_data_bus[410]), .A2(n10407), .B1(
        i_data_bus[442]), .B2(n10405), .ZN(n8865) );
  ND2D1BWP30P140LVT U12926 ( .A1(n8866), .A2(n8865), .ZN(N9417) );
  AOI22D1BWP30P140LVT U12927 ( .A1(i_data_bus[505]), .A2(n10406), .B1(
        i_data_bus[473]), .B2(n10408), .ZN(n8868) );
  AOI22D1BWP30P140LVT U12928 ( .A1(i_data_bus[409]), .A2(n10407), .B1(
        i_data_bus[441]), .B2(n10405), .ZN(n8867) );
  ND2D1BWP30P140LVT U12929 ( .A1(n8868), .A2(n8867), .ZN(N9416) );
  AOI22D1BWP30P140LVT U12930 ( .A1(i_data_bus[501]), .A2(n10406), .B1(
        i_data_bus[469]), .B2(n10408), .ZN(n8870) );
  AOI22D1BWP30P140LVT U12931 ( .A1(i_data_bus[405]), .A2(n10407), .B1(
        i_data_bus[437]), .B2(n10405), .ZN(n8869) );
  ND2D1BWP30P140LVT U12932 ( .A1(n8870), .A2(n8869), .ZN(N9412) );
  AOI22D1BWP30P140LVT U12933 ( .A1(i_data_bus[502]), .A2(n10406), .B1(
        i_data_bus[438]), .B2(n10405), .ZN(n8872) );
  AOI22D1BWP30P140LVT U12934 ( .A1(i_data_bus[406]), .A2(n10407), .B1(
        i_data_bus[470]), .B2(n10408), .ZN(n8871) );
  ND2D1BWP30P140LVT U12935 ( .A1(n8872), .A2(n8871), .ZN(N9413) );
  AOI22D1BWP30P140LVT U12936 ( .A1(i_data_bus[446]), .A2(n10405), .B1(
        i_data_bus[510]), .B2(n10406), .ZN(n8874) );
  AOI22D1BWP30P140LVT U12937 ( .A1(i_data_bus[414]), .A2(n10407), .B1(
        i_data_bus[478]), .B2(n10408), .ZN(n8873) );
  ND2D1BWP30P140LVT U12938 ( .A1(n8874), .A2(n8873), .ZN(N9421) );
  AOI22D1BWP30P140LVT U12939 ( .A1(i_data_bus[426]), .A2(n10405), .B1(
        i_data_bus[490]), .B2(n10406), .ZN(n8876) );
  AOI22D1BWP30P140LVT U12940 ( .A1(i_data_bus[394]), .A2(n10407), .B1(
        i_data_bus[458]), .B2(n10408), .ZN(n8875) );
  ND2D1BWP30P140LVT U12941 ( .A1(n8876), .A2(n8875), .ZN(N9401) );
  AOI22D1BWP30P140LVT U12942 ( .A1(i_data_bus[422]), .A2(n10405), .B1(
        i_data_bus[486]), .B2(n10406), .ZN(n8878) );
  AOI22D1BWP30P140LVT U12943 ( .A1(i_data_bus[390]), .A2(n10407), .B1(
        i_data_bus[454]), .B2(n10408), .ZN(n8877) );
  ND2D1BWP30P140LVT U12944 ( .A1(n8878), .A2(n8877), .ZN(N9397) );
  AOI22D1BWP30P140LVT U12945 ( .A1(i_data_bus[482]), .A2(n10406), .B1(
        i_data_bus[418]), .B2(n10405), .ZN(n8880) );
  AOI22D1BWP30P140LVT U12946 ( .A1(i_data_bus[386]), .A2(n10407), .B1(
        i_data_bus[450]), .B2(n10408), .ZN(n8879) );
  ND2D1BWP30P140LVT U12947 ( .A1(n8880), .A2(n8879), .ZN(N9393) );
  AOI22D1BWP30P140LVT U12948 ( .A1(i_data_bus[429]), .A2(n10405), .B1(
        i_data_bus[493]), .B2(n10406), .ZN(n8882) );
  AOI22D1BWP30P140LVT U12949 ( .A1(i_data_bus[397]), .A2(n10407), .B1(
        i_data_bus[461]), .B2(n10408), .ZN(n8881) );
  ND2D1BWP30P140LVT U12950 ( .A1(n8882), .A2(n8881), .ZN(N9404) );
  AOI22D1BWP30P140LVT U12951 ( .A1(i_data_bus[360]), .A2(n9773), .B1(
        i_data_bus[296]), .B2(n9775), .ZN(n8884) );
  AOI22D1BWP30P140LVT U12952 ( .A1(i_data_bus[328]), .A2(n9774), .B1(
        i_data_bus[264]), .B2(n6216), .ZN(n8883) );
  ND2D1BWP30P140LVT U12953 ( .A1(n8884), .A2(n8883), .ZN(N2501) );
  AOI22D1BWP30P140LVT U12954 ( .A1(i_data_bus[87]), .A2(n9790), .B1(
        i_data_bus[119]), .B2(n9792), .ZN(n8886) );
  AOI22D1BWP30P140LVT U12955 ( .A1(i_data_bus[55]), .A2(n9791), .B1(
        i_data_bus[23]), .B2(n6223), .ZN(n8885) );
  ND2D1BWP30P140LVT U12956 ( .A1(n8886), .A2(n8885), .ZN(N8766) );
  AOI22D1BWP30P140LVT U12957 ( .A1(i_data_bus[317]), .A2(n9843), .B1(
        i_data_bus[381]), .B2(n9845), .ZN(n8888) );
  AOI22D1BWP30P140LVT U12958 ( .A1(i_data_bus[349]), .A2(n9844), .B1(
        i_data_bus[285]), .B2(n9846), .ZN(n8887) );
  ND2D1BWP30P140LVT U12959 ( .A1(n8888), .A2(n8887), .ZN(N7970) );
  AOI22D1BWP30P140LVT U12960 ( .A1(i_data_bus[428]), .A2(n10427), .B1(
        i_data_bus[492]), .B2(n10428), .ZN(n8890) );
  AOI22D1BWP30P140LVT U12961 ( .A1(i_data_bus[396]), .A2(n10429), .B1(
        i_data_bus[460]), .B2(n10430), .ZN(n8889) );
  ND2D1BWP30P140LVT U12962 ( .A1(n8890), .A2(n8889), .ZN(N6679) );
  AOI22D1BWP30P140LVT U12963 ( .A1(i_data_bus[423]), .A2(n10427), .B1(
        i_data_bus[487]), .B2(n10428), .ZN(n8892) );
  AOI22D1BWP30P140LVT U12964 ( .A1(i_data_bus[391]), .A2(n10429), .B1(
        i_data_bus[455]), .B2(n10430), .ZN(n8891) );
  ND2D1BWP30P140LVT U12965 ( .A1(n8892), .A2(n8891), .ZN(N6674) );
  AOI22D1BWP30P140LVT U12966 ( .A1(i_data_bus[485]), .A2(n10428), .B1(
        i_data_bus[421]), .B2(n10427), .ZN(n8894) );
  AOI22D1BWP30P140LVT U12967 ( .A1(i_data_bus[389]), .A2(n10429), .B1(
        i_data_bus[453]), .B2(n10430), .ZN(n8893) );
  ND2D1BWP30P140LVT U12968 ( .A1(n8894), .A2(n8893), .ZN(N6672) );
  AOI22D1BWP30P140LVT U12969 ( .A1(i_data_bus[505]), .A2(n10428), .B1(
        i_data_bus[473]), .B2(n10430), .ZN(n8896) );
  AOI22D1BWP30P140LVT U12970 ( .A1(i_data_bus[409]), .A2(n10429), .B1(
        i_data_bus[441]), .B2(n10427), .ZN(n8895) );
  ND2D1BWP30P140LVT U12971 ( .A1(n8896), .A2(n8895), .ZN(N6692) );
  AOI22D1BWP30P140LVT U12972 ( .A1(i_data_bus[477]), .A2(n10430), .B1(
        i_data_bus[445]), .B2(n10427), .ZN(n8898) );
  AOI22D1BWP30P140LVT U12973 ( .A1(i_data_bus[413]), .A2(n10429), .B1(
        i_data_bus[509]), .B2(n10428), .ZN(n8897) );
  ND2D1BWP30P140LVT U12974 ( .A1(n8898), .A2(n8897), .ZN(N6696) );
  AOI22D1BWP30P140LVT U12975 ( .A1(i_data_bus[464]), .A2(n10430), .B1(
        i_data_bus[432]), .B2(n10427), .ZN(n8900) );
  AOI22D1BWP30P140LVT U12976 ( .A1(i_data_bus[400]), .A2(n10429), .B1(
        i_data_bus[496]), .B2(n10428), .ZN(n8899) );
  ND2D1BWP30P140LVT U12977 ( .A1(n8900), .A2(n8899), .ZN(N6683) );
  AOI22D1BWP30P140LVT U12978 ( .A1(i_data_bus[452]), .A2(n10430), .B1(
        i_data_bus[420]), .B2(n10427), .ZN(n8902) );
  AOI22D1BWP30P140LVT U12979 ( .A1(i_data_bus[388]), .A2(n10429), .B1(
        i_data_bus[484]), .B2(n10428), .ZN(n8901) );
  ND2D1BWP30P140LVT U12980 ( .A1(n8902), .A2(n8901), .ZN(N6671) );
  AOI22D1BWP30P140LVT U12981 ( .A1(i_data_bus[422]), .A2(n10427), .B1(
        i_data_bus[454]), .B2(n10430), .ZN(n8904) );
  AOI22D1BWP30P140LVT U12982 ( .A1(i_data_bus[390]), .A2(n10429), .B1(
        i_data_bus[486]), .B2(n10428), .ZN(n8903) );
  ND2D1BWP30P140LVT U12983 ( .A1(n8904), .A2(n8903), .ZN(N6673) );
  AOI22D1BWP30P140LVT U12984 ( .A1(i_data_bus[450]), .A2(n10430), .B1(
        i_data_bus[418]), .B2(n10427), .ZN(n8906) );
  AOI22D1BWP30P140LVT U12985 ( .A1(i_data_bus[386]), .A2(n10429), .B1(
        i_data_bus[482]), .B2(n10428), .ZN(n8905) );
  ND2D1BWP30P140LVT U12986 ( .A1(n8906), .A2(n8905), .ZN(N6669) );
  AOI22D1BWP30P140LVT U12987 ( .A1(i_data_bus[340]), .A2(n9879), .B1(
        i_data_bus[308]), .B2(n9878), .ZN(n8908) );
  AOI22D1BWP30P140LVT U12988 ( .A1(i_data_bus[372]), .A2(n9877), .B1(
        i_data_bus[276]), .B2(n6217), .ZN(n8907) );
  ND2D1BWP30P140LVT U12989 ( .A1(n8908), .A2(n8907), .ZN(N10685) );
  AOI22D1BWP30P140LVT U12990 ( .A1(i_data_bus[378]), .A2(n9877), .B1(
        i_data_bus[314]), .B2(n9878), .ZN(n8910) );
  AOI22D1BWP30P140LVT U12991 ( .A1(i_data_bus[346]), .A2(n9879), .B1(
        i_data_bus[282]), .B2(n6217), .ZN(n8909) );
  ND2D1BWP30P140LVT U12992 ( .A1(n8910), .A2(n8909), .ZN(N10691) );
  AOI22D1BWP30P140LVT U12993 ( .A1(i_data_bus[363]), .A2(n9877), .B1(
        i_data_bus[299]), .B2(n9878), .ZN(n8912) );
  AOI22D1BWP30P140LVT U12994 ( .A1(i_data_bus[331]), .A2(n9879), .B1(
        i_data_bus[267]), .B2(n6217), .ZN(n8911) );
  ND2D1BWP30P140LVT U12995 ( .A1(n8912), .A2(n8911), .ZN(N10676) );
  AOI22D1BWP30P140LVT U12996 ( .A1(i_data_bus[529]), .A2(n10272), .B1(
        i_data_bus[593]), .B2(n10269), .ZN(n8914) );
  AOI22D1BWP30P140LVT U12997 ( .A1(i_data_bus[561]), .A2(n10271), .B1(
        i_data_bus[625]), .B2(n10270), .ZN(n8913) );
  ND2D1BWP30P140LVT U12998 ( .A1(n8914), .A2(n8913), .ZN(N8134) );
  AOI22D1BWP30P140LVT U12999 ( .A1(i_data_bus[590]), .A2(n10269), .B1(
        i_data_bus[526]), .B2(n10272), .ZN(n8916) );
  AOI22D1BWP30P140LVT U13000 ( .A1(i_data_bus[558]), .A2(n10271), .B1(
        i_data_bus[622]), .B2(n10270), .ZN(n8915) );
  ND2D1BWP30P140LVT U13001 ( .A1(n8916), .A2(n8915), .ZN(N8131) );
  AOI22D1BWP30P140LVT U13002 ( .A1(i_data_bus[516]), .A2(n10272), .B1(
        i_data_bus[580]), .B2(n10269), .ZN(n8918) );
  AOI22D1BWP30P140LVT U13003 ( .A1(i_data_bus[548]), .A2(n10271), .B1(
        i_data_bus[612]), .B2(n10270), .ZN(n8917) );
  ND2D1BWP30P140LVT U13004 ( .A1(n8918), .A2(n8917), .ZN(N8121) );
  AOI22D1BWP30P140LVT U13005 ( .A1(i_data_bus[578]), .A2(n9936), .B1(
        i_data_bus[546]), .B2(n9935), .ZN(n8920) );
  AOI22D1BWP30P140LVT U13006 ( .A1(i_data_bus[610]), .A2(n9933), .B1(
        i_data_bus[514]), .B2(n9934), .ZN(n8919) );
  ND2D1BWP30P140LVT U13007 ( .A1(n8920), .A2(n8919), .ZN(N5395) );
  AOI22D1BWP30P140LVT U13008 ( .A1(i_data_bus[639]), .A2(n9933), .B1(
        i_data_bus[575]), .B2(n9935), .ZN(n8922) );
  AOI22D1BWP30P140LVT U13009 ( .A1(i_data_bus[607]), .A2(n9936), .B1(
        i_data_bus[543]), .B2(n9934), .ZN(n8921) );
  ND2D1BWP30P140LVT U13010 ( .A1(n8922), .A2(n8921), .ZN(N5424) );
  AOI22D1BWP30P140LVT U13011 ( .A1(i_data_bus[616]), .A2(n9933), .B1(
        i_data_bus[552]), .B2(n9935), .ZN(n8924) );
  AOI22D1BWP30P140LVT U13012 ( .A1(i_data_bus[584]), .A2(n9936), .B1(
        i_data_bus[520]), .B2(n9934), .ZN(n8923) );
  ND2D1BWP30P140LVT U13013 ( .A1(n8924), .A2(n8923), .ZN(N5401) );
  AOI22D1BWP30P140LVT U13014 ( .A1(i_data_bus[74]), .A2(n9914), .B1(
        i_data_bus[42]), .B2(n9916), .ZN(n8926) );
  AOI22D1BWP30P140LVT U13015 ( .A1(i_data_bus[106]), .A2(n9915), .B1(
        i_data_bus[10]), .B2(n6218), .ZN(n8925) );
  ND2D1BWP30P140LVT U13016 ( .A1(n8926), .A2(n8925), .ZN(N3305) );
  AOI22D1BWP30P140LVT U13017 ( .A1(i_data_bus[95]), .A2(n9914), .B1(
        i_data_bus[63]), .B2(n9916), .ZN(n8928) );
  AOI22D1BWP30P140LVT U13018 ( .A1(i_data_bus[127]), .A2(n9915), .B1(
        i_data_bus[31]), .B2(n6218), .ZN(n8927) );
  ND2D1BWP30P140LVT U13019 ( .A1(n8928), .A2(n8927), .ZN(N3326) );
  INR4D1BWP30P140LVT U13020 ( .A1(i_cmd[20]), .B1(i_cmd[4]), .B2(n10632), .B3(
        n11046), .ZN(n10095) );
  NR4D1BWP30P140LVT U13021 ( .A1(i_cmd[12]), .A2(n8929), .A3(n10630), .A4(
        n11049), .ZN(n10098) );
  AOI22D1BWP30P140LVT U13022 ( .A1(i_data_bus[82]), .A2(n10095), .B1(
        i_data_bus[114]), .B2(n10098), .ZN(n8931) );
  NR4D1BWP30P140LVT U13023 ( .A1(i_cmd[28]), .A2(n8929), .A3(n10634), .A4(
        n11048), .ZN(n10097) );
  NR3D0P7BWP30P140LVT U13024 ( .A1(i_cmd[20]), .A2(i_cmd[28]), .A3(i_cmd[12]), 
        .ZN(n11045) );
  AOI22D1BWP30P140LVT U13025 ( .A1(i_data_bus[50]), .A2(n10097), .B1(
        i_data_bus[18]), .B2(n10096), .ZN(n8930) );
  ND2D1BWP30P140LVT U13026 ( .A1(n8931), .A2(n8930), .ZN(N6037) );
  AOI22D1BWP30P140LVT U13027 ( .A1(i_data_bus[73]), .A2(n9976), .B1(
        i_data_bus[105]), .B2(n9978), .ZN(n8933) );
  AOI22D1BWP30P140LVT U13028 ( .A1(i_data_bus[41]), .A2(n9977), .B1(
        i_data_bus[9]), .B2(n9969), .ZN(n8932) );
  ND2D1BWP30P140LVT U13029 ( .A1(n8933), .A2(n8932), .ZN(N2326) );
  AOI22D1BWP30P140LVT U13030 ( .A1(i_data_bus[118]), .A2(n9915), .B1(
        i_data_bus[54]), .B2(n9916), .ZN(n8935) );
  AOI22D1BWP30P140LVT U13031 ( .A1(i_data_bus[86]), .A2(n9914), .B1(
        i_data_bus[22]), .B2(n6218), .ZN(n8934) );
  ND2D1BWP30P140LVT U13032 ( .A1(n8935), .A2(n8934), .ZN(N3317) );
  AOI22D1BWP30P140LVT U13033 ( .A1(i_data_bus[61]), .A2(n9977), .B1(
        i_data_bus[125]), .B2(n9978), .ZN(n8937) );
  AOI22D1BWP30P140LVT U13034 ( .A1(i_data_bus[93]), .A2(n9976), .B1(
        i_data_bus[29]), .B2(n9969), .ZN(n8936) );
  ND2D1BWP30P140LVT U13035 ( .A1(n8937), .A2(n8936), .ZN(N2346) );
  AOI22D1BWP30P140LVT U13036 ( .A1(i_data_bus[50]), .A2(n9977), .B1(
        i_data_bus[114]), .B2(n9978), .ZN(n8939) );
  AOI22D1BWP30P140LVT U13037 ( .A1(i_data_bus[82]), .A2(n9976), .B1(
        i_data_bus[18]), .B2(n9969), .ZN(n8938) );
  ND2D1BWP30P140LVT U13038 ( .A1(n8939), .A2(n8938), .ZN(N2335) );
  AOI22D1BWP30P140LVT U13039 ( .A1(i_data_bus[629]), .A2(n9933), .B1(
        i_data_bus[565]), .B2(n9935), .ZN(n8941) );
  AOI22D1BWP30P140LVT U13040 ( .A1(i_data_bus[533]), .A2(n9934), .B1(
        i_data_bus[597]), .B2(n9936), .ZN(n8940) );
  ND2D1BWP30P140LVT U13041 ( .A1(n8941), .A2(n8940), .ZN(N5414) );
  AOI22D1BWP30P140LVT U13042 ( .A1(i_data_bus[623]), .A2(n9933), .B1(
        i_data_bus[559]), .B2(n9935), .ZN(n8943) );
  AOI22D1BWP30P140LVT U13043 ( .A1(i_data_bus[527]), .A2(n9934), .B1(
        i_data_bus[591]), .B2(n9936), .ZN(n8942) );
  ND2D1BWP30P140LVT U13044 ( .A1(n8943), .A2(n8942), .ZN(N5408) );
  AOI22D1BWP30P140LVT U13045 ( .A1(i_data_bus[607]), .A2(n10001), .B1(
        i_data_bus[575]), .B2(n10002), .ZN(n8945) );
  AOI22D1BWP30P140LVT U13046 ( .A1(i_data_bus[639]), .A2(n10003), .B1(
        i_data_bus[543]), .B2(n6222), .ZN(n8944) );
  ND2D1BWP30P140LVT U13047 ( .A1(n8945), .A2(n8944), .ZN(N4190) );
  AOI22D1BWP30P140LVT U13048 ( .A1(i_data_bus[628]), .A2(n10003), .B1(
        i_data_bus[564]), .B2(n10002), .ZN(n8947) );
  AOI22D1BWP30P140LVT U13049 ( .A1(i_data_bus[596]), .A2(n10001), .B1(
        i_data_bus[532]), .B2(n6222), .ZN(n8946) );
  ND2D1BWP30P140LVT U13050 ( .A1(n8947), .A2(n8946), .ZN(N4179) );
  AOI22D1BWP30P140LVT U13051 ( .A1(i_data_bus[616]), .A2(n10003), .B1(
        i_data_bus[552]), .B2(n10002), .ZN(n8949) );
  AOI22D1BWP30P140LVT U13052 ( .A1(i_data_bus[584]), .A2(n10001), .B1(
        i_data_bus[520]), .B2(n6222), .ZN(n8948) );
  ND2D1BWP30P140LVT U13053 ( .A1(n8949), .A2(n8948), .ZN(N4167) );
  AOI22D1BWP30P140LVT U13054 ( .A1(i_data_bus[639]), .A2(n10011), .B1(
        i_data_bus[575]), .B2(n10012), .ZN(n8951) );
  AOI22D1BWP30P140LVT U13055 ( .A1(i_data_bus[607]), .A2(n10013), .B1(
        i_data_bus[543]), .B2(n10006), .ZN(n8950) );
  ND2D1BWP30P140LVT U13056 ( .A1(n8951), .A2(n8950), .ZN(N2700) );
  AOI22D1BWP30P140LVT U13057 ( .A1(i_data_bus[522]), .A2(n6222), .B1(
        i_data_bus[554]), .B2(n10002), .ZN(n8953) );
  AOI22D1BWP30P140LVT U13058 ( .A1(i_data_bus[586]), .A2(n10001), .B1(
        i_data_bus[618]), .B2(n10003), .ZN(n8952) );
  ND2D1BWP30P140LVT U13059 ( .A1(n8953), .A2(n8952), .ZN(N4169) );
  AOI22D1BWP30P140LVT U13060 ( .A1(i_data_bus[512]), .A2(n6222), .B1(
        i_data_bus[544]), .B2(n10002), .ZN(n8955) );
  AOI22D1BWP30P140LVT U13061 ( .A1(i_data_bus[576]), .A2(n10001), .B1(
        i_data_bus[608]), .B2(n10003), .ZN(n8954) );
  ND2D1BWP30P140LVT U13062 ( .A1(n8955), .A2(n8954), .ZN(N4159) );
  AOI22D1BWP30P140LVT U13063 ( .A1(i_data_bus[590]), .A2(n10001), .B1(
        i_data_bus[558]), .B2(n10002), .ZN(n8957) );
  AOI22D1BWP30P140LVT U13064 ( .A1(i_data_bus[526]), .A2(n6222), .B1(
        i_data_bus[622]), .B2(n10003), .ZN(n8956) );
  ND2D1BWP30P140LVT U13065 ( .A1(n8957), .A2(n8956), .ZN(N4173) );
  AOI22D1BWP30P140LVT U13066 ( .A1(i_data_bus[522]), .A2(n10006), .B1(
        i_data_bus[554]), .B2(n10012), .ZN(n8959) );
  AOI22D1BWP30P140LVT U13067 ( .A1(i_data_bus[586]), .A2(n10013), .B1(
        i_data_bus[618]), .B2(n10011), .ZN(n8958) );
  ND2D1BWP30P140LVT U13068 ( .A1(n8959), .A2(n8958), .ZN(N2679) );
  AOI22D1BWP30P140LVT U13069 ( .A1(i_data_bus[581]), .A2(n10013), .B1(
        i_data_bus[549]), .B2(n10012), .ZN(n8961) );
  AOI22D1BWP30P140LVT U13070 ( .A1(i_data_bus[517]), .A2(n10006), .B1(
        i_data_bus[613]), .B2(n10011), .ZN(n8960) );
  ND2D1BWP30P140LVT U13071 ( .A1(n8961), .A2(n8960), .ZN(N2674) );
  AOI22D1BWP30P140LVT U13072 ( .A1(i_data_bus[514]), .A2(n10006), .B1(
        i_data_bus[546]), .B2(n10012), .ZN(n8963) );
  AOI22D1BWP30P140LVT U13073 ( .A1(i_data_bus[578]), .A2(n10013), .B1(
        i_data_bus[610]), .B2(n10011), .ZN(n8962) );
  ND2D1BWP30P140LVT U13074 ( .A1(n8963), .A2(n8962), .ZN(N2671) );
  AOI22D1BWP30P140LVT U13075 ( .A1(i_data_bus[531]), .A2(n6222), .B1(
        i_data_bus[563]), .B2(n10002), .ZN(n8965) );
  AOI22D1BWP30P140LVT U13076 ( .A1(i_data_bus[627]), .A2(n10003), .B1(
        i_data_bus[595]), .B2(n10001), .ZN(n8964) );
  ND2D1BWP30P140LVT U13077 ( .A1(n8965), .A2(n8964), .ZN(N4178) );
  AOI22D1BWP30P140LVT U13078 ( .A1(i_data_bus[623]), .A2(n10003), .B1(
        i_data_bus[559]), .B2(n10002), .ZN(n8967) );
  AOI22D1BWP30P140LVT U13079 ( .A1(i_data_bus[527]), .A2(n6222), .B1(
        i_data_bus[591]), .B2(n10001), .ZN(n8966) );
  ND2D1BWP30P140LVT U13080 ( .A1(n8967), .A2(n8966), .ZN(N4174) );
  AOI22D1BWP30P140LVT U13081 ( .A1(i_data_bus[637]), .A2(n10011), .B1(
        i_data_bus[573]), .B2(n10012), .ZN(n8969) );
  AOI22D1BWP30P140LVT U13082 ( .A1(i_data_bus[541]), .A2(n10006), .B1(
        i_data_bus[605]), .B2(n10013), .ZN(n8968) );
  ND2D1BWP30P140LVT U13083 ( .A1(n8969), .A2(n8968), .ZN(N2698) );
  AOI22D1BWP30P140LVT U13084 ( .A1(i_data_bus[623]), .A2(n10011), .B1(
        i_data_bus[559]), .B2(n10012), .ZN(n8971) );
  AOI22D1BWP30P140LVT U13085 ( .A1(i_data_bus[527]), .A2(n10006), .B1(
        i_data_bus[591]), .B2(n10013), .ZN(n8970) );
  ND2D1BWP30P140LVT U13086 ( .A1(n8971), .A2(n8970), .ZN(N2684) );
  AOI22D1BWP30P140LVT U13087 ( .A1(i_data_bus[525]), .A2(n10006), .B1(
        i_data_bus[557]), .B2(n10012), .ZN(n8973) );
  AOI22D1BWP30P140LVT U13088 ( .A1(i_data_bus[621]), .A2(n10011), .B1(
        i_data_bus[589]), .B2(n10013), .ZN(n8972) );
  ND2D1BWP30P140LVT U13089 ( .A1(n8973), .A2(n8972), .ZN(N2682) );
  AOI22D1BWP30P140LVT U13090 ( .A1(i_data_bus[532]), .A2(n10006), .B1(
        i_data_bus[564]), .B2(n10012), .ZN(n8975) );
  AOI22D1BWP30P140LVT U13091 ( .A1(i_data_bus[628]), .A2(n10011), .B1(
        i_data_bus[596]), .B2(n10013), .ZN(n8974) );
  ND2D1BWP30P140LVT U13092 ( .A1(n8975), .A2(n8974), .ZN(N2689) );
  AOI22D1BWP30P140LVT U13093 ( .A1(i_data_bus[337]), .A2(n10054), .B1(
        i_data_bus[305]), .B2(n10053), .ZN(n8977) );
  AOI22D1BWP30P140LVT U13094 ( .A1(i_data_bus[369]), .A2(n10051), .B1(
        i_data_bus[273]), .B2(n10052), .ZN(n8976) );
  ND2D1BWP30P140LVT U13095 ( .A1(n8977), .A2(n8976), .ZN(N6468) );
  AOI22D1BWP30P140LVT U13096 ( .A1(i_data_bus[349]), .A2(n10054), .B1(
        i_data_bus[317]), .B2(n10053), .ZN(n8979) );
  AOI22D1BWP30P140LVT U13097 ( .A1(i_data_bus[381]), .A2(n10051), .B1(
        i_data_bus[285]), .B2(n10052), .ZN(n8978) );
  ND2D1BWP30P140LVT U13098 ( .A1(n8979), .A2(n8978), .ZN(N6480) );
  AOI22D1BWP30P140LVT U13099 ( .A1(i_data_bus[197]), .A2(n10033), .B1(
        i_data_bus[165]), .B2(n10034), .ZN(n8981) );
  AOI22D1BWP30P140LVT U13100 ( .A1(i_data_bus[229]), .A2(n10035), .B1(
        i_data_bus[133]), .B2(n10026), .ZN(n8980) );
  ND2D1BWP30P140LVT U13101 ( .A1(n8981), .A2(n8980), .ZN(N3516) );
  AOI22D1BWP30P140LVT U13102 ( .A1(i_data_bus[223]), .A2(n10039), .B1(
        i_data_bus[191]), .B2(n10040), .ZN(n8983) );
  AOI22D1BWP30P140LVT U13103 ( .A1(i_data_bus[255]), .A2(n10038), .B1(
        i_data_bus[159]), .B2(n9318), .ZN(n8982) );
  ND2D1BWP30P140LVT U13104 ( .A1(n8983), .A2(n8982), .ZN(N8990) );
  AOI22D1BWP30P140LVT U13105 ( .A1(i_data_bus[222]), .A2(n10039), .B1(
        i_data_bus[190]), .B2(n10040), .ZN(n8985) );
  AOI22D1BWP30P140LVT U13106 ( .A1(i_data_bus[254]), .A2(n10038), .B1(
        i_data_bus[158]), .B2(n9318), .ZN(n8984) );
  ND2D1BWP30P140LVT U13107 ( .A1(n8985), .A2(n8984), .ZN(N8989) );
  AOI22D1BWP30P140LVT U13108 ( .A1(i_data_bus[212]), .A2(n10039), .B1(
        i_data_bus[180]), .B2(n10040), .ZN(n8987) );
  AOI22D1BWP30P140LVT U13109 ( .A1(i_data_bus[244]), .A2(n10038), .B1(
        i_data_bus[148]), .B2(n9318), .ZN(n8986) );
  ND2D1BWP30P140LVT U13110 ( .A1(n8987), .A2(n8986), .ZN(N8979) );
  AOI22D1BWP30P140LVT U13111 ( .A1(i_data_bus[205]), .A2(n10039), .B1(
        i_data_bus[173]), .B2(n10040), .ZN(n8989) );
  AOI22D1BWP30P140LVT U13112 ( .A1(i_data_bus[237]), .A2(n10038), .B1(
        i_data_bus[141]), .B2(n9318), .ZN(n8988) );
  ND2D1BWP30P140LVT U13113 ( .A1(n8989), .A2(n8988), .ZN(N8972) );
  AOI22D1BWP30P140LVT U13114 ( .A1(i_data_bus[76]), .A2(n10095), .B1(
        i_data_bus[44]), .B2(n10097), .ZN(n8991) );
  AOI22D1BWP30P140LVT U13115 ( .A1(i_data_bus[108]), .A2(n10098), .B1(
        i_data_bus[12]), .B2(n10096), .ZN(n8990) );
  ND2D1BWP30P140LVT U13116 ( .A1(n8991), .A2(n8990), .ZN(N6031) );
  AOI22D1BWP30P140LVT U13117 ( .A1(i_data_bus[74]), .A2(n10095), .B1(
        i_data_bus[42]), .B2(n10097), .ZN(n8993) );
  AOI22D1BWP30P140LVT U13118 ( .A1(i_data_bus[106]), .A2(n10098), .B1(
        i_data_bus[10]), .B2(n10096), .ZN(n8992) );
  ND2D1BWP30P140LVT U13119 ( .A1(n8993), .A2(n8992), .ZN(N6029) );
  AOI22D1BWP30P140LVT U13120 ( .A1(i_data_bus[93]), .A2(n10086), .B1(
        i_data_bus[61]), .B2(n10087), .ZN(n8995) );
  AOI22D1BWP30P140LVT U13121 ( .A1(i_data_bus[125]), .A2(n10085), .B1(
        i_data_bus[29]), .B2(n10088), .ZN(n8994) );
  ND2D1BWP30P140LVT U13122 ( .A1(n8995), .A2(n8994), .ZN(N5070) );
  AOI22D1BWP30P140LVT U13123 ( .A1(i_data_bus[249]), .A2(n10038), .B1(
        i_data_bus[185]), .B2(n10040), .ZN(n8997) );
  AOI22D1BWP30P140LVT U13124 ( .A1(i_data_bus[217]), .A2(n10039), .B1(
        i_data_bus[153]), .B2(n9318), .ZN(n8996) );
  ND2D1BWP30P140LVT U13125 ( .A1(n8997), .A2(n8996), .ZN(N8984) );
  AOI22D1BWP30P140LVT U13126 ( .A1(i_data_bus[363]), .A2(n10051), .B1(
        i_data_bus[299]), .B2(n10053), .ZN(n8999) );
  AOI22D1BWP30P140LVT U13127 ( .A1(i_data_bus[331]), .A2(n10054), .B1(
        i_data_bus[267]), .B2(n10052), .ZN(n8998) );
  ND2D1BWP30P140LVT U13128 ( .A1(n8999), .A2(n8998), .ZN(N6462) );
  AOI22D1BWP30P140LVT U13129 ( .A1(i_data_bus[118]), .A2(n10098), .B1(
        i_data_bus[54]), .B2(n10097), .ZN(n9001) );
  AOI22D1BWP30P140LVT U13130 ( .A1(i_data_bus[86]), .A2(n10095), .B1(
        i_data_bus[22]), .B2(n10096), .ZN(n9000) );
  ND2D1BWP30P140LVT U13131 ( .A1(n9001), .A2(n9000), .ZN(N6041) );
  AOI22D1BWP30P140LVT U13132 ( .A1(i_data_bus[93]), .A2(n10115), .B1(
        i_data_bus[125]), .B2(n10117), .ZN(n9003) );
  AOI22D1BWP30P140LVT U13133 ( .A1(i_data_bus[61]), .A2(n10118), .B1(
        i_data_bus[29]), .B2(n10116), .ZN(n9002) );
  ND2D1BWP30P140LVT U13134 ( .A1(n9003), .A2(n9002), .ZN(N7794) );
  AOI22D1BWP30P140LVT U13135 ( .A1(i_data_bus[87]), .A2(n10115), .B1(
        i_data_bus[119]), .B2(n10117), .ZN(n9005) );
  AOI22D1BWP30P140LVT U13136 ( .A1(i_data_bus[55]), .A2(n10118), .B1(
        i_data_bus[23]), .B2(n10116), .ZN(n9004) );
  ND2D1BWP30P140LVT U13137 ( .A1(n9005), .A2(n9004), .ZN(N7788) );
  AOI22D1BWP30P140LVT U13138 ( .A1(i_data_bus[127]), .A2(n10085), .B1(
        i_data_bus[63]), .B2(n10087), .ZN(n9007) );
  AOI22D1BWP30P140LVT U13139 ( .A1(i_data_bus[95]), .A2(n10086), .B1(
        i_data_bus[31]), .B2(n10088), .ZN(n9006) );
  ND2D1BWP30P140LVT U13140 ( .A1(n9007), .A2(n9006), .ZN(N5072) );
  AOI22D1BWP30P140LVT U13141 ( .A1(i_data_bus[216]), .A2(n10033), .B1(
        i_data_bus[184]), .B2(n10034), .ZN(n9009) );
  AOI22D1BWP30P140LVT U13142 ( .A1(i_data_bus[152]), .A2(n10026), .B1(
        i_data_bus[248]), .B2(n10035), .ZN(n9008) );
  ND2D1BWP30P140LVT U13143 ( .A1(n9009), .A2(n9008), .ZN(N3535) );
  AOI22D1BWP30P140LVT U13144 ( .A1(i_data_bus[215]), .A2(n10033), .B1(
        i_data_bus[183]), .B2(n10034), .ZN(n9011) );
  AOI22D1BWP30P140LVT U13145 ( .A1(i_data_bus[151]), .A2(n10026), .B1(
        i_data_bus[247]), .B2(n10035), .ZN(n9010) );
  ND2D1BWP30P140LVT U13146 ( .A1(n9011), .A2(n9010), .ZN(N3534) );
  AOI22D1BWP30P140LVT U13147 ( .A1(i_data_bus[206]), .A2(n10033), .B1(
        i_data_bus[174]), .B2(n10034), .ZN(n9013) );
  AOI22D1BWP30P140LVT U13148 ( .A1(i_data_bus[142]), .A2(n10026), .B1(
        i_data_bus[238]), .B2(n10035), .ZN(n9012) );
  ND2D1BWP30P140LVT U13149 ( .A1(n9013), .A2(n9012), .ZN(N3525) );
  AOI22D1BWP30P140LVT U13150 ( .A1(i_data_bus[216]), .A2(n10039), .B1(
        i_data_bus[184]), .B2(n10040), .ZN(n9015) );
  AOI22D1BWP30P140LVT U13151 ( .A1(i_data_bus[152]), .A2(n9318), .B1(
        i_data_bus[248]), .B2(n10038), .ZN(n9014) );
  ND2D1BWP30P140LVT U13152 ( .A1(n9015), .A2(n9014), .ZN(N8983) );
  AOI22D1BWP30P140LVT U13153 ( .A1(i_data_bus[214]), .A2(n10039), .B1(
        i_data_bus[182]), .B2(n10040), .ZN(n9017) );
  AOI22D1BWP30P140LVT U13154 ( .A1(i_data_bus[150]), .A2(n9318), .B1(
        i_data_bus[246]), .B2(n10038), .ZN(n9016) );
  ND2D1BWP30P140LVT U13155 ( .A1(n9017), .A2(n9016), .ZN(N8981) );
  AOI22D1BWP30P140LVT U13156 ( .A1(i_data_bus[146]), .A2(n9318), .B1(
        i_data_bus[178]), .B2(n10040), .ZN(n9019) );
  AOI22D1BWP30P140LVT U13157 ( .A1(i_data_bus[210]), .A2(n10039), .B1(
        i_data_bus[242]), .B2(n10038), .ZN(n9018) );
  ND2D1BWP30P140LVT U13158 ( .A1(n9019), .A2(n9018), .ZN(N8977) );
  AOI22D1BWP30P140LVT U13159 ( .A1(i_data_bus[133]), .A2(n9318), .B1(
        i_data_bus[165]), .B2(n10040), .ZN(n9021) );
  AOI22D1BWP30P140LVT U13160 ( .A1(i_data_bus[197]), .A2(n10039), .B1(
        i_data_bus[229]), .B2(n10038), .ZN(n9020) );
  ND2D1BWP30P140LVT U13161 ( .A1(n9021), .A2(n9020), .ZN(N8964) );
  AOI22D1BWP30P140LVT U13162 ( .A1(i_data_bus[154]), .A2(n9318), .B1(
        i_data_bus[186]), .B2(n10040), .ZN(n9023) );
  AOI22D1BWP30P140LVT U13163 ( .A1(i_data_bus[218]), .A2(n10039), .B1(
        i_data_bus[250]), .B2(n10038), .ZN(n9022) );
  ND2D1BWP30P140LVT U13164 ( .A1(n9023), .A2(n9022), .ZN(N8985) );
  AOI22D1BWP30P140LVT U13165 ( .A1(i_data_bus[266]), .A2(n6217), .B1(
        i_data_bus[330]), .B2(n9879), .ZN(n9025) );
  AOI22D1BWP30P140LVT U13166 ( .A1(i_data_bus[298]), .A2(n9878), .B1(
        i_data_bus[362]), .B2(n9877), .ZN(n9024) );
  ND2D1BWP30P140LVT U13167 ( .A1(n9025), .A2(n9024), .ZN(N10675) );
  AOI22D1BWP30P140LVT U13168 ( .A1(i_data_bus[332]), .A2(n9879), .B1(
        i_data_bus[300]), .B2(n9878), .ZN(n9027) );
  AOI22D1BWP30P140LVT U13169 ( .A1(i_data_bus[268]), .A2(n6217), .B1(
        i_data_bus[364]), .B2(n9877), .ZN(n9026) );
  ND2D1BWP30P140LVT U13170 ( .A1(n9027), .A2(n9026), .ZN(N10677) );
  AOI22D1BWP30P140LVT U13171 ( .A1(i_data_bus[302]), .A2(n9878), .B1(
        i_data_bus[334]), .B2(n9879), .ZN(n9029) );
  AOI22D1BWP30P140LVT U13172 ( .A1(i_data_bus[270]), .A2(n6217), .B1(
        i_data_bus[366]), .B2(n9877), .ZN(n9028) );
  ND2D1BWP30P140LVT U13173 ( .A1(n9029), .A2(n9028), .ZN(N10679) );
  AOI22D1BWP30P140LVT U13174 ( .A1(i_data_bus[286]), .A2(n6227), .B1(
        i_data_bus[318]), .B2(n10276), .ZN(n9031) );
  AOI22D1BWP30P140LVT U13175 ( .A1(i_data_bus[350]), .A2(n10275), .B1(
        i_data_bus[382]), .B2(n10277), .ZN(n9030) );
  ND2D1BWP30P140LVT U13176 ( .A1(n9031), .A2(n9030), .ZN(N9205) );
  AOI22D1BWP30P140LVT U13177 ( .A1(i_data_bus[274]), .A2(n6227), .B1(
        i_data_bus[306]), .B2(n10276), .ZN(n9033) );
  AOI22D1BWP30P140LVT U13178 ( .A1(i_data_bus[338]), .A2(n10275), .B1(
        i_data_bus[370]), .B2(n10277), .ZN(n9032) );
  ND2D1BWP30P140LVT U13179 ( .A1(n9033), .A2(n9032), .ZN(N9193) );
  AOI22D1BWP30P140LVT U13180 ( .A1(i_data_bus[302]), .A2(n10276), .B1(
        i_data_bus[334]), .B2(n10275), .ZN(n9035) );
  AOI22D1BWP30P140LVT U13181 ( .A1(i_data_bus[270]), .A2(n6227), .B1(
        i_data_bus[366]), .B2(n10277), .ZN(n9034) );
  ND2D1BWP30P140LVT U13182 ( .A1(n9035), .A2(n9034), .ZN(N9189) );
  AOI22D1BWP30P140LVT U13183 ( .A1(i_data_bus[266]), .A2(n6227), .B1(
        i_data_bus[298]), .B2(n10276), .ZN(n9037) );
  AOI22D1BWP30P140LVT U13184 ( .A1(i_data_bus[330]), .A2(n10275), .B1(
        i_data_bus[362]), .B2(n10277), .ZN(n9036) );
  ND2D1BWP30P140LVT U13185 ( .A1(n9037), .A2(n9036), .ZN(N9185) );
  AOI22D1BWP30P140LVT U13186 ( .A1(i_data_bus[256]), .A2(n6227), .B1(
        i_data_bus[320]), .B2(n10275), .ZN(n9039) );
  AOI22D1BWP30P140LVT U13187 ( .A1(i_data_bus[288]), .A2(n10276), .B1(
        i_data_bus[352]), .B2(n10277), .ZN(n9038) );
  ND2D1BWP30P140LVT U13188 ( .A1(n9039), .A2(n9038), .ZN(N9175) );
  AOI22D1BWP30P140LVT U13189 ( .A1(i_data_bus[311]), .A2(n9878), .B1(
        i_data_bus[343]), .B2(n9879), .ZN(n9041) );
  AOI22D1BWP30P140LVT U13190 ( .A1(i_data_bus[279]), .A2(n6217), .B1(
        i_data_bus[375]), .B2(n9877), .ZN(n9040) );
  ND2D1BWP30P140LVT U13191 ( .A1(n9041), .A2(n9040), .ZN(N10688) );
  AOI22D1BWP30P140LVT U13192 ( .A1(i_data_bus[350]), .A2(n9879), .B1(
        i_data_bus[318]), .B2(n9878), .ZN(n9043) );
  AOI22D1BWP30P140LVT U13193 ( .A1(i_data_bus[286]), .A2(n6217), .B1(
        i_data_bus[382]), .B2(n9877), .ZN(n9042) );
  ND2D1BWP30P140LVT U13194 ( .A1(n9043), .A2(n9042), .ZN(N10695) );
  AOI22D1BWP30P140LVT U13195 ( .A1(i_data_bus[273]), .A2(n6217), .B1(
        i_data_bus[305]), .B2(n9878), .ZN(n9045) );
  AOI22D1BWP30P140LVT U13196 ( .A1(i_data_bus[337]), .A2(n9879), .B1(
        i_data_bus[369]), .B2(n9877), .ZN(n9044) );
  ND2D1BWP30P140LVT U13197 ( .A1(n9045), .A2(n9044), .ZN(N10682) );
  AOI22D1BWP30P140LVT U13198 ( .A1(i_data_bus[303]), .A2(n9878), .B1(
        i_data_bus[335]), .B2(n9879), .ZN(n9047) );
  AOI22D1BWP30P140LVT U13199 ( .A1(i_data_bus[271]), .A2(n6217), .B1(
        i_data_bus[367]), .B2(n9877), .ZN(n9046) );
  ND2D1BWP30P140LVT U13200 ( .A1(n9047), .A2(n9046), .ZN(N10680) );
  AOI22D1BWP30P140LVT U13201 ( .A1(i_data_bus[295]), .A2(n9878), .B1(
        i_data_bus[327]), .B2(n9879), .ZN(n9049) );
  AOI22D1BWP30P140LVT U13202 ( .A1(i_data_bus[263]), .A2(n6217), .B1(
        i_data_bus[359]), .B2(n9877), .ZN(n9048) );
  ND2D1BWP30P140LVT U13203 ( .A1(n9049), .A2(n9048), .ZN(N10672) );
  AOI22D1BWP30P140LVT U13204 ( .A1(i_data_bus[317]), .A2(n9878), .B1(
        i_data_bus[285]), .B2(n6217), .ZN(n9051) );
  AOI22D1BWP30P140LVT U13205 ( .A1(i_data_bus[349]), .A2(n9879), .B1(
        i_data_bus[381]), .B2(n9877), .ZN(n9050) );
  ND2D1BWP30P140LVT U13206 ( .A1(n9051), .A2(n9050), .ZN(N10694) );
  AOI22D1BWP30P140LVT U13207 ( .A1(i_data_bus[315]), .A2(n9878), .B1(
        i_data_bus[347]), .B2(n9879), .ZN(n9053) );
  AOI22D1BWP30P140LVT U13208 ( .A1(i_data_bus[283]), .A2(n6217), .B1(
        i_data_bus[379]), .B2(n9877), .ZN(n9052) );
  ND2D1BWP30P140LVT U13209 ( .A1(n9053), .A2(n9052), .ZN(N10692) );
  AOI22D1BWP30P140LVT U13210 ( .A1(i_data_bus[316]), .A2(n9878), .B1(
        i_data_bus[348]), .B2(n9879), .ZN(n9055) );
  AOI22D1BWP30P140LVT U13211 ( .A1(i_data_bus[284]), .A2(n6217), .B1(
        i_data_bus[380]), .B2(n9877), .ZN(n9054) );
  ND2D1BWP30P140LVT U13212 ( .A1(n9055), .A2(n9054), .ZN(N10693) );
  AOI22D1BWP30P140LVT U13213 ( .A1(i_data_bus[212]), .A2(n10132), .B1(
        i_data_bus[180]), .B2(n10133), .ZN(n9057) );
  AOI22D1BWP30P140LVT U13214 ( .A1(i_data_bus[244]), .A2(n10131), .B1(
        i_data_bus[148]), .B2(n10134), .ZN(n9056) );
  ND2D1BWP30P140LVT U13215 ( .A1(n9057), .A2(n9056), .ZN(N7873) );
  AOI22D1BWP30P140LVT U13216 ( .A1(i_data_bus[197]), .A2(n10132), .B1(
        i_data_bus[165]), .B2(n10133), .ZN(n9059) );
  AOI22D1BWP30P140LVT U13217 ( .A1(i_data_bus[229]), .A2(n10131), .B1(
        i_data_bus[133]), .B2(n10134), .ZN(n9058) );
  ND2D1BWP30P140LVT U13218 ( .A1(n9059), .A2(n9058), .ZN(N7858) );
  AOI22D1BWP30P140LVT U13219 ( .A1(i_data_bus[216]), .A2(n10132), .B1(
        i_data_bus[184]), .B2(n10133), .ZN(n9061) );
  AOI22D1BWP30P140LVT U13220 ( .A1(i_data_bus[152]), .A2(n10134), .B1(
        i_data_bus[248]), .B2(n10131), .ZN(n9060) );
  ND2D1BWP30P140LVT U13221 ( .A1(n9061), .A2(n9060), .ZN(N7877) );
  AOI22D1BWP30P140LVT U13222 ( .A1(i_data_bus[151]), .A2(n10134), .B1(
        i_data_bus[183]), .B2(n10133), .ZN(n9063) );
  AOI22D1BWP30P140LVT U13223 ( .A1(i_data_bus[215]), .A2(n10132), .B1(
        i_data_bus[247]), .B2(n10131), .ZN(n9062) );
  ND2D1BWP30P140LVT U13224 ( .A1(n9063), .A2(n9062), .ZN(N7876) );
  AOI22D1BWP30P140LVT U13225 ( .A1(i_data_bus[146]), .A2(n10134), .B1(
        i_data_bus[178]), .B2(n10133), .ZN(n9065) );
  AOI22D1BWP30P140LVT U13226 ( .A1(i_data_bus[210]), .A2(n10132), .B1(
        i_data_bus[242]), .B2(n10131), .ZN(n9064) );
  ND2D1BWP30P140LVT U13227 ( .A1(n9065), .A2(n9064), .ZN(N7871) );
  AOI22D1BWP30P140LVT U13228 ( .A1(i_data_bus[350]), .A2(n9755), .B1(
        i_data_bus[382]), .B2(n9757), .ZN(n9067) );
  AOI22D1BWP30P140LVT U13229 ( .A1(i_data_bus[286]), .A2(n9756), .B1(
        i_data_bus[318]), .B2(n9758), .ZN(n9066) );
  ND2D1BWP30P140LVT U13230 ( .A1(n9067), .A2(n9066), .ZN(N5247) );
  AOI22D1BWP30P140LVT U13231 ( .A1(i_data_bus[259]), .A2(n9756), .B1(
        i_data_bus[323]), .B2(n9755), .ZN(n9069) );
  AOI22D1BWP30P140LVT U13232 ( .A1(i_data_bus[355]), .A2(n9757), .B1(
        i_data_bus[291]), .B2(n9758), .ZN(n9068) );
  ND2D1BWP30P140LVT U13233 ( .A1(n9069), .A2(n9068), .ZN(N5220) );
  AOI22D1BWP30P140LVT U13234 ( .A1(i_data_bus[380]), .A2(n9757), .B1(
        i_data_bus[348]), .B2(n9755), .ZN(n9071) );
  AOI22D1BWP30P140LVT U13235 ( .A1(i_data_bus[284]), .A2(n9756), .B1(
        i_data_bus[316]), .B2(n9758), .ZN(n9070) );
  ND2D1BWP30P140LVT U13236 ( .A1(n9071), .A2(n9070), .ZN(N5245) );
  AOI22D1BWP30P140LVT U13237 ( .A1(i_data_bus[280]), .A2(n9756), .B1(
        i_data_bus[344]), .B2(n9755), .ZN(n9073) );
  AOI22D1BWP30P140LVT U13238 ( .A1(i_data_bus[376]), .A2(n9757), .B1(
        i_data_bus[312]), .B2(n9758), .ZN(n9072) );
  ND2D1BWP30P140LVT U13239 ( .A1(n9073), .A2(n9072), .ZN(N5241) );
  AOI22D1BWP30P140LVT U13240 ( .A1(i_data_bus[371]), .A2(n9757), .B1(
        i_data_bus[339]), .B2(n9755), .ZN(n9075) );
  AOI22D1BWP30P140LVT U13241 ( .A1(i_data_bus[275]), .A2(n9756), .B1(
        i_data_bus[307]), .B2(n9758), .ZN(n9074) );
  ND2D1BWP30P140LVT U13242 ( .A1(n9075), .A2(n9074), .ZN(N5236) );
  AOI22D1BWP30P140LVT U13243 ( .A1(i_data_bus[364]), .A2(n9757), .B1(
        i_data_bus[332]), .B2(n9755), .ZN(n9077) );
  AOI22D1BWP30P140LVT U13244 ( .A1(i_data_bus[268]), .A2(n9756), .B1(
        i_data_bus[300]), .B2(n9758), .ZN(n9076) );
  ND2D1BWP30P140LVT U13245 ( .A1(n9077), .A2(n9076), .ZN(N5229) );
  AOI22D1BWP30P140LVT U13246 ( .A1(i_data_bus[262]), .A2(n9756), .B1(
        i_data_bus[326]), .B2(n9755), .ZN(n9079) );
  AOI22D1BWP30P140LVT U13247 ( .A1(i_data_bus[358]), .A2(n9757), .B1(
        i_data_bus[294]), .B2(n9758), .ZN(n9078) );
  ND2D1BWP30P140LVT U13248 ( .A1(n9079), .A2(n9078), .ZN(N5223) );
  AOI22D1BWP30P140LVT U13249 ( .A1(i_data_bus[256]), .A2(n9756), .B1(
        i_data_bus[352]), .B2(n9757), .ZN(n9081) );
  AOI22D1BWP30P140LVT U13250 ( .A1(i_data_bus[320]), .A2(n9755), .B1(
        i_data_bus[288]), .B2(n9758), .ZN(n9080) );
  ND2D1BWP30P140LVT U13251 ( .A1(n9081), .A2(n9080), .ZN(N5217) );
  AOI22D1BWP30P140LVT U13252 ( .A1(i_data_bus[95]), .A2(n10115), .B1(
        i_data_bus[31]), .B2(n10116), .ZN(n9083) );
  AOI22D1BWP30P140LVT U13253 ( .A1(i_data_bus[127]), .A2(n10117), .B1(
        i_data_bus[63]), .B2(n10118), .ZN(n9082) );
  ND2D1BWP30P140LVT U13254 ( .A1(n9083), .A2(n9082), .ZN(N7796) );
  AOI22D1BWP30P140LVT U13255 ( .A1(i_data_bus[27]), .A2(n10116), .B1(
        i_data_bus[123]), .B2(n10117), .ZN(n9085) );
  AOI22D1BWP30P140LVT U13256 ( .A1(i_data_bus[91]), .A2(n10115), .B1(
        i_data_bus[59]), .B2(n10118), .ZN(n9084) );
  ND2D1BWP30P140LVT U13257 ( .A1(n9085), .A2(n9084), .ZN(N7792) );
  AOI22D1BWP30P140LVT U13258 ( .A1(i_data_bus[121]), .A2(n10117), .B1(
        i_data_bus[89]), .B2(n10115), .ZN(n9087) );
  AOI22D1BWP30P140LVT U13259 ( .A1(i_data_bus[25]), .A2(n10116), .B1(
        i_data_bus[57]), .B2(n10118), .ZN(n9086) );
  ND2D1BWP30P140LVT U13260 ( .A1(n9087), .A2(n9086), .ZN(N7790) );
  AOI22D1BWP30P140LVT U13261 ( .A1(i_data_bus[15]), .A2(n10116), .B1(
        i_data_bus[111]), .B2(n10117), .ZN(n9089) );
  AOI22D1BWP30P140LVT U13262 ( .A1(i_data_bus[79]), .A2(n10115), .B1(
        i_data_bus[47]), .B2(n10118), .ZN(n9088) );
  ND2D1BWP30P140LVT U13263 ( .A1(n9089), .A2(n9088), .ZN(N7780) );
  AOI22D1BWP30P140LVT U13264 ( .A1(i_data_bus[77]), .A2(n10115), .B1(
        i_data_bus[109]), .B2(n10117), .ZN(n9091) );
  AOI22D1BWP30P140LVT U13265 ( .A1(i_data_bus[13]), .A2(n10116), .B1(
        i_data_bus[45]), .B2(n10118), .ZN(n9090) );
  ND2D1BWP30P140LVT U13266 ( .A1(n9091), .A2(n9090), .ZN(N7778) );
  AOI22D1BWP30P140LVT U13267 ( .A1(i_data_bus[74]), .A2(n10115), .B1(
        i_data_bus[10]), .B2(n10116), .ZN(n9093) );
  AOI22D1BWP30P140LVT U13268 ( .A1(i_data_bus[106]), .A2(n10117), .B1(
        i_data_bus[42]), .B2(n10118), .ZN(n9092) );
  ND2D1BWP30P140LVT U13269 ( .A1(n9093), .A2(n9092), .ZN(N7775) );
  AOI22D1BWP30P140LVT U13270 ( .A1(i_data_bus[102]), .A2(n10117), .B1(
        i_data_bus[70]), .B2(n10115), .ZN(n9095) );
  AOI22D1BWP30P140LVT U13271 ( .A1(i_data_bus[6]), .A2(n10116), .B1(
        i_data_bus[38]), .B2(n10118), .ZN(n9094) );
  ND2D1BWP30P140LVT U13272 ( .A1(n9095), .A2(n9094), .ZN(N7771) );
  AOI22D1BWP30P140LVT U13273 ( .A1(i_data_bus[5]), .A2(n10116), .B1(
        i_data_bus[101]), .B2(n10117), .ZN(n9097) );
  AOI22D1BWP30P140LVT U13274 ( .A1(i_data_bus[69]), .A2(n10115), .B1(
        i_data_bus[37]), .B2(n10118), .ZN(n9096) );
  ND2D1BWP30P140LVT U13275 ( .A1(n9097), .A2(n9096), .ZN(N7770) );
  AOI22D1BWP30P140LVT U13276 ( .A1(i_data_bus[3]), .A2(n10116), .B1(
        i_data_bus[67]), .B2(n10115), .ZN(n9099) );
  AOI22D1BWP30P140LVT U13277 ( .A1(i_data_bus[99]), .A2(n10117), .B1(
        i_data_bus[35]), .B2(n10118), .ZN(n9098) );
  ND2D1BWP30P140LVT U13278 ( .A1(n9099), .A2(n9098), .ZN(N7768) );
  AOI22D1BWP30P140LVT U13279 ( .A1(i_data_bus[95]), .A2(n9790), .B1(
        i_data_bus[31]), .B2(n6223), .ZN(n9101) );
  AOI22D1BWP30P140LVT U13280 ( .A1(i_data_bus[127]), .A2(n9792), .B1(
        i_data_bus[63]), .B2(n9791), .ZN(n9100) );
  ND2D1BWP30P140LVT U13281 ( .A1(n9101), .A2(n9100), .ZN(N8774) );
  AOI22D1BWP30P140LVT U13282 ( .A1(i_data_bus[84]), .A2(n9790), .B1(
        i_data_bus[116]), .B2(n9792), .ZN(n9103) );
  AOI22D1BWP30P140LVT U13283 ( .A1(i_data_bus[20]), .A2(n6223), .B1(
        i_data_bus[52]), .B2(n9791), .ZN(n9102) );
  ND2D1BWP30P140LVT U13284 ( .A1(n9103), .A2(n9102), .ZN(N8763) );
  AOI22D1BWP30P140LVT U13285 ( .A1(i_data_bus[15]), .A2(n6223), .B1(
        i_data_bus[79]), .B2(n9790), .ZN(n9105) );
  AOI22D1BWP30P140LVT U13286 ( .A1(i_data_bus[111]), .A2(n9792), .B1(
        i_data_bus[47]), .B2(n9791), .ZN(n9104) );
  ND2D1BWP30P140LVT U13287 ( .A1(n9105), .A2(n9104), .ZN(N8758) );
  AOI22D1BWP30P140LVT U13288 ( .A1(i_data_bus[9]), .A2(n6223), .B1(
        i_data_bus[105]), .B2(n9792), .ZN(n9107) );
  AOI22D1BWP30P140LVT U13289 ( .A1(i_data_bus[73]), .A2(n9790), .B1(
        i_data_bus[41]), .B2(n9791), .ZN(n9106) );
  ND2D1BWP30P140LVT U13290 ( .A1(n9107), .A2(n9106), .ZN(N8752) );
  AOI22D1BWP30P140LVT U13291 ( .A1(i_data_bus[101]), .A2(n9792), .B1(
        i_data_bus[69]), .B2(n9790), .ZN(n9109) );
  AOI22D1BWP30P140LVT U13292 ( .A1(i_data_bus[5]), .A2(n6223), .B1(
        i_data_bus[37]), .B2(n9791), .ZN(n9108) );
  ND2D1BWP30P140LVT U13293 ( .A1(n9109), .A2(n9108), .ZN(N8748) );
  AOI22D1BWP30P140LVT U13294 ( .A1(i_data_bus[78]), .A2(n9790), .B1(
        i_data_bus[110]), .B2(n9792), .ZN(n9111) );
  AOI22D1BWP30P140LVT U13295 ( .A1(i_data_bus[14]), .A2(n6223), .B1(
        i_data_bus[46]), .B2(n9791), .ZN(n9110) );
  ND2D1BWP30P140LVT U13296 ( .A1(n9111), .A2(n9110), .ZN(N8757) );
  AOI22D1BWP30P140LVT U13297 ( .A1(i_data_bus[24]), .A2(n6218), .B1(
        i_data_bus[88]), .B2(n9914), .ZN(n9113) );
  AOI22D1BWP30P140LVT U13298 ( .A1(i_data_bus[56]), .A2(n9916), .B1(
        i_data_bus[120]), .B2(n9915), .ZN(n9112) );
  ND2D1BWP30P140LVT U13299 ( .A1(n9113), .A2(n9112), .ZN(N3319) );
  AOI22D1BWP30P140LVT U13300 ( .A1(i_data_bus[50]), .A2(n9916), .B1(
        i_data_bus[82]), .B2(n9914), .ZN(n9115) );
  AOI22D1BWP30P140LVT U13301 ( .A1(i_data_bus[18]), .A2(n6218), .B1(
        i_data_bus[114]), .B2(n9915), .ZN(n9114) );
  ND2D1BWP30P140LVT U13302 ( .A1(n9115), .A2(n9114), .ZN(N3313) );
  AOI22D1BWP30P140LVT U13303 ( .A1(i_data_bus[16]), .A2(n6218), .B1(
        i_data_bus[80]), .B2(n9914), .ZN(n9117) );
  AOI22D1BWP30P140LVT U13304 ( .A1(i_data_bus[48]), .A2(n9916), .B1(
        i_data_bus[112]), .B2(n9915), .ZN(n9116) );
  ND2D1BWP30P140LVT U13305 ( .A1(n9117), .A2(n9116), .ZN(N3311) );
  AOI22D1BWP30P140LVT U13306 ( .A1(i_data_bus[43]), .A2(n9916), .B1(
        i_data_bus[75]), .B2(n9914), .ZN(n9119) );
  AOI22D1BWP30P140LVT U13307 ( .A1(i_data_bus[11]), .A2(n6218), .B1(
        i_data_bus[107]), .B2(n9915), .ZN(n9118) );
  ND2D1BWP30P140LVT U13308 ( .A1(n9119), .A2(n9118), .ZN(N3306) );
  AOI22D1BWP30P140LVT U13309 ( .A1(i_data_bus[73]), .A2(n9914), .B1(
        i_data_bus[41]), .B2(n9916), .ZN(n9121) );
  AOI22D1BWP30P140LVT U13310 ( .A1(i_data_bus[9]), .A2(n6218), .B1(
        i_data_bus[105]), .B2(n9915), .ZN(n9120) );
  ND2D1BWP30P140LVT U13311 ( .A1(n9121), .A2(n9120), .ZN(N3304) );
  AOI22D1BWP30P140LVT U13312 ( .A1(i_data_bus[4]), .A2(n6218), .B1(
        i_data_bus[68]), .B2(n9914), .ZN(n9123) );
  AOI22D1BWP30P140LVT U13313 ( .A1(i_data_bus[36]), .A2(n9916), .B1(
        i_data_bus[100]), .B2(n9915), .ZN(n9122) );
  ND2D1BWP30P140LVT U13314 ( .A1(n9123), .A2(n9122), .ZN(N3299) );
  AOI22D1BWP30P140LVT U13315 ( .A1(i_data_bus[32]), .A2(n9916), .B1(
        i_data_bus[64]), .B2(n9914), .ZN(n9125) );
  AOI22D1BWP30P140LVT U13316 ( .A1(i_data_bus[0]), .A2(n6218), .B1(
        i_data_bus[96]), .B2(n9915), .ZN(n9124) );
  ND2D1BWP30P140LVT U13317 ( .A1(n9125), .A2(n9124), .ZN(N3295) );
  AOI22D1BWP30P140LVT U13318 ( .A1(i_data_bus[606]), .A2(n10183), .B1(
        i_data_bus[574]), .B2(n10184), .ZN(n9127) );
  AOI22D1BWP30P140LVT U13319 ( .A1(i_data_bus[638]), .A2(n10185), .B1(
        i_data_bus[542]), .B2(n10182), .ZN(n9126) );
  ND2D1BWP30P140LVT U13320 ( .A1(n9127), .A2(n9126), .ZN(N6913) );
  AOI22D1BWP30P140LVT U13321 ( .A1(i_data_bus[587]), .A2(n10183), .B1(
        i_data_bus[555]), .B2(n10184), .ZN(n9129) );
  AOI22D1BWP30P140LVT U13322 ( .A1(i_data_bus[619]), .A2(n10185), .B1(
        i_data_bus[523]), .B2(n10182), .ZN(n9128) );
  ND2D1BWP30P140LVT U13323 ( .A1(n9129), .A2(n9128), .ZN(N6894) );
  AOI22D1BWP30P140LVT U13324 ( .A1(i_data_bus[380]), .A2(n9845), .B1(
        i_data_bus[348]), .B2(n9844), .ZN(n9131) );
  AOI22D1BWP30P140LVT U13325 ( .A1(i_data_bus[284]), .A2(n9846), .B1(
        i_data_bus[316]), .B2(n9843), .ZN(n9130) );
  ND2D1BWP30P140LVT U13326 ( .A1(n9131), .A2(n9130), .ZN(N7969) );
  AOI22D1BWP30P140LVT U13327 ( .A1(i_data_bus[346]), .A2(n9844), .B1(
        i_data_bus[378]), .B2(n9845), .ZN(n9133) );
  AOI22D1BWP30P140LVT U13328 ( .A1(i_data_bus[282]), .A2(n9846), .B1(
        i_data_bus[314]), .B2(n9843), .ZN(n9132) );
  ND2D1BWP30P140LVT U13329 ( .A1(n9133), .A2(n9132), .ZN(N7967) );
  AOI22D1BWP30P140LVT U13330 ( .A1(i_data_bus[340]), .A2(n9844), .B1(
        i_data_bus[372]), .B2(n9845), .ZN(n9135) );
  AOI22D1BWP30P140LVT U13331 ( .A1(i_data_bus[276]), .A2(n9846), .B1(
        i_data_bus[308]), .B2(n9843), .ZN(n9134) );
  ND2D1BWP30P140LVT U13332 ( .A1(n9135), .A2(n9134), .ZN(N7961) );
  AOI22D1BWP30P140LVT U13333 ( .A1(i_data_bus[368]), .A2(n9845), .B1(
        i_data_bus[336]), .B2(n9844), .ZN(n9137) );
  AOI22D1BWP30P140LVT U13334 ( .A1(i_data_bus[272]), .A2(n9846), .B1(
        i_data_bus[304]), .B2(n9843), .ZN(n9136) );
  ND2D1BWP30P140LVT U13335 ( .A1(n9137), .A2(n9136), .ZN(N7957) );
  AOI22D1BWP30P140LVT U13336 ( .A1(i_data_bus[331]), .A2(n9844), .B1(
        i_data_bus[267]), .B2(n9846), .ZN(n9139) );
  AOI22D1BWP30P140LVT U13337 ( .A1(i_data_bus[363]), .A2(n9845), .B1(
        i_data_bus[299]), .B2(n9843), .ZN(n9138) );
  ND2D1BWP30P140LVT U13338 ( .A1(n9139), .A2(n9138), .ZN(N7952) );
  AOI22D1BWP30P140LVT U13339 ( .A1(i_data_bus[356]), .A2(n9845), .B1(
        i_data_bus[324]), .B2(n9844), .ZN(n9141) );
  AOI22D1BWP30P140LVT U13340 ( .A1(i_data_bus[260]), .A2(n9846), .B1(
        i_data_bus[292]), .B2(n9843), .ZN(n9140) );
  ND2D1BWP30P140LVT U13341 ( .A1(n9141), .A2(n9140), .ZN(N7945) );
  AOI22D1BWP30P140LVT U13342 ( .A1(i_data_bus[355]), .A2(n9845), .B1(
        i_data_bus[323]), .B2(n9844), .ZN(n9143) );
  AOI22D1BWP30P140LVT U13343 ( .A1(i_data_bus[259]), .A2(n9846), .B1(
        i_data_bus[291]), .B2(n9843), .ZN(n9142) );
  ND2D1BWP30P140LVT U13344 ( .A1(n9143), .A2(n9142), .ZN(N7944) );
  AOI22D1BWP30P140LVT U13345 ( .A1(i_data_bus[27]), .A2(n9969), .B1(
        i_data_bus[123]), .B2(n9978), .ZN(n9145) );
  AOI22D1BWP30P140LVT U13346 ( .A1(i_data_bus[91]), .A2(n9976), .B1(
        i_data_bus[59]), .B2(n9977), .ZN(n9144) );
  ND2D1BWP30P140LVT U13347 ( .A1(n9145), .A2(n9144), .ZN(N2344) );
  AOI22D1BWP30P140LVT U13348 ( .A1(i_data_bus[81]), .A2(n9976), .B1(
        i_data_bus[113]), .B2(n9978), .ZN(n9147) );
  AOI22D1BWP30P140LVT U13349 ( .A1(i_data_bus[17]), .A2(n9969), .B1(
        i_data_bus[49]), .B2(n9977), .ZN(n9146) );
  ND2D1BWP30P140LVT U13350 ( .A1(n9147), .A2(n9146), .ZN(N2334) );
  AOI22D1BWP30P140LVT U13351 ( .A1(i_data_bus[111]), .A2(n9978), .B1(
        i_data_bus[79]), .B2(n9976), .ZN(n9149) );
  AOI22D1BWP30P140LVT U13352 ( .A1(i_data_bus[15]), .A2(n9969), .B1(
        i_data_bus[47]), .B2(n9977), .ZN(n9148) );
  ND2D1BWP30P140LVT U13353 ( .A1(n9149), .A2(n9148), .ZN(N2332) );
  AOI22D1BWP30P140LVT U13354 ( .A1(i_data_bus[76]), .A2(n9976), .B1(
        i_data_bus[108]), .B2(n9978), .ZN(n9151) );
  AOI22D1BWP30P140LVT U13355 ( .A1(i_data_bus[12]), .A2(n9969), .B1(
        i_data_bus[44]), .B2(n9977), .ZN(n9150) );
  ND2D1BWP30P140LVT U13356 ( .A1(n9151), .A2(n9150), .ZN(N2329) );
  AOI22D1BWP30P140LVT U13357 ( .A1(i_data_bus[74]), .A2(n9976), .B1(
        i_data_bus[10]), .B2(n9969), .ZN(n9153) );
  AOI22D1BWP30P140LVT U13358 ( .A1(i_data_bus[106]), .A2(n9978), .B1(
        i_data_bus[42]), .B2(n9977), .ZN(n9152) );
  ND2D1BWP30P140LVT U13359 ( .A1(n9153), .A2(n9152), .ZN(N2327) );
  AOI22D1BWP30P140LVT U13360 ( .A1(i_data_bus[64]), .A2(n9976), .B1(
        i_data_bus[96]), .B2(n9978), .ZN(n9155) );
  AOI22D1BWP30P140LVT U13361 ( .A1(i_data_bus[0]), .A2(n9969), .B1(
        i_data_bus[32]), .B2(n9977), .ZN(n9154) );
  ND2D1BWP30P140LVT U13362 ( .A1(n9155), .A2(n9154), .ZN(N2317) );
  AOI22D1BWP30P140LVT U13363 ( .A1(i_data_bus[112]), .A2(n9978), .B1(
        i_data_bus[80]), .B2(n9976), .ZN(n9157) );
  AOI22D1BWP30P140LVT U13364 ( .A1(i_data_bus[16]), .A2(n9969), .B1(
        i_data_bus[48]), .B2(n9977), .ZN(n9156) );
  ND2D1BWP30P140LVT U13365 ( .A1(n9157), .A2(n9156), .ZN(N2333) );
  AOI22D1BWP30P140LVT U13366 ( .A1(i_data_bus[95]), .A2(n9976), .B1(
        i_data_bus[31]), .B2(n9969), .ZN(n9159) );
  AOI22D1BWP30P140LVT U13367 ( .A1(i_data_bus[127]), .A2(n9978), .B1(
        i_data_bus[63]), .B2(n9977), .ZN(n9158) );
  ND2D1BWP30P140LVT U13368 ( .A1(n9159), .A2(n9158), .ZN(N2348) );
  AOI22D1BWP30P140LVT U13369 ( .A1(i_data_bus[26]), .A2(n9969), .B1(
        i_data_bus[122]), .B2(n9978), .ZN(n9161) );
  AOI22D1BWP30P140LVT U13370 ( .A1(i_data_bus[90]), .A2(n9976), .B1(
        i_data_bus[58]), .B2(n9977), .ZN(n9160) );
  ND2D1BWP30P140LVT U13371 ( .A1(n9161), .A2(n9160), .ZN(N2343) );
  AOI22D1BWP30P140LVT U13372 ( .A1(i_data_bus[143]), .A2(n10134), .B1(
        i_data_bus[175]), .B2(n10133), .ZN(n9163) );
  AOI22D1BWP30P140LVT U13373 ( .A1(i_data_bus[239]), .A2(n10131), .B1(
        i_data_bus[207]), .B2(n10132), .ZN(n9162) );
  ND2D1BWP30P140LVT U13374 ( .A1(n9163), .A2(n9162), .ZN(N7868) );
  AOI22D1BWP30P140LVT U13375 ( .A1(i_data_bus[188]), .A2(n10225), .B1(
        i_data_bus[156]), .B2(n10224), .ZN(n9165) );
  AOI22D1BWP30P140LVT U13376 ( .A1(i_data_bus[252]), .A2(n10226), .B1(
        i_data_bus[220]), .B2(n10223), .ZN(n9164) );
  ND2D1BWP30P140LVT U13377 ( .A1(n9165), .A2(n9164), .ZN(N6263) );
  AOI22D1BWP30P140LVT U13378 ( .A1(i_data_bus[179]), .A2(n10225), .B1(
        i_data_bus[147]), .B2(n10224), .ZN(n9167) );
  AOI22D1BWP30P140LVT U13379 ( .A1(i_data_bus[243]), .A2(n10226), .B1(
        i_data_bus[211]), .B2(n10223), .ZN(n9166) );
  ND2D1BWP30P140LVT U13380 ( .A1(n9167), .A2(n9166), .ZN(N6254) );
  AOI22D1BWP30P140LVT U13381 ( .A1(i_data_bus[176]), .A2(n10225), .B1(
        i_data_bus[240]), .B2(n10226), .ZN(n9169) );
  AOI22D1BWP30P140LVT U13382 ( .A1(i_data_bus[144]), .A2(n10224), .B1(
        i_data_bus[208]), .B2(n10223), .ZN(n9168) );
  ND2D1BWP30P140LVT U13383 ( .A1(n9169), .A2(n9168), .ZN(N6251) );
  AOI22D1BWP30P140LVT U13384 ( .A1(i_data_bus[143]), .A2(n10224), .B1(
        i_data_bus[239]), .B2(n10226), .ZN(n9171) );
  AOI22D1BWP30P140LVT U13385 ( .A1(i_data_bus[175]), .A2(n10225), .B1(
        i_data_bus[207]), .B2(n10223), .ZN(n9170) );
  ND2D1BWP30P140LVT U13386 ( .A1(n9171), .A2(n9170), .ZN(N6250) );
  AOI22D1BWP30P140LVT U13387 ( .A1(i_data_bus[161]), .A2(n10225), .B1(
        i_data_bus[129]), .B2(n10224), .ZN(n9173) );
  AOI22D1BWP30P140LVT U13388 ( .A1(i_data_bus[225]), .A2(n10226), .B1(
        i_data_bus[193]), .B2(n10223), .ZN(n9172) );
  ND2D1BWP30P140LVT U13389 ( .A1(n9173), .A2(n9172), .ZN(N6236) );
  AOI22D1BWP30P140LVT U13390 ( .A1(i_data_bus[179]), .A2(n10133), .B1(
        i_data_bus[147]), .B2(n10134), .ZN(n9175) );
  AOI22D1BWP30P140LVT U13391 ( .A1(i_data_bus[243]), .A2(n10131), .B1(
        i_data_bus[211]), .B2(n10132), .ZN(n9174) );
  ND2D1BWP30P140LVT U13392 ( .A1(n9175), .A2(n9174), .ZN(N7872) );
  AOI22D1BWP30P140LVT U13393 ( .A1(i_data_bus[172]), .A2(n10133), .B1(
        i_data_bus[236]), .B2(n10131), .ZN(n9177) );
  AOI22D1BWP30P140LVT U13394 ( .A1(i_data_bus[140]), .A2(n10134), .B1(
        i_data_bus[204]), .B2(n10132), .ZN(n9176) );
  ND2D1BWP30P140LVT U13395 ( .A1(n9177), .A2(n9176), .ZN(N7865) );
  AOI22D1BWP30P140LVT U13396 ( .A1(i_data_bus[160]), .A2(n10133), .B1(
        i_data_bus[128]), .B2(n10134), .ZN(n9179) );
  AOI22D1BWP30P140LVT U13397 ( .A1(i_data_bus[224]), .A2(n10131), .B1(
        i_data_bus[192]), .B2(n10132), .ZN(n9178) );
  ND2D1BWP30P140LVT U13398 ( .A1(n9179), .A2(n9178), .ZN(N7853) );
  AOI22D1BWP30P140LVT U13399 ( .A1(i_data_bus[153]), .A2(n10134), .B1(
        i_data_bus[185]), .B2(n10133), .ZN(n9181) );
  AOI22D1BWP30P140LVT U13400 ( .A1(i_data_bus[249]), .A2(n10131), .B1(
        i_data_bus[217]), .B2(n10132), .ZN(n9180) );
  ND2D1BWP30P140LVT U13401 ( .A1(n9181), .A2(n9180), .ZN(N7878) );
  AOI22D1BWP30P140LVT U13402 ( .A1(i_data_bus[131]), .A2(n10134), .B1(
        i_data_bus[163]), .B2(n10133), .ZN(n9183) );
  AOI22D1BWP30P140LVT U13403 ( .A1(i_data_bus[227]), .A2(n10131), .B1(
        i_data_bus[195]), .B2(n10132), .ZN(n9182) );
  ND2D1BWP30P140LVT U13404 ( .A1(n9183), .A2(n9182), .ZN(N7856) );
  AOI22D1BWP30P140LVT U13405 ( .A1(i_data_bus[253]), .A2(n10131), .B1(
        i_data_bus[189]), .B2(n10133), .ZN(n9185) );
  AOI22D1BWP30P140LVT U13406 ( .A1(i_data_bus[157]), .A2(n10134), .B1(
        i_data_bus[221]), .B2(n10132), .ZN(n9184) );
  ND2D1BWP30P140LVT U13407 ( .A1(n9185), .A2(n9184), .ZN(N7882) );
  AOI22D1BWP30P140LVT U13408 ( .A1(i_data_bus[155]), .A2(n10134), .B1(
        i_data_bus[187]), .B2(n10133), .ZN(n9187) );
  AOI22D1BWP30P140LVT U13409 ( .A1(i_data_bus[251]), .A2(n10131), .B1(
        i_data_bus[219]), .B2(n10132), .ZN(n9186) );
  ND2D1BWP30P140LVT U13410 ( .A1(n9187), .A2(n9186), .ZN(N7880) );
  AOI22D1BWP30P140LVT U13411 ( .A1(i_data_bus[154]), .A2(n9522), .B1(
        i_data_bus[250]), .B2(n9520), .ZN(n9189) );
  AOI22D1BWP30P140LVT U13412 ( .A1(i_data_bus[218]), .A2(n9521), .B1(
        i_data_bus[186]), .B2(n9519), .ZN(n9188) );
  ND2D1BWP30P140LVT U13413 ( .A1(n9189), .A2(n9188), .ZN(N5155) );
  AOI22D1BWP30P140LVT U13414 ( .A1(i_data_bus[152]), .A2(n9522), .B1(
        i_data_bus[248]), .B2(n9520), .ZN(n9191) );
  AOI22D1BWP30P140LVT U13415 ( .A1(i_data_bus[216]), .A2(n9521), .B1(
        i_data_bus[184]), .B2(n9519), .ZN(n9190) );
  ND2D1BWP30P140LVT U13416 ( .A1(n9191), .A2(n9190), .ZN(N5153) );
  AOI22D1BWP30P140LVT U13417 ( .A1(i_data_bus[151]), .A2(n9522), .B1(
        i_data_bus[215]), .B2(n9521), .ZN(n9193) );
  AOI22D1BWP30P140LVT U13418 ( .A1(i_data_bus[247]), .A2(n9520), .B1(
        i_data_bus[183]), .B2(n9519), .ZN(n9192) );
  ND2D1BWP30P140LVT U13419 ( .A1(n9193), .A2(n9192), .ZN(N5152) );
  AOI22D1BWP30P140LVT U13420 ( .A1(i_data_bus[213]), .A2(n9521), .B1(
        i_data_bus[245]), .B2(n9520), .ZN(n9195) );
  AOI22D1BWP30P140LVT U13421 ( .A1(i_data_bus[149]), .A2(n9522), .B1(
        i_data_bus[181]), .B2(n9519), .ZN(n9194) );
  ND2D1BWP30P140LVT U13422 ( .A1(n9195), .A2(n9194), .ZN(N5150) );
  AOI22D1BWP30P140LVT U13423 ( .A1(i_data_bus[210]), .A2(n9521), .B1(
        i_data_bus[242]), .B2(n9520), .ZN(n9197) );
  AOI22D1BWP30P140LVT U13424 ( .A1(i_data_bus[146]), .A2(n9522), .B1(
        i_data_bus[178]), .B2(n9519), .ZN(n9196) );
  ND2D1BWP30P140LVT U13425 ( .A1(n9197), .A2(n9196), .ZN(N5147) );
  AOI22D1BWP30P140LVT U13426 ( .A1(i_data_bus[71]), .A2(n10086), .B1(
        i_data_bus[39]), .B2(n10087), .ZN(n9199) );
  AOI22D1BWP30P140LVT U13427 ( .A1(i_data_bus[7]), .A2(n10088), .B1(
        i_data_bus[103]), .B2(n10085), .ZN(n9198) );
  ND2D1BWP30P140LVT U13428 ( .A1(n9199), .A2(n9198), .ZN(N5048) );
  AOI22D1BWP30P140LVT U13429 ( .A1(i_data_bus[70]), .A2(n10086), .B1(
        i_data_bus[38]), .B2(n10087), .ZN(n9201) );
  AOI22D1BWP30P140LVT U13430 ( .A1(i_data_bus[6]), .A2(n10088), .B1(
        i_data_bus[102]), .B2(n10085), .ZN(n9200) );
  ND2D1BWP30P140LVT U13431 ( .A1(n9201), .A2(n9200), .ZN(N5047) );
  AOI22D1BWP30P140LVT U13432 ( .A1(i_data_bus[82]), .A2(n10086), .B1(
        i_data_bus[18]), .B2(n10088), .ZN(n9203) );
  AOI22D1BWP30P140LVT U13433 ( .A1(i_data_bus[50]), .A2(n10087), .B1(
        i_data_bus[114]), .B2(n10085), .ZN(n9202) );
  ND2D1BWP30P140LVT U13434 ( .A1(n9203), .A2(n9202), .ZN(N5059) );
  AOI22D1BWP30P140LVT U13435 ( .A1(i_data_bus[20]), .A2(n10088), .B1(
        i_data_bus[84]), .B2(n10086), .ZN(n9205) );
  AOI22D1BWP30P140LVT U13436 ( .A1(i_data_bus[52]), .A2(n10087), .B1(
        i_data_bus[116]), .B2(n10085), .ZN(n9204) );
  ND2D1BWP30P140LVT U13437 ( .A1(n9205), .A2(n9204), .ZN(N5061) );
  AOI22D1BWP30P140LVT U13438 ( .A1(i_data_bus[10]), .A2(n10088), .B1(
        i_data_bus[42]), .B2(n10087), .ZN(n9207) );
  AOI22D1BWP30P140LVT U13439 ( .A1(i_data_bus[74]), .A2(n10086), .B1(
        i_data_bus[106]), .B2(n10085), .ZN(n9206) );
  ND2D1BWP30P140LVT U13440 ( .A1(n9207), .A2(n9206), .ZN(N5051) );
  AOI22D1BWP30P140LVT U13441 ( .A1(i_data_bus[92]), .A2(n10086), .B1(
        i_data_bus[28]), .B2(n10088), .ZN(n9209) );
  AOI22D1BWP30P140LVT U13442 ( .A1(i_data_bus[60]), .A2(n10087), .B1(
        i_data_bus[124]), .B2(n10085), .ZN(n9208) );
  ND2D1BWP30P140LVT U13443 ( .A1(n9209), .A2(n9208), .ZN(N5069) );
  AOI22D1BWP30P140LVT U13444 ( .A1(i_data_bus[11]), .A2(n10088), .B1(
        i_data_bus[75]), .B2(n10086), .ZN(n9211) );
  AOI22D1BWP30P140LVT U13445 ( .A1(i_data_bus[43]), .A2(n10087), .B1(
        i_data_bus[107]), .B2(n10085), .ZN(n9210) );
  ND2D1BWP30P140LVT U13446 ( .A1(n9211), .A2(n9210), .ZN(N5052) );
  AOI22D1BWP30P140LVT U13447 ( .A1(i_data_bus[282]), .A2(n6216), .B1(
        i_data_bus[314]), .B2(n9775), .ZN(n9213) );
  AOI22D1BWP30P140LVT U13448 ( .A1(i_data_bus[346]), .A2(n9774), .B1(
        i_data_bus[378]), .B2(n9773), .ZN(n9212) );
  ND2D1BWP30P140LVT U13449 ( .A1(n9213), .A2(n9212), .ZN(N2519) );
  AOI22D1BWP30P140LVT U13450 ( .A1(i_data_bus[350]), .A2(n9774), .B1(
        i_data_bus[318]), .B2(n9775), .ZN(n9215) );
  AOI22D1BWP30P140LVT U13451 ( .A1(i_data_bus[286]), .A2(n6216), .B1(
        i_data_bus[382]), .B2(n9773), .ZN(n9214) );
  ND2D1BWP30P140LVT U13452 ( .A1(n9215), .A2(n9214), .ZN(N2523) );
  AOI22D1BWP30P140LVT U13453 ( .A1(i_data_bus[278]), .A2(n6216), .B1(
        i_data_bus[310]), .B2(n9775), .ZN(n9217) );
  AOI22D1BWP30P140LVT U13454 ( .A1(i_data_bus[342]), .A2(n9774), .B1(
        i_data_bus[374]), .B2(n9773), .ZN(n9216) );
  ND2D1BWP30P140LVT U13455 ( .A1(n9217), .A2(n9216), .ZN(N2515) );
  AOI22D1BWP30P140LVT U13456 ( .A1(i_data_bus[303]), .A2(n9775), .B1(
        i_data_bus[271]), .B2(n6216), .ZN(n9219) );
  AOI22D1BWP30P140LVT U13457 ( .A1(i_data_bus[335]), .A2(n9774), .B1(
        i_data_bus[367]), .B2(n9773), .ZN(n9218) );
  ND2D1BWP30P140LVT U13458 ( .A1(n9219), .A2(n9218), .ZN(N2508) );
  AOI22D1BWP30P140LVT U13459 ( .A1(i_data_bus[332]), .A2(n9774), .B1(
        i_data_bus[300]), .B2(n9775), .ZN(n9221) );
  AOI22D1BWP30P140LVT U13460 ( .A1(i_data_bus[268]), .A2(n6216), .B1(
        i_data_bus[364]), .B2(n9773), .ZN(n9220) );
  ND2D1BWP30P140LVT U13461 ( .A1(n9221), .A2(n9220), .ZN(N2505) );
  AOI22D1BWP30P140LVT U13462 ( .A1(i_data_bus[293]), .A2(n9775), .B1(
        i_data_bus[325]), .B2(n9774), .ZN(n9223) );
  AOI22D1BWP30P140LVT U13463 ( .A1(i_data_bus[261]), .A2(n6216), .B1(
        i_data_bus[357]), .B2(n9773), .ZN(n9222) );
  ND2D1BWP30P140LVT U13464 ( .A1(n9223), .A2(n9222), .ZN(N2498) );
  AOI22D1BWP30P140LVT U13465 ( .A1(i_data_bus[322]), .A2(n9774), .B1(
        i_data_bus[290]), .B2(n9775), .ZN(n9225) );
  AOI22D1BWP30P140LVT U13466 ( .A1(i_data_bus[258]), .A2(n6216), .B1(
        i_data_bus[354]), .B2(n9773), .ZN(n9224) );
  ND2D1BWP30P140LVT U13467 ( .A1(n9225), .A2(n9224), .ZN(N2495) );
  AOI22D1BWP30P140LVT U13468 ( .A1(i_data_bus[289]), .A2(n9775), .B1(
        i_data_bus[257]), .B2(n6216), .ZN(n9227) );
  AOI22D1BWP30P140LVT U13469 ( .A1(i_data_bus[321]), .A2(n9774), .B1(
        i_data_bus[353]), .B2(n9773), .ZN(n9226) );
  ND2D1BWP30P140LVT U13470 ( .A1(n9227), .A2(n9226), .ZN(N2494) );
  AOI22D1BWP30P140LVT U13471 ( .A1(i_data_bus[209]), .A2(n9521), .B1(
        i_data_bus[145]), .B2(n9522), .ZN(n9229) );
  AOI22D1BWP30P140LVT U13472 ( .A1(i_data_bus[177]), .A2(n9519), .B1(
        i_data_bus[241]), .B2(n9520), .ZN(n9228) );
  ND2D1BWP30P140LVT U13473 ( .A1(n9229), .A2(n9228), .ZN(N5146) );
  AOI22D1BWP30P140LVT U13474 ( .A1(i_data_bus[173]), .A2(n9519), .B1(
        i_data_bus[141]), .B2(n9522), .ZN(n9231) );
  AOI22D1BWP30P140LVT U13475 ( .A1(i_data_bus[205]), .A2(n9521), .B1(
        i_data_bus[237]), .B2(n9520), .ZN(n9230) );
  ND2D1BWP30P140LVT U13476 ( .A1(n9231), .A2(n9230), .ZN(N5142) );
  AOI22D1BWP30P140LVT U13477 ( .A1(i_data_bus[143]), .A2(n9522), .B1(
        i_data_bus[207]), .B2(n9521), .ZN(n9233) );
  AOI22D1BWP30P140LVT U13478 ( .A1(i_data_bus[175]), .A2(n9519), .B1(
        i_data_bus[239]), .B2(n9520), .ZN(n9232) );
  ND2D1BWP30P140LVT U13479 ( .A1(n9233), .A2(n9232), .ZN(N5144) );
  AOI22D1BWP30P140LVT U13480 ( .A1(i_data_bus[191]), .A2(n9519), .B1(
        i_data_bus[159]), .B2(n9522), .ZN(n9235) );
  AOI22D1BWP30P140LVT U13481 ( .A1(i_data_bus[223]), .A2(n9521), .B1(
        i_data_bus[255]), .B2(n9520), .ZN(n9234) );
  ND2D1BWP30P140LVT U13482 ( .A1(n9235), .A2(n9234), .ZN(N5160) );
  AOI22D1BWP30P140LVT U13483 ( .A1(i_data_bus[214]), .A2(n9521), .B1(
        i_data_bus[182]), .B2(n9519), .ZN(n9237) );
  AOI22D1BWP30P140LVT U13484 ( .A1(i_data_bus[150]), .A2(n9522), .B1(
        i_data_bus[246]), .B2(n9520), .ZN(n9236) );
  ND2D1BWP30P140LVT U13485 ( .A1(n9237), .A2(n9236), .ZN(N5151) );
  AOI22D1BWP30P140LVT U13486 ( .A1(i_data_bus[147]), .A2(n9522), .B1(
        i_data_bus[211]), .B2(n9521), .ZN(n9239) );
  AOI22D1BWP30P140LVT U13487 ( .A1(i_data_bus[179]), .A2(n9519), .B1(
        i_data_bus[243]), .B2(n9520), .ZN(n9238) );
  ND2D1BWP30P140LVT U13488 ( .A1(n9239), .A2(n9238), .ZN(N5148) );
  AOI22D1BWP30P140LVT U13489 ( .A1(i_data_bus[194]), .A2(n9521), .B1(
        i_data_bus[130]), .B2(n9522), .ZN(n9241) );
  AOI22D1BWP30P140LVT U13490 ( .A1(i_data_bus[162]), .A2(n9519), .B1(
        i_data_bus[226]), .B2(n9520), .ZN(n9240) );
  ND2D1BWP30P140LVT U13491 ( .A1(n9241), .A2(n9240), .ZN(N5131) );
  AOI22D1BWP30P140LVT U13492 ( .A1(i_data_bus[137]), .A2(n9522), .B1(
        i_data_bus[201]), .B2(n9521), .ZN(n9243) );
  AOI22D1BWP30P140LVT U13493 ( .A1(i_data_bus[169]), .A2(n9519), .B1(
        i_data_bus[233]), .B2(n9520), .ZN(n9242) );
  ND2D1BWP30P140LVT U13494 ( .A1(n9243), .A2(n9242), .ZN(N5138) );
  AOI22D1BWP30P140LVT U13495 ( .A1(i_data_bus[213]), .A2(n10218), .B1(
        i_data_bus[181]), .B2(n10219), .ZN(n9245) );
  AOI22D1BWP30P140LVT U13496 ( .A1(i_data_bus[245]), .A2(n10220), .B1(
        i_data_bus[149]), .B2(n6213), .ZN(n9244) );
  ND2D1BWP30P140LVT U13497 ( .A1(n9245), .A2(n9244), .ZN(N2426) );
  AOI22D1BWP30P140LVT U13498 ( .A1(i_data_bus[197]), .A2(n10218), .B1(
        i_data_bus[165]), .B2(n10219), .ZN(n9247) );
  AOI22D1BWP30P140LVT U13499 ( .A1(i_data_bus[229]), .A2(n10220), .B1(
        i_data_bus[133]), .B2(n6213), .ZN(n9246) );
  ND2D1BWP30P140LVT U13500 ( .A1(n9247), .A2(n9246), .ZN(N2410) );
  AOI22D1BWP30P140LVT U13501 ( .A1(i_data_bus[213]), .A2(n10223), .B1(
        i_data_bus[181]), .B2(n10225), .ZN(n9249) );
  AOI22D1BWP30P140LVT U13502 ( .A1(i_data_bus[245]), .A2(n10226), .B1(
        i_data_bus[149]), .B2(n10224), .ZN(n9248) );
  ND2D1BWP30P140LVT U13503 ( .A1(n9249), .A2(n9248), .ZN(N6256) );
  AOI22D1BWP30P140LVT U13504 ( .A1(i_data_bus[229]), .A2(n10226), .B1(
        i_data_bus[165]), .B2(n10225), .ZN(n9251) );
  AOI22D1BWP30P140LVT U13505 ( .A1(i_data_bus[197]), .A2(n10223), .B1(
        i_data_bus[133]), .B2(n10224), .ZN(n9250) );
  ND2D1BWP30P140LVT U13506 ( .A1(n9251), .A2(n9250), .ZN(N6240) );
  AOI22D1BWP30P140LVT U13507 ( .A1(i_data_bus[254]), .A2(n10220), .B1(
        i_data_bus[190]), .B2(n10219), .ZN(n9253) );
  AOI22D1BWP30P140LVT U13508 ( .A1(i_data_bus[222]), .A2(n10218), .B1(
        i_data_bus[158]), .B2(n6213), .ZN(n9252) );
  ND2D1BWP30P140LVT U13509 ( .A1(n9253), .A2(n9252), .ZN(N2435) );
  AOI22D1BWP30P140LVT U13510 ( .A1(i_data_bus[154]), .A2(n6213), .B1(
        i_data_bus[186]), .B2(n10219), .ZN(n9255) );
  AOI22D1BWP30P140LVT U13511 ( .A1(i_data_bus[218]), .A2(n10218), .B1(
        i_data_bus[250]), .B2(n10220), .ZN(n9254) );
  ND2D1BWP30P140LVT U13512 ( .A1(n9255), .A2(n9254), .ZN(N2431) );
  AOI22D1BWP30P140LVT U13513 ( .A1(i_data_bus[152]), .A2(n6213), .B1(
        i_data_bus[184]), .B2(n10219), .ZN(n9257) );
  AOI22D1BWP30P140LVT U13514 ( .A1(i_data_bus[216]), .A2(n10218), .B1(
        i_data_bus[248]), .B2(n10220), .ZN(n9256) );
  ND2D1BWP30P140LVT U13515 ( .A1(n9257), .A2(n9256), .ZN(N2429) );
  AOI22D1BWP30P140LVT U13516 ( .A1(i_data_bus[214]), .A2(n10218), .B1(
        i_data_bus[182]), .B2(n10219), .ZN(n9259) );
  AOI22D1BWP30P140LVT U13517 ( .A1(i_data_bus[150]), .A2(n6213), .B1(
        i_data_bus[246]), .B2(n10220), .ZN(n9258) );
  ND2D1BWP30P140LVT U13518 ( .A1(n9259), .A2(n9258), .ZN(N2427) );
  AOI22D1BWP30P140LVT U13519 ( .A1(i_data_bus[195]), .A2(n10218), .B1(
        i_data_bus[163]), .B2(n10219), .ZN(n9261) );
  AOI22D1BWP30P140LVT U13520 ( .A1(i_data_bus[131]), .A2(n6213), .B1(
        i_data_bus[227]), .B2(n10220), .ZN(n9260) );
  ND2D1BWP30P140LVT U13521 ( .A1(n9261), .A2(n9260), .ZN(N2408) );
  AOI22D1BWP30P140LVT U13522 ( .A1(i_data_bus[154]), .A2(n10224), .B1(
        i_data_bus[186]), .B2(n10225), .ZN(n9263) );
  AOI22D1BWP30P140LVT U13523 ( .A1(i_data_bus[218]), .A2(n10223), .B1(
        i_data_bus[250]), .B2(n10226), .ZN(n9262) );
  ND2D1BWP30P140LVT U13524 ( .A1(n9263), .A2(n9262), .ZN(N6261) );
  AOI22D1BWP30P140LVT U13525 ( .A1(i_data_bus[216]), .A2(n10223), .B1(
        i_data_bus[184]), .B2(n10225), .ZN(n9265) );
  AOI22D1BWP30P140LVT U13526 ( .A1(i_data_bus[152]), .A2(n10224), .B1(
        i_data_bus[248]), .B2(n10226), .ZN(n9264) );
  ND2D1BWP30P140LVT U13527 ( .A1(n9265), .A2(n9264), .ZN(N6259) );
  AOI22D1BWP30P140LVT U13528 ( .A1(i_data_bus[210]), .A2(n10223), .B1(
        i_data_bus[178]), .B2(n10225), .ZN(n9267) );
  AOI22D1BWP30P140LVT U13529 ( .A1(i_data_bus[146]), .A2(n10224), .B1(
        i_data_bus[242]), .B2(n10226), .ZN(n9266) );
  ND2D1BWP30P140LVT U13530 ( .A1(n9267), .A2(n9266), .ZN(N6253) );
  AOI22D1BWP30P140LVT U13531 ( .A1(i_data_bus[151]), .A2(n10224), .B1(
        i_data_bus[183]), .B2(n10225), .ZN(n9269) );
  AOI22D1BWP30P140LVT U13532 ( .A1(i_data_bus[215]), .A2(n10223), .B1(
        i_data_bus[247]), .B2(n10226), .ZN(n9268) );
  ND2D1BWP30P140LVT U13533 ( .A1(n9269), .A2(n9268), .ZN(N6258) );
  AOI22D1BWP30P140LVT U13534 ( .A1(i_data_bus[135]), .A2(n10224), .B1(
        i_data_bus[167]), .B2(n10225), .ZN(n9271) );
  AOI22D1BWP30P140LVT U13535 ( .A1(i_data_bus[231]), .A2(n10226), .B1(
        i_data_bus[199]), .B2(n10223), .ZN(n9270) );
  ND2D1BWP30P140LVT U13536 ( .A1(n9271), .A2(n9270), .ZN(N6242) );
  AOI22D1BWP30P140LVT U13537 ( .A1(i_data_bus[234]), .A2(n10226), .B1(
        i_data_bus[170]), .B2(n10225), .ZN(n9273) );
  AOI22D1BWP30P140LVT U13538 ( .A1(i_data_bus[138]), .A2(n10224), .B1(
        i_data_bus[202]), .B2(n10223), .ZN(n9272) );
  ND2D1BWP30P140LVT U13539 ( .A1(n9273), .A2(n9272), .ZN(N6245) );
  AOI22D1BWP30P140LVT U13540 ( .A1(i_data_bus[232]), .A2(n10226), .B1(
        i_data_bus[168]), .B2(n10225), .ZN(n9275) );
  AOI22D1BWP30P140LVT U13541 ( .A1(i_data_bus[136]), .A2(n10224), .B1(
        i_data_bus[200]), .B2(n10223), .ZN(n9274) );
  ND2D1BWP30P140LVT U13542 ( .A1(n9275), .A2(n9274), .ZN(N6243) );
  AOI22D1BWP30P140LVT U13543 ( .A1(i_data_bus[174]), .A2(n10040), .B1(
        i_data_bus[238]), .B2(n10038), .ZN(n9277) );
  AOI22D1BWP30P140LVT U13544 ( .A1(i_data_bus[142]), .A2(n9318), .B1(
        i_data_bus[206]), .B2(n10039), .ZN(n9276) );
  ND2D1BWP30P140LVT U13545 ( .A1(n9277), .A2(n9276), .ZN(N8973) );
  AOI22D1BWP30P140LVT U13546 ( .A1(i_data_bus[30]), .A2(n10096), .B1(
        i_data_bus[62]), .B2(n10097), .ZN(n9279) );
  AOI22D1BWP30P140LVT U13547 ( .A1(i_data_bus[126]), .A2(n10098), .B1(
        i_data_bus[94]), .B2(n10095), .ZN(n9278) );
  ND2D1BWP30P140LVT U13548 ( .A1(n9279), .A2(n9278), .ZN(N6049) );
  AOI22D1BWP30P140LVT U13549 ( .A1(i_data_bus[21]), .A2(n10096), .B1(
        i_data_bus[53]), .B2(n10097), .ZN(n9281) );
  AOI22D1BWP30P140LVT U13550 ( .A1(i_data_bus[117]), .A2(n10098), .B1(
        i_data_bus[85]), .B2(n10095), .ZN(n9280) );
  ND2D1BWP30P140LVT U13551 ( .A1(n9281), .A2(n9280), .ZN(N6040) );
  AOI22D1BWP30P140LVT U13552 ( .A1(i_data_bus[51]), .A2(n10097), .B1(
        i_data_bus[115]), .B2(n10098), .ZN(n9283) );
  AOI22D1BWP30P140LVT U13553 ( .A1(i_data_bus[19]), .A2(n10096), .B1(
        i_data_bus[83]), .B2(n10095), .ZN(n9282) );
  ND2D1BWP30P140LVT U13554 ( .A1(n9283), .A2(n9282), .ZN(N6038) );
  AOI22D1BWP30P140LVT U13555 ( .A1(i_data_bus[1]), .A2(n10096), .B1(
        i_data_bus[33]), .B2(n10097), .ZN(n9285) );
  AOI22D1BWP30P140LVT U13556 ( .A1(i_data_bus[97]), .A2(n10098), .B1(
        i_data_bus[65]), .B2(n10095), .ZN(n9284) );
  ND2D1BWP30P140LVT U13557 ( .A1(n9285), .A2(n9284), .ZN(N6020) );
  AOI22D1BWP30P140LVT U13558 ( .A1(i_data_bus[0]), .A2(n10096), .B1(
        i_data_bus[96]), .B2(n10098), .ZN(n9287) );
  AOI22D1BWP30P140LVT U13559 ( .A1(i_data_bus[32]), .A2(n10097), .B1(
        i_data_bus[64]), .B2(n10095), .ZN(n9286) );
  ND2D1BWP30P140LVT U13560 ( .A1(n9287), .A2(n9286), .ZN(N6019) );
  AOI22D1BWP30P140LVT U13561 ( .A1(i_data_bus[136]), .A2(n9318), .B1(
        i_data_bus[232]), .B2(n10038), .ZN(n9289) );
  AOI22D1BWP30P140LVT U13562 ( .A1(i_data_bus[168]), .A2(n10040), .B1(
        i_data_bus[200]), .B2(n10039), .ZN(n9288) );
  ND2D1BWP30P140LVT U13563 ( .A1(n9289), .A2(n9288), .ZN(N8967) );
  AOI22D1BWP30P140LVT U13564 ( .A1(i_data_bus[35]), .A2(n10097), .B1(
        i_data_bus[3]), .B2(n10096), .ZN(n9291) );
  AOI22D1BWP30P140LVT U13565 ( .A1(i_data_bus[99]), .A2(n10098), .B1(
        i_data_bus[67]), .B2(n10095), .ZN(n9290) );
  ND2D1BWP30P140LVT U13566 ( .A1(n9291), .A2(n9290), .ZN(N6022) );
  AOI22D1BWP30P140LVT U13567 ( .A1(i_data_bus[230]), .A2(n10038), .B1(
        i_data_bus[134]), .B2(n9318), .ZN(n9293) );
  AOI22D1BWP30P140LVT U13568 ( .A1(i_data_bus[166]), .A2(n10040), .B1(
        i_data_bus[198]), .B2(n10039), .ZN(n9292) );
  ND2D1BWP30P140LVT U13569 ( .A1(n9293), .A2(n9292), .ZN(N8965) );
  AOI22D1BWP30P140LVT U13570 ( .A1(i_data_bus[316]), .A2(n9775), .B1(
        i_data_bus[380]), .B2(n9773), .ZN(n9295) );
  AOI22D1BWP30P140LVT U13571 ( .A1(i_data_bus[284]), .A2(n6216), .B1(
        i_data_bus[348]), .B2(n9774), .ZN(n9294) );
  ND2D1BWP30P140LVT U13572 ( .A1(n9295), .A2(n9294), .ZN(N2521) );
  AOI22D1BWP30P140LVT U13573 ( .A1(i_data_bus[283]), .A2(n6216), .B1(
        i_data_bus[379]), .B2(n9773), .ZN(n9297) );
  AOI22D1BWP30P140LVT U13574 ( .A1(i_data_bus[315]), .A2(n9775), .B1(
        i_data_bus[347]), .B2(n9774), .ZN(n9296) );
  ND2D1BWP30P140LVT U13575 ( .A1(n9297), .A2(n9296), .ZN(N2520) );
  AOI22D1BWP30P140LVT U13576 ( .A1(i_data_bus[377]), .A2(n9773), .B1(
        i_data_bus[281]), .B2(n6216), .ZN(n9299) );
  AOI22D1BWP30P140LVT U13577 ( .A1(i_data_bus[313]), .A2(n9775), .B1(
        i_data_bus[345]), .B2(n9774), .ZN(n9298) );
  ND2D1BWP30P140LVT U13578 ( .A1(n9299), .A2(n9298), .ZN(N2518) );
  AOI22D1BWP30P140LVT U13579 ( .A1(i_data_bus[272]), .A2(n6216), .B1(
        i_data_bus[368]), .B2(n9773), .ZN(n9301) );
  AOI22D1BWP30P140LVT U13580 ( .A1(i_data_bus[304]), .A2(n9775), .B1(
        i_data_bus[336]), .B2(n9774), .ZN(n9300) );
  ND2D1BWP30P140LVT U13581 ( .A1(n9301), .A2(n9300), .ZN(N2509) );
  AOI22D1BWP30P140LVT U13582 ( .A1(i_data_bus[363]), .A2(n9773), .B1(
        i_data_bus[267]), .B2(n6216), .ZN(n9303) );
  AOI22D1BWP30P140LVT U13583 ( .A1(i_data_bus[299]), .A2(n9775), .B1(
        i_data_bus[331]), .B2(n9774), .ZN(n9302) );
  ND2D1BWP30P140LVT U13584 ( .A1(n9303), .A2(n9302), .ZN(N2504) );
  AOI22D1BWP30P140LVT U13585 ( .A1(i_data_bus[266]), .A2(n6216), .B1(
        i_data_bus[362]), .B2(n9773), .ZN(n9305) );
  AOI22D1BWP30P140LVT U13586 ( .A1(i_data_bus[298]), .A2(n9775), .B1(
        i_data_bus[330]), .B2(n9774), .ZN(n9304) );
  ND2D1BWP30P140LVT U13587 ( .A1(n9305), .A2(n9304), .ZN(N2503) );
  AOI22D1BWP30P140LVT U13588 ( .A1(i_data_bus[295]), .A2(n9775), .B1(
        i_data_bus[359]), .B2(n9773), .ZN(n9307) );
  AOI22D1BWP30P140LVT U13589 ( .A1(i_data_bus[263]), .A2(n6216), .B1(
        i_data_bus[327]), .B2(n9774), .ZN(n9306) );
  ND2D1BWP30P140LVT U13590 ( .A1(n9307), .A2(n9306), .ZN(N2500) );
  AOI22D1BWP30P140LVT U13591 ( .A1(i_data_bus[131]), .A2(n9318), .B1(
        i_data_bus[163]), .B2(n10040), .ZN(n9309) );
  AOI22D1BWP30P140LVT U13592 ( .A1(i_data_bus[227]), .A2(n10038), .B1(
        i_data_bus[195]), .B2(n10039), .ZN(n9308) );
  ND2D1BWP30P140LVT U13593 ( .A1(n9309), .A2(n9308), .ZN(N8962) );
  AOI22D1BWP30P140LVT U13594 ( .A1(i_data_bus[260]), .A2(n6216), .B1(
        i_data_bus[356]), .B2(n9773), .ZN(n9311) );
  AOI22D1BWP30P140LVT U13595 ( .A1(i_data_bus[292]), .A2(n9775), .B1(
        i_data_bus[324]), .B2(n9774), .ZN(n9310) );
  ND2D1BWP30P140LVT U13596 ( .A1(n9311), .A2(n9310), .ZN(N2497) );
  AOI22D1BWP30P140LVT U13597 ( .A1(i_data_bus[355]), .A2(n9773), .B1(
        i_data_bus[291]), .B2(n9775), .ZN(n9313) );
  AOI22D1BWP30P140LVT U13598 ( .A1(i_data_bus[259]), .A2(n6216), .B1(
        i_data_bus[323]), .B2(n9774), .ZN(n9312) );
  ND2D1BWP30P140LVT U13599 ( .A1(n9313), .A2(n9312), .ZN(N2496) );
  AOI22D1BWP30P140LVT U13600 ( .A1(i_data_bus[8]), .A2(n10096), .B1(
        i_data_bus[40]), .B2(n10097), .ZN(n9315) );
  AOI22D1BWP30P140LVT U13601 ( .A1(i_data_bus[104]), .A2(n10098), .B1(
        i_data_bus[72]), .B2(n10095), .ZN(n9314) );
  ND2D1BWP30P140LVT U13602 ( .A1(n9315), .A2(n9314), .ZN(N6027) );
  AOI22D1BWP30P140LVT U13603 ( .A1(i_data_bus[279]), .A2(n6216), .B1(
        i_data_bus[311]), .B2(n9775), .ZN(n9317) );
  AOI22D1BWP30P140LVT U13604 ( .A1(i_data_bus[375]), .A2(n9773), .B1(
        i_data_bus[343]), .B2(n9774), .ZN(n9316) );
  ND2D1BWP30P140LVT U13605 ( .A1(n9317), .A2(n9316), .ZN(N2516) );
  AOI22D1BWP30P140LVT U13606 ( .A1(i_data_bus[252]), .A2(n10038), .B1(
        i_data_bus[156]), .B2(n9318), .ZN(n9320) );
  AOI22D1BWP30P140LVT U13607 ( .A1(i_data_bus[188]), .A2(n10040), .B1(
        i_data_bus[220]), .B2(n10039), .ZN(n9319) );
  ND2D1BWP30P140LVT U13608 ( .A1(n9320), .A2(n9319), .ZN(N8987) );
  AOI22D1BWP30P140LVT U13609 ( .A1(i_data_bus[169]), .A2(n10040), .B1(
        i_data_bus[233]), .B2(n10038), .ZN(n9322) );
  AOI22D1BWP30P140LVT U13610 ( .A1(i_data_bus[137]), .A2(n9318), .B1(
        i_data_bus[201]), .B2(n10039), .ZN(n9321) );
  ND2D1BWP30P140LVT U13611 ( .A1(n9322), .A2(n9321), .ZN(N8968) );
  AOI22D1BWP30P140LVT U13612 ( .A1(i_data_bus[34]), .A2(n10097), .B1(
        i_data_bus[98]), .B2(n10098), .ZN(n9324) );
  AOI22D1BWP30P140LVT U13613 ( .A1(i_data_bus[2]), .A2(n10096), .B1(
        i_data_bus[66]), .B2(n10095), .ZN(n9323) );
  ND2D1BWP30P140LVT U13614 ( .A1(n9324), .A2(n9323), .ZN(N6021) );
  AOI22D1BWP30P140LVT U13615 ( .A1(i_data_bus[155]), .A2(n9318), .B1(
        i_data_bus[251]), .B2(n10038), .ZN(n9326) );
  AOI22D1BWP30P140LVT U13616 ( .A1(i_data_bus[187]), .A2(n10040), .B1(
        i_data_bus[219]), .B2(n10039), .ZN(n9325) );
  ND2D1BWP30P140LVT U13617 ( .A1(n9326), .A2(n9325), .ZN(N8986) );
  AOI22D1BWP30P140LVT U13618 ( .A1(i_data_bus[350]), .A2(n9731), .B1(
        i_data_bus[318]), .B2(n9732), .ZN(n9328) );
  AOI22D1BWP30P140LVT U13619 ( .A1(i_data_bus[286]), .A2(n6219), .B1(
        i_data_bus[382]), .B2(n9730), .ZN(n9327) );
  ND2D1BWP30P140LVT U13620 ( .A1(n9328), .A2(n9327), .ZN(N3757) );
  AOI22D1BWP30P140LVT U13621 ( .A1(i_data_bus[311]), .A2(n9732), .B1(
        i_data_bus[343]), .B2(n9731), .ZN(n9330) );
  AOI22D1BWP30P140LVT U13622 ( .A1(i_data_bus[279]), .A2(n6219), .B1(
        i_data_bus[375]), .B2(n9730), .ZN(n9329) );
  ND2D1BWP30P140LVT U13623 ( .A1(n9330), .A2(n9329), .ZN(N3750) );
  AOI22D1BWP30P140LVT U13624 ( .A1(i_data_bus[278]), .A2(n6219), .B1(
        i_data_bus[342]), .B2(n9731), .ZN(n9332) );
  AOI22D1BWP30P140LVT U13625 ( .A1(i_data_bus[310]), .A2(n9732), .B1(
        i_data_bus[374]), .B2(n9730), .ZN(n9331) );
  ND2D1BWP30P140LVT U13626 ( .A1(n9332), .A2(n9331), .ZN(N3749) );
  AOI22D1BWP30P140LVT U13627 ( .A1(i_data_bus[339]), .A2(n9731), .B1(
        i_data_bus[307]), .B2(n9732), .ZN(n9334) );
  AOI22D1BWP30P140LVT U13628 ( .A1(i_data_bus[275]), .A2(n6219), .B1(
        i_data_bus[371]), .B2(n9730), .ZN(n9333) );
  ND2D1BWP30P140LVT U13629 ( .A1(n9334), .A2(n9333), .ZN(N3746) );
  AOI22D1BWP30P140LVT U13630 ( .A1(i_data_bus[304]), .A2(n9732), .B1(
        i_data_bus[336]), .B2(n9731), .ZN(n9336) );
  AOI22D1BWP30P140LVT U13631 ( .A1(i_data_bus[272]), .A2(n6219), .B1(
        i_data_bus[368]), .B2(n9730), .ZN(n9335) );
  ND2D1BWP30P140LVT U13632 ( .A1(n9336), .A2(n9335), .ZN(N3743) );
  AOI22D1BWP30P140LVT U13633 ( .A1(i_data_bus[302]), .A2(n9732), .B1(
        i_data_bus[334]), .B2(n9731), .ZN(n9338) );
  AOI22D1BWP30P140LVT U13634 ( .A1(i_data_bus[270]), .A2(n6219), .B1(
        i_data_bus[366]), .B2(n9730), .ZN(n9337) );
  ND2D1BWP30P140LVT U13635 ( .A1(n9338), .A2(n9337), .ZN(N3741) );
  AOI22D1BWP30P140LVT U13636 ( .A1(i_data_bus[266]), .A2(n6219), .B1(
        i_data_bus[298]), .B2(n9732), .ZN(n9340) );
  AOI22D1BWP30P140LVT U13637 ( .A1(i_data_bus[330]), .A2(n9731), .B1(
        i_data_bus[362]), .B2(n9730), .ZN(n9339) );
  ND2D1BWP30P140LVT U13638 ( .A1(n9340), .A2(n9339), .ZN(N3737) );
  AOI22D1BWP30P140LVT U13639 ( .A1(i_data_bus[263]), .A2(n6219), .B1(
        i_data_bus[327]), .B2(n9731), .ZN(n9342) );
  AOI22D1BWP30P140LVT U13640 ( .A1(i_data_bus[295]), .A2(n9732), .B1(
        i_data_bus[359]), .B2(n9730), .ZN(n9341) );
  ND2D1BWP30P140LVT U13641 ( .A1(n9342), .A2(n9341), .ZN(N3734) );
  AOI22D1BWP30P140LVT U13642 ( .A1(i_data_bus[260]), .A2(n6219), .B1(
        i_data_bus[324]), .B2(n9731), .ZN(n9344) );
  AOI22D1BWP30P140LVT U13643 ( .A1(i_data_bus[292]), .A2(n9732), .B1(
        i_data_bus[356]), .B2(n9730), .ZN(n9343) );
  ND2D1BWP30P140LVT U13644 ( .A1(n9344), .A2(n9343), .ZN(N3731) );
  AOI22D1BWP30P140LVT U13645 ( .A1(i_data_bus[290]), .A2(n9732), .B1(
        i_data_bus[258]), .B2(n6219), .ZN(n9346) );
  AOI22D1BWP30P140LVT U13646 ( .A1(i_data_bus[322]), .A2(n9731), .B1(
        i_data_bus[354]), .B2(n9730), .ZN(n9345) );
  ND2D1BWP30P140LVT U13647 ( .A1(n9346), .A2(n9345), .ZN(N3729) );
  AOI22D1BWP30P140LVT U13648 ( .A1(i_data_bus[321]), .A2(n9731), .B1(
        i_data_bus[257]), .B2(n6219), .ZN(n9348) );
  AOI22D1BWP30P140LVT U13649 ( .A1(i_data_bus[289]), .A2(n9732), .B1(
        i_data_bus[353]), .B2(n9730), .ZN(n9347) );
  ND2D1BWP30P140LVT U13650 ( .A1(n9348), .A2(n9347), .ZN(N3728) );
  AOI22D1BWP30P140LVT U13651 ( .A1(i_data_bus[628]), .A2(n10254), .B1(
        i_data_bus[564]), .B2(n10253), .ZN(n9350) );
  AOI22D1BWP30P140LVT U13652 ( .A1(i_data_bus[596]), .A2(n10252), .B1(
        i_data_bus[532]), .B2(n10245), .ZN(n9349) );
  ND2D1BWP30P140LVT U13653 ( .A1(n9350), .A2(n9349), .ZN(N9627) );
  AOI22D1BWP30P140LVT U13654 ( .A1(i_data_bus[530]), .A2(n10245), .B1(
        i_data_bus[562]), .B2(n10253), .ZN(n9352) );
  AOI22D1BWP30P140LVT U13655 ( .A1(i_data_bus[594]), .A2(n10252), .B1(
        i_data_bus[626]), .B2(n10254), .ZN(n9351) );
  ND2D1BWP30P140LVT U13656 ( .A1(n9352), .A2(n9351), .ZN(N9625) );
  AOI22D1BWP30P140LVT U13657 ( .A1(i_data_bus[543]), .A2(n10245), .B1(
        i_data_bus[575]), .B2(n10253), .ZN(n9354) );
  AOI22D1BWP30P140LVT U13658 ( .A1(i_data_bus[607]), .A2(n10252), .B1(
        i_data_bus[639]), .B2(n10254), .ZN(n9353) );
  ND2D1BWP30P140LVT U13659 ( .A1(n9354), .A2(n9353), .ZN(N9638) );
  AOI22D1BWP30P140LVT U13660 ( .A1(i_data_bus[517]), .A2(n10245), .B1(
        i_data_bus[549]), .B2(n10253), .ZN(n9356) );
  AOI22D1BWP30P140LVT U13661 ( .A1(i_data_bus[581]), .A2(n10252), .B1(
        i_data_bus[613]), .B2(n10254), .ZN(n9355) );
  ND2D1BWP30P140LVT U13662 ( .A1(n9356), .A2(n9355), .ZN(N9612) );
  AOI22D1BWP30P140LVT U13663 ( .A1(i_data_bus[633]), .A2(n10254), .B1(
        i_data_bus[569]), .B2(n10253), .ZN(n9358) );
  AOI22D1BWP30P140LVT U13664 ( .A1(i_data_bus[537]), .A2(n10245), .B1(
        i_data_bus[601]), .B2(n10252), .ZN(n9357) );
  ND2D1BWP30P140LVT U13665 ( .A1(n9358), .A2(n9357), .ZN(N9632) );
  AOI22D1BWP30P140LVT U13666 ( .A1(i_data_bus[525]), .A2(n10245), .B1(
        i_data_bus[557]), .B2(n10253), .ZN(n9360) );
  AOI22D1BWP30P140LVT U13667 ( .A1(i_data_bus[621]), .A2(n10254), .B1(
        i_data_bus[589]), .B2(n10252), .ZN(n9359) );
  ND2D1BWP30P140LVT U13668 ( .A1(n9360), .A2(n9359), .ZN(N9620) );
  AOI22D1BWP30P140LVT U13669 ( .A1(i_data_bus[630]), .A2(n10254), .B1(
        i_data_bus[566]), .B2(n10253), .ZN(n9362) );
  AOI22D1BWP30P140LVT U13670 ( .A1(i_data_bus[534]), .A2(n10245), .B1(
        i_data_bus[598]), .B2(n10252), .ZN(n9361) );
  ND2D1BWP30P140LVT U13671 ( .A1(n9362), .A2(n9361), .ZN(N9629) );
  AOI22D1BWP30P140LVT U13672 ( .A1(i_data_bus[606]), .A2(n10269), .B1(
        i_data_bus[574]), .B2(n10271), .ZN(n9364) );
  AOI22D1BWP30P140LVT U13673 ( .A1(i_data_bus[638]), .A2(n10270), .B1(
        i_data_bus[542]), .B2(n10272), .ZN(n9363) );
  ND2D1BWP30P140LVT U13674 ( .A1(n9364), .A2(n9363), .ZN(N8147) );
  AOI22D1BWP30P140LVT U13675 ( .A1(i_data_bus[579]), .A2(n10269), .B1(
        i_data_bus[547]), .B2(n10271), .ZN(n9366) );
  AOI22D1BWP30P140LVT U13676 ( .A1(i_data_bus[611]), .A2(n10270), .B1(
        i_data_bus[515]), .B2(n10272), .ZN(n9365) );
  ND2D1BWP30P140LVT U13677 ( .A1(n9366), .A2(n9365), .ZN(N8120) );
  AOI22D1BWP30P140LVT U13678 ( .A1(i_data_bus[530]), .A2(n10272), .B1(
        i_data_bus[562]), .B2(n10271), .ZN(n9368) );
  AOI22D1BWP30P140LVT U13679 ( .A1(i_data_bus[594]), .A2(n10269), .B1(
        i_data_bus[626]), .B2(n10270), .ZN(n9367) );
  ND2D1BWP30P140LVT U13680 ( .A1(n9368), .A2(n9367), .ZN(N8135) );
  AOI22D1BWP30P140LVT U13681 ( .A1(i_data_bus[520]), .A2(n10272), .B1(
        i_data_bus[552]), .B2(n10271), .ZN(n9370) );
  AOI22D1BWP30P140LVT U13682 ( .A1(i_data_bus[584]), .A2(n10269), .B1(
        i_data_bus[616]), .B2(n10270), .ZN(n9369) );
  ND2D1BWP30P140LVT U13683 ( .A1(n9370), .A2(n9369), .ZN(N8125) );
  AOI22D1BWP30P140LVT U13684 ( .A1(i_data_bus[543]), .A2(n10272), .B1(
        i_data_bus[575]), .B2(n10271), .ZN(n9372) );
  AOI22D1BWP30P140LVT U13685 ( .A1(i_data_bus[607]), .A2(n10269), .B1(
        i_data_bus[639]), .B2(n10270), .ZN(n9371) );
  ND2D1BWP30P140LVT U13686 ( .A1(n9372), .A2(n9371), .ZN(N8148) );
  AOI22D1BWP30P140LVT U13687 ( .A1(i_data_bus[571]), .A2(n10184), .B1(
        i_data_bus[603]), .B2(n10183), .ZN(n9374) );
  AOI22D1BWP30P140LVT U13688 ( .A1(i_data_bus[539]), .A2(n10182), .B1(
        i_data_bus[635]), .B2(n10185), .ZN(n9373) );
  ND2D1BWP30P140LVT U13689 ( .A1(n9374), .A2(n9373), .ZN(N6910) );
  AOI22D1BWP30P140LVT U13690 ( .A1(i_data_bus[522]), .A2(n10182), .B1(
        i_data_bus[554]), .B2(n10184), .ZN(n9376) );
  AOI22D1BWP30P140LVT U13691 ( .A1(i_data_bus[586]), .A2(n10183), .B1(
        i_data_bus[618]), .B2(n10185), .ZN(n9375) );
  ND2D1BWP30P140LVT U13692 ( .A1(n9376), .A2(n9375), .ZN(N6893) );
  AOI22D1BWP30P140LVT U13693 ( .A1(i_data_bus[529]), .A2(n10182), .B1(
        i_data_bus[593]), .B2(n10183), .ZN(n9378) );
  AOI22D1BWP30P140LVT U13694 ( .A1(i_data_bus[561]), .A2(n10184), .B1(
        i_data_bus[625]), .B2(n10185), .ZN(n9377) );
  ND2D1BWP30P140LVT U13695 ( .A1(n9378), .A2(n9377), .ZN(N6900) );
  AOI22D1BWP30P140LVT U13696 ( .A1(i_data_bus[521]), .A2(n10182), .B1(
        i_data_bus[553]), .B2(n10184), .ZN(n9380) );
  AOI22D1BWP30P140LVT U13697 ( .A1(i_data_bus[585]), .A2(n10183), .B1(
        i_data_bus[617]), .B2(n10185), .ZN(n9379) );
  ND2D1BWP30P140LVT U13698 ( .A1(n9380), .A2(n9379), .ZN(N6892) );
  AOI22D1BWP30P140LVT U13699 ( .A1(i_data_bus[637]), .A2(n10270), .B1(
        i_data_bus[573]), .B2(n10271), .ZN(n9382) );
  AOI22D1BWP30P140LVT U13700 ( .A1(i_data_bus[541]), .A2(n10272), .B1(
        i_data_bus[605]), .B2(n10269), .ZN(n9381) );
  ND2D1BWP30P140LVT U13701 ( .A1(n9382), .A2(n9381), .ZN(N8146) );
  AOI22D1BWP30P140LVT U13702 ( .A1(i_data_bus[538]), .A2(n10272), .B1(
        i_data_bus[570]), .B2(n10271), .ZN(n9384) );
  AOI22D1BWP30P140LVT U13703 ( .A1(i_data_bus[634]), .A2(n10270), .B1(
        i_data_bus[602]), .B2(n10269), .ZN(n9383) );
  ND2D1BWP30P140LVT U13704 ( .A1(n9384), .A2(n9383), .ZN(N8143) );
  AOI22D1BWP30P140LVT U13705 ( .A1(i_data_bus[633]), .A2(n10270), .B1(
        i_data_bus[569]), .B2(n10271), .ZN(n9386) );
  AOI22D1BWP30P140LVT U13706 ( .A1(i_data_bus[537]), .A2(n10272), .B1(
        i_data_bus[601]), .B2(n10269), .ZN(n9385) );
  ND2D1BWP30P140LVT U13707 ( .A1(n9386), .A2(n9385), .ZN(N8142) );
  AOI22D1BWP30P140LVT U13708 ( .A1(i_data_bus[630]), .A2(n10270), .B1(
        i_data_bus[566]), .B2(n10271), .ZN(n9388) );
  AOI22D1BWP30P140LVT U13709 ( .A1(i_data_bus[534]), .A2(n10272), .B1(
        i_data_bus[598]), .B2(n10269), .ZN(n9387) );
  ND2D1BWP30P140LVT U13710 ( .A1(n9388), .A2(n9387), .ZN(N8139) );
  AOI22D1BWP30P140LVT U13711 ( .A1(i_data_bus[629]), .A2(n10270), .B1(
        i_data_bus[565]), .B2(n10271), .ZN(n9390) );
  AOI22D1BWP30P140LVT U13712 ( .A1(i_data_bus[533]), .A2(n10272), .B1(
        i_data_bus[597]), .B2(n10269), .ZN(n9389) );
  ND2D1BWP30P140LVT U13713 ( .A1(n9390), .A2(n9389), .ZN(N8138) );
  AOI22D1BWP30P140LVT U13714 ( .A1(i_data_bus[525]), .A2(n10272), .B1(
        i_data_bus[557]), .B2(n10271), .ZN(n9392) );
  AOI22D1BWP30P140LVT U13715 ( .A1(i_data_bus[621]), .A2(n10270), .B1(
        i_data_bus[589]), .B2(n10269), .ZN(n9391) );
  ND2D1BWP30P140LVT U13716 ( .A1(n9392), .A2(n9391), .ZN(N8130) );
  AOI22D1BWP30P140LVT U13717 ( .A1(i_data_bus[518]), .A2(n10272), .B1(
        i_data_bus[550]), .B2(n10271), .ZN(n9394) );
  AOI22D1BWP30P140LVT U13718 ( .A1(i_data_bus[614]), .A2(n10270), .B1(
        i_data_bus[582]), .B2(n10269), .ZN(n9393) );
  ND2D1BWP30P140LVT U13719 ( .A1(n9394), .A2(n9393), .ZN(N8123) );
  AOI22D1BWP30P140LVT U13720 ( .A1(i_data_bus[570]), .A2(n9935), .B1(
        i_data_bus[602]), .B2(n9936), .ZN(n9396) );
  AOI22D1BWP30P140LVT U13721 ( .A1(i_data_bus[538]), .A2(n9934), .B1(
        i_data_bus[634]), .B2(n9933), .ZN(n9395) );
  ND2D1BWP30P140LVT U13722 ( .A1(n9396), .A2(n9395), .ZN(N5419) );
  AOI22D1BWP30P140LVT U13723 ( .A1(i_data_bus[563]), .A2(n9935), .B1(
        i_data_bus[595]), .B2(n9936), .ZN(n9398) );
  AOI22D1BWP30P140LVT U13724 ( .A1(i_data_bus[531]), .A2(n9934), .B1(
        i_data_bus[627]), .B2(n9933), .ZN(n9397) );
  ND2D1BWP30P140LVT U13725 ( .A1(n9398), .A2(n9397), .ZN(N5412) );
  AOI22D1BWP30P140LVT U13726 ( .A1(i_data_bus[529]), .A2(n9934), .B1(
        i_data_bus[593]), .B2(n9936), .ZN(n9400) );
  AOI22D1BWP30P140LVT U13727 ( .A1(i_data_bus[561]), .A2(n9935), .B1(
        i_data_bus[625]), .B2(n9933), .ZN(n9399) );
  ND2D1BWP30P140LVT U13728 ( .A1(n9400), .A2(n9399), .ZN(N5410) );
  AOI22D1BWP30P140LVT U13729 ( .A1(i_data_bus[521]), .A2(n9934), .B1(
        i_data_bus[553]), .B2(n9935), .ZN(n9402) );
  AOI22D1BWP30P140LVT U13730 ( .A1(i_data_bus[585]), .A2(n9936), .B1(
        i_data_bus[617]), .B2(n9933), .ZN(n9401) );
  ND2D1BWP30P140LVT U13731 ( .A1(n9402), .A2(n9401), .ZN(N5402) );
  AOI22D1BWP30P140LVT U13732 ( .A1(i_data_bus[516]), .A2(n9934), .B1(
        i_data_bus[580]), .B2(n9936), .ZN(n9404) );
  AOI22D1BWP30P140LVT U13733 ( .A1(i_data_bus[548]), .A2(n9935), .B1(
        i_data_bus[612]), .B2(n9933), .ZN(n9403) );
  ND2D1BWP30P140LVT U13734 ( .A1(n9404), .A2(n9403), .ZN(N5397) );
  AOI22D1BWP30P140LVT U13735 ( .A1(i_data_bus[45]), .A2(n10087), .B1(
        i_data_bus[109]), .B2(n10085), .ZN(n9406) );
  AOI22D1BWP30P140LVT U13736 ( .A1(i_data_bus[13]), .A2(n10088), .B1(
        i_data_bus[77]), .B2(n10086), .ZN(n9405) );
  ND2D1BWP30P140LVT U13737 ( .A1(n9406), .A2(n9405), .ZN(N5054) );
  AOI22D1BWP30P140LVT U13738 ( .A1(i_data_bus[103]), .A2(n10117), .B1(
        i_data_bus[39]), .B2(n10118), .ZN(n9408) );
  AOI22D1BWP30P140LVT U13739 ( .A1(i_data_bus[7]), .A2(n10116), .B1(
        i_data_bus[71]), .B2(n10115), .ZN(n9407) );
  ND2D1BWP30P140LVT U13740 ( .A1(n9408), .A2(n9407), .ZN(N7772) );
  AOI22D1BWP30P140LVT U13741 ( .A1(i_data_bus[56]), .A2(n9977), .B1(
        i_data_bus[120]), .B2(n9978), .ZN(n9410) );
  AOI22D1BWP30P140LVT U13742 ( .A1(i_data_bus[24]), .A2(n9969), .B1(
        i_data_bus[88]), .B2(n9976), .ZN(n9409) );
  ND2D1BWP30P140LVT U13743 ( .A1(n9410), .A2(n9409), .ZN(N2341) );
  AOI22D1BWP30P140LVT U13744 ( .A1(i_data_bus[51]), .A2(n9977), .B1(
        i_data_bus[115]), .B2(n9978), .ZN(n9412) );
  AOI22D1BWP30P140LVT U13745 ( .A1(i_data_bus[19]), .A2(n9969), .B1(
        i_data_bus[83]), .B2(n9976), .ZN(n9411) );
  ND2D1BWP30P140LVT U13746 ( .A1(n9412), .A2(n9411), .ZN(N2336) );
  AOI22D1BWP30P140LVT U13747 ( .A1(i_data_bus[139]), .A2(n9522), .B1(
        i_data_bus[235]), .B2(n9520), .ZN(n9414) );
  AOI22D1BWP30P140LVT U13748 ( .A1(i_data_bus[171]), .A2(n9519), .B1(
        i_data_bus[203]), .B2(n9521), .ZN(n9413) );
  ND2D1BWP30P140LVT U13749 ( .A1(n9414), .A2(n9413), .ZN(N5140) );
  AOI22D1BWP30P140LVT U13750 ( .A1(i_data_bus[98]), .A2(n10085), .B1(
        i_data_bus[2]), .B2(n10088), .ZN(n9416) );
  AOI22D1BWP30P140LVT U13751 ( .A1(i_data_bus[34]), .A2(n10087), .B1(
        i_data_bus[66]), .B2(n10086), .ZN(n9415) );
  ND2D1BWP30P140LVT U13752 ( .A1(n9416), .A2(n9415), .ZN(N5043) );
  AOI22D1BWP30P140LVT U13753 ( .A1(i_data_bus[278]), .A2(n6227), .B1(
        i_data_bus[374]), .B2(n10277), .ZN(n9418) );
  AOI22D1BWP30P140LVT U13754 ( .A1(i_data_bus[310]), .A2(n10276), .B1(
        i_data_bus[342]), .B2(n10275), .ZN(n9417) );
  ND2D1BWP30P140LVT U13755 ( .A1(n9418), .A2(n9417), .ZN(N9197) );
  AOI22D1BWP30P140LVT U13756 ( .A1(i_data_bus[98]), .A2(n10117), .B1(
        i_data_bus[2]), .B2(n10116), .ZN(n9420) );
  AOI22D1BWP30P140LVT U13757 ( .A1(i_data_bus[34]), .A2(n10118), .B1(
        i_data_bus[66]), .B2(n10115), .ZN(n9419) );
  ND2D1BWP30P140LVT U13758 ( .A1(n9420), .A2(n9419), .ZN(N7767) );
  AOI22D1BWP30P140LVT U13759 ( .A1(i_data_bus[103]), .A2(n9978), .B1(
        i_data_bus[39]), .B2(n9977), .ZN(n9422) );
  AOI22D1BWP30P140LVT U13760 ( .A1(i_data_bus[7]), .A2(n9969), .B1(
        i_data_bus[71]), .B2(n9976), .ZN(n9421) );
  ND2D1BWP30P140LVT U13761 ( .A1(n9422), .A2(n9421), .ZN(N2324) );
  AOI22D1BWP30P140LVT U13762 ( .A1(i_data_bus[102]), .A2(n9978), .B1(
        i_data_bus[38]), .B2(n9977), .ZN(n9424) );
  AOI22D1BWP30P140LVT U13763 ( .A1(i_data_bus[6]), .A2(n9969), .B1(
        i_data_bus[70]), .B2(n9976), .ZN(n9423) );
  ND2D1BWP30P140LVT U13764 ( .A1(n9424), .A2(n9423), .ZN(N2323) );
  AOI22D1BWP30P140LVT U13765 ( .A1(i_data_bus[5]), .A2(n9969), .B1(
        i_data_bus[37]), .B2(n9977), .ZN(n9426) );
  AOI22D1BWP30P140LVT U13766 ( .A1(i_data_bus[101]), .A2(n9978), .B1(
        i_data_bus[69]), .B2(n9976), .ZN(n9425) );
  ND2D1BWP30P140LVT U13767 ( .A1(n9426), .A2(n9425), .ZN(N2322) );
  AOI22D1BWP30P140LVT U13768 ( .A1(i_data_bus[28]), .A2(n10116), .B1(
        i_data_bus[124]), .B2(n10117), .ZN(n9428) );
  AOI22D1BWP30P140LVT U13769 ( .A1(i_data_bus[60]), .A2(n10118), .B1(
        i_data_bus[92]), .B2(n10115), .ZN(n9427) );
  ND2D1BWP30P140LVT U13770 ( .A1(n9428), .A2(n9427), .ZN(N7793) );
  AOI22D1BWP30P140LVT U13771 ( .A1(i_data_bus[34]), .A2(n9977), .B1(
        i_data_bus[2]), .B2(n9969), .ZN(n9430) );
  AOI22D1BWP30P140LVT U13772 ( .A1(i_data_bus[98]), .A2(n9978), .B1(
        i_data_bus[66]), .B2(n9976), .ZN(n9429) );
  ND2D1BWP30P140LVT U13773 ( .A1(n9430), .A2(n9429), .ZN(N2319) );
  AOI22D1BWP30P140LVT U13774 ( .A1(i_data_bus[35]), .A2(n9977), .B1(
        i_data_bus[3]), .B2(n9969), .ZN(n9432) );
  AOI22D1BWP30P140LVT U13775 ( .A1(i_data_bus[99]), .A2(n9978), .B1(
        i_data_bus[67]), .B2(n9976), .ZN(n9431) );
  ND2D1BWP30P140LVT U13776 ( .A1(n9432), .A2(n9431), .ZN(N2320) );
  AOI22D1BWP30P140LVT U13777 ( .A1(i_data_bus[1]), .A2(n9969), .B1(
        i_data_bus[33]), .B2(n9977), .ZN(n9434) );
  AOI22D1BWP30P140LVT U13778 ( .A1(i_data_bus[97]), .A2(n9978), .B1(
        i_data_bus[65]), .B2(n9976), .ZN(n9433) );
  ND2D1BWP30P140LVT U13779 ( .A1(n9434), .A2(n9433), .ZN(N2318) );
  AOI22D1BWP30P140LVT U13780 ( .A1(i_data_bus[155]), .A2(n6213), .B1(
        i_data_bus[251]), .B2(n10220), .ZN(n9436) );
  AOI22D1BWP30P140LVT U13781 ( .A1(i_data_bus[187]), .A2(n10219), .B1(
        i_data_bus[219]), .B2(n10218), .ZN(n9435) );
  ND2D1BWP30P140LVT U13782 ( .A1(n9436), .A2(n9435), .ZN(N2432) );
  AOI22D1BWP30P140LVT U13783 ( .A1(i_data_bus[153]), .A2(n6213), .B1(
        i_data_bus[185]), .B2(n10219), .ZN(n9438) );
  AOI22D1BWP30P140LVT U13784 ( .A1(i_data_bus[249]), .A2(n10220), .B1(
        i_data_bus[217]), .B2(n10218), .ZN(n9437) );
  ND2D1BWP30P140LVT U13785 ( .A1(n9438), .A2(n9437), .ZN(N2430) );
  AOI22D1BWP30P140LVT U13786 ( .A1(i_data_bus[30]), .A2(n9969), .B1(
        i_data_bus[126]), .B2(n9978), .ZN(n9440) );
  AOI22D1BWP30P140LVT U13787 ( .A1(i_data_bus[62]), .A2(n9977), .B1(
        i_data_bus[94]), .B2(n9976), .ZN(n9439) );
  ND2D1BWP30P140LVT U13788 ( .A1(n9440), .A2(n9439), .ZN(N2347) );
  AOI22D1BWP30P140LVT U13789 ( .A1(i_data_bus[174]), .A2(n10219), .B1(
        i_data_bus[238]), .B2(n10220), .ZN(n9442) );
  AOI22D1BWP30P140LVT U13790 ( .A1(i_data_bus[142]), .A2(n6213), .B1(
        i_data_bus[206]), .B2(n10218), .ZN(n9441) );
  ND2D1BWP30P140LVT U13791 ( .A1(n9442), .A2(n9441), .ZN(N2419) );
  AOI22D1BWP30P140LVT U13792 ( .A1(i_data_bus[139]), .A2(n6213), .B1(
        i_data_bus[171]), .B2(n10219), .ZN(n9444) );
  AOI22D1BWP30P140LVT U13793 ( .A1(i_data_bus[235]), .A2(n10220), .B1(
        i_data_bus[203]), .B2(n10218), .ZN(n9443) );
  ND2D1BWP30P140LVT U13794 ( .A1(n9444), .A2(n9443), .ZN(N2416) );
  AOI22D1BWP30P140LVT U13795 ( .A1(i_data_bus[138]), .A2(n6213), .B1(
        i_data_bus[234]), .B2(n10220), .ZN(n9446) );
  AOI22D1BWP30P140LVT U13796 ( .A1(i_data_bus[170]), .A2(n10219), .B1(
        i_data_bus[202]), .B2(n10218), .ZN(n9445) );
  ND2D1BWP30P140LVT U13797 ( .A1(n9446), .A2(n9445), .ZN(N2415) );
  AOI22D1BWP30P140LVT U13798 ( .A1(i_data_bus[230]), .A2(n10220), .B1(
        i_data_bus[166]), .B2(n10219), .ZN(n9448) );
  AOI22D1BWP30P140LVT U13799 ( .A1(i_data_bus[134]), .A2(n6213), .B1(
        i_data_bus[198]), .B2(n10218), .ZN(n9447) );
  ND2D1BWP30P140LVT U13800 ( .A1(n9448), .A2(n9447), .ZN(N2411) );
  AOI22D1BWP30P140LVT U13801 ( .A1(i_data_bus[226]), .A2(n10220), .B1(
        i_data_bus[130]), .B2(n6213), .ZN(n9450) );
  AOI22D1BWP30P140LVT U13802 ( .A1(i_data_bus[162]), .A2(n10219), .B1(
        i_data_bus[194]), .B2(n10218), .ZN(n9449) );
  ND2D1BWP30P140LVT U13803 ( .A1(n9450), .A2(n9449), .ZN(N2407) );
  AOI22D1BWP30P140LVT U13804 ( .A1(i_data_bus[160]), .A2(n10219), .B1(
        i_data_bus[128]), .B2(n6213), .ZN(n9452) );
  AOI22D1BWP30P140LVT U13805 ( .A1(i_data_bus[224]), .A2(n10220), .B1(
        i_data_bus[192]), .B2(n10218), .ZN(n9451) );
  ND2D1BWP30P140LVT U13806 ( .A1(n9452), .A2(n9451), .ZN(N2405) );
  AOI22D1BWP30P140LVT U13807 ( .A1(i_data_bus[113]), .A2(n10117), .B1(
        i_data_bus[49]), .B2(n10118), .ZN(n9454) );
  AOI22D1BWP30P140LVT U13808 ( .A1(i_data_bus[17]), .A2(n10116), .B1(
        i_data_bus[81]), .B2(n10115), .ZN(n9453) );
  ND2D1BWP30P140LVT U13809 ( .A1(n9454), .A2(n9453), .ZN(N7782) );
  AOI22D1BWP30P140LVT U13810 ( .A1(i_data_bus[97]), .A2(n10117), .B1(
        i_data_bus[33]), .B2(n10118), .ZN(n9456) );
  AOI22D1BWP30P140LVT U13811 ( .A1(i_data_bus[1]), .A2(n10116), .B1(
        i_data_bus[65]), .B2(n10115), .ZN(n9455) );
  ND2D1BWP30P140LVT U13812 ( .A1(n9456), .A2(n9455), .ZN(N7766) );
  AOI22D1BWP30P140LVT U13813 ( .A1(i_data_bus[136]), .A2(n9522), .B1(
        i_data_bus[232]), .B2(n9520), .ZN(n9458) );
  AOI22D1BWP30P140LVT U13814 ( .A1(i_data_bus[168]), .A2(n9519), .B1(
        i_data_bus[200]), .B2(n9521), .ZN(n9457) );
  ND2D1BWP30P140LVT U13815 ( .A1(n9458), .A2(n9457), .ZN(N5137) );
  AOI22D1BWP30P140LVT U13816 ( .A1(i_data_bus[21]), .A2(n9969), .B1(
        i_data_bus[53]), .B2(n9977), .ZN(n9460) );
  AOI22D1BWP30P140LVT U13817 ( .A1(i_data_bus[117]), .A2(n9978), .B1(
        i_data_bus[85]), .B2(n9976), .ZN(n9459) );
  ND2D1BWP30P140LVT U13818 ( .A1(n9460), .A2(n9459), .ZN(N2338) );
  AOI22D1BWP30P140LVT U13819 ( .A1(i_data_bus[48]), .A2(n10118), .B1(
        i_data_bus[112]), .B2(n10117), .ZN(n9462) );
  AOI22D1BWP30P140LVT U13820 ( .A1(i_data_bus[16]), .A2(n10116), .B1(
        i_data_bus[80]), .B2(n10115), .ZN(n9461) );
  ND2D1BWP30P140LVT U13821 ( .A1(n9462), .A2(n9461), .ZN(N7781) );
  AOI22D1BWP30P140LVT U13822 ( .A1(i_data_bus[279]), .A2(n6227), .B1(
        i_data_bus[311]), .B2(n10276), .ZN(n9464) );
  AOI22D1BWP30P140LVT U13823 ( .A1(i_data_bus[375]), .A2(n10277), .B1(
        i_data_bus[343]), .B2(n10275), .ZN(n9463) );
  ND2D1BWP30P140LVT U13824 ( .A1(n9464), .A2(n9463), .ZN(N9198) );
  AOI22D1BWP30P140LVT U13825 ( .A1(i_data_bus[56]), .A2(n10118), .B1(
        i_data_bus[120]), .B2(n10117), .ZN(n9466) );
  AOI22D1BWP30P140LVT U13826 ( .A1(i_data_bus[24]), .A2(n10116), .B1(
        i_data_bus[88]), .B2(n10115), .ZN(n9465) );
  ND2D1BWP30P140LVT U13827 ( .A1(n9466), .A2(n9465), .ZN(N7789) );
  AOI22D1BWP30P140LVT U13828 ( .A1(i_data_bus[268]), .A2(n6227), .B1(
        i_data_bus[300]), .B2(n10276), .ZN(n9468) );
  AOI22D1BWP30P140LVT U13829 ( .A1(i_data_bus[364]), .A2(n10277), .B1(
        i_data_bus[332]), .B2(n10275), .ZN(n9467) );
  ND2D1BWP30P140LVT U13830 ( .A1(n9468), .A2(n9467), .ZN(N9187) );
  AOI22D1BWP30P140LVT U13831 ( .A1(i_data_bus[316]), .A2(n10276), .B1(
        i_data_bus[380]), .B2(n10277), .ZN(n9470) );
  AOI22D1BWP30P140LVT U13832 ( .A1(i_data_bus[284]), .A2(n6227), .B1(
        i_data_bus[348]), .B2(n10275), .ZN(n9469) );
  ND2D1BWP30P140LVT U13833 ( .A1(n9470), .A2(n9469), .ZN(N9203) );
  AOI22D1BWP30P140LVT U13834 ( .A1(i_data_bus[357]), .A2(n10277), .B1(
        i_data_bus[293]), .B2(n10276), .ZN(n9472) );
  AOI22D1BWP30P140LVT U13835 ( .A1(i_data_bus[261]), .A2(n6227), .B1(
        i_data_bus[325]), .B2(n10275), .ZN(n9471) );
  ND2D1BWP30P140LVT U13836 ( .A1(n9472), .A2(n9471), .ZN(N9180) );
  AOI22D1BWP30P140LVT U13837 ( .A1(i_data_bus[30]), .A2(n10088), .B1(
        i_data_bus[126]), .B2(n10085), .ZN(n9474) );
  AOI22D1BWP30P140LVT U13838 ( .A1(i_data_bus[62]), .A2(n10087), .B1(
        i_data_bus[94]), .B2(n10086), .ZN(n9473) );
  ND2D1BWP30P140LVT U13839 ( .A1(n9474), .A2(n9473), .ZN(N5071) );
  AOI22D1BWP30P140LVT U13840 ( .A1(i_data_bus[11]), .A2(n10116), .B1(
        i_data_bus[43]), .B2(n10118), .ZN(n9476) );
  AOI22D1BWP30P140LVT U13841 ( .A1(i_data_bus[107]), .A2(n10117), .B1(
        i_data_bus[75]), .B2(n10115), .ZN(n9475) );
  ND2D1BWP30P140LVT U13842 ( .A1(n9476), .A2(n9475), .ZN(N7776) );
  AOI22D1BWP30P140LVT U13843 ( .A1(i_data_bus[123]), .A2(n10085), .B1(
        i_data_bus[59]), .B2(n10087), .ZN(n9478) );
  AOI22D1BWP30P140LVT U13844 ( .A1(i_data_bus[27]), .A2(n10088), .B1(
        i_data_bus[91]), .B2(n10086), .ZN(n9477) );
  ND2D1BWP30P140LVT U13845 ( .A1(n9478), .A2(n9477), .ZN(N5068) );
  AOI22D1BWP30P140LVT U13846 ( .A1(i_data_bus[25]), .A2(n10088), .B1(
        i_data_bus[57]), .B2(n10087), .ZN(n9480) );
  AOI22D1BWP30P140LVT U13847 ( .A1(i_data_bus[121]), .A2(n10085), .B1(
        i_data_bus[89]), .B2(n10086), .ZN(n9479) );
  ND2D1BWP30P140LVT U13848 ( .A1(n9480), .A2(n9479), .ZN(N5066) );
  AOI22D1BWP30P140LVT U13849 ( .A1(i_data_bus[23]), .A2(n10088), .B1(
        i_data_bus[119]), .B2(n10085), .ZN(n9482) );
  AOI22D1BWP30P140LVT U13850 ( .A1(i_data_bus[55]), .A2(n10087), .B1(
        i_data_bus[87]), .B2(n10086), .ZN(n9481) );
  ND2D1BWP30P140LVT U13851 ( .A1(n9482), .A2(n9481), .ZN(N5064) );
  AOI22D1BWP30P140LVT U13852 ( .A1(i_data_bus[22]), .A2(n10088), .B1(
        i_data_bus[54]), .B2(n10087), .ZN(n9484) );
  AOI22D1BWP30P140LVT U13853 ( .A1(i_data_bus[118]), .A2(n10085), .B1(
        i_data_bus[86]), .B2(n10086), .ZN(n9483) );
  ND2D1BWP30P140LVT U13854 ( .A1(n9484), .A2(n9483), .ZN(N5063) );
  AOI22D1BWP30P140LVT U13855 ( .A1(i_data_bus[21]), .A2(n10088), .B1(
        i_data_bus[53]), .B2(n10087), .ZN(n9486) );
  AOI22D1BWP30P140LVT U13856 ( .A1(i_data_bus[117]), .A2(n10085), .B1(
        i_data_bus[85]), .B2(n10086), .ZN(n9485) );
  ND2D1BWP30P140LVT U13857 ( .A1(n9486), .A2(n9485), .ZN(N5062) );
  AOI22D1BWP30P140LVT U13858 ( .A1(i_data_bus[16]), .A2(n10088), .B1(
        i_data_bus[112]), .B2(n10085), .ZN(n9488) );
  AOI22D1BWP30P140LVT U13859 ( .A1(i_data_bus[48]), .A2(n10087), .B1(
        i_data_bus[80]), .B2(n10086), .ZN(n9487) );
  ND2D1BWP30P140LVT U13860 ( .A1(n9488), .A2(n9487), .ZN(N5057) );
  AOI22D1BWP30P140LVT U13861 ( .A1(i_data_bus[22]), .A2(n9969), .B1(
        i_data_bus[54]), .B2(n9977), .ZN(n9490) );
  AOI22D1BWP30P140LVT U13862 ( .A1(i_data_bus[118]), .A2(n9978), .B1(
        i_data_bus[86]), .B2(n9976), .ZN(n9489) );
  ND2D1BWP30P140LVT U13863 ( .A1(n9490), .A2(n9489), .ZN(N2339) );
  AOI22D1BWP30P140LVT U13864 ( .A1(i_data_bus[283]), .A2(n6227), .B1(
        i_data_bus[379]), .B2(n10277), .ZN(n9492) );
  AOI22D1BWP30P140LVT U13865 ( .A1(i_data_bus[315]), .A2(n10276), .B1(
        i_data_bus[347]), .B2(n10275), .ZN(n9491) );
  ND2D1BWP30P140LVT U13866 ( .A1(n9492), .A2(n9491), .ZN(N9202) );
  AOI22D1BWP30P140LVT U13867 ( .A1(i_data_bus[157]), .A2(n9522), .B1(
        i_data_bus[189]), .B2(n9519), .ZN(n9494) );
  AOI22D1BWP30P140LVT U13868 ( .A1(i_data_bus[253]), .A2(n9520), .B1(
        i_data_bus[221]), .B2(n9521), .ZN(n9493) );
  ND2D1BWP30P140LVT U13869 ( .A1(n9494), .A2(n9493), .ZN(N5158) );
  AOI22D1BWP30P140LVT U13870 ( .A1(i_data_bus[36]), .A2(n10118), .B1(
        i_data_bus[4]), .B2(n10116), .ZN(n9496) );
  AOI22D1BWP30P140LVT U13871 ( .A1(i_data_bus[100]), .A2(n10117), .B1(
        i_data_bus[68]), .B2(n10115), .ZN(n9495) );
  ND2D1BWP30P140LVT U13872 ( .A1(n9496), .A2(n9495), .ZN(N7769) );
  AOI22D1BWP30P140LVT U13873 ( .A1(i_data_bus[187]), .A2(n9519), .B1(
        i_data_bus[251]), .B2(n9520), .ZN(n9498) );
  AOI22D1BWP30P140LVT U13874 ( .A1(i_data_bus[155]), .A2(n9522), .B1(
        i_data_bus[219]), .B2(n9521), .ZN(n9497) );
  ND2D1BWP30P140LVT U13875 ( .A1(n9498), .A2(n9497), .ZN(N5156) );
  AOI22D1BWP30P140LVT U13876 ( .A1(i_data_bus[295]), .A2(n10276), .B1(
        i_data_bus[359]), .B2(n10277), .ZN(n9500) );
  AOI22D1BWP30P140LVT U13877 ( .A1(i_data_bus[263]), .A2(n6227), .B1(
        i_data_bus[327]), .B2(n10275), .ZN(n9499) );
  ND2D1BWP30P140LVT U13878 ( .A1(n9500), .A2(n9499), .ZN(N9182) );
  AOI22D1BWP30P140LVT U13879 ( .A1(i_data_bus[176]), .A2(n9519), .B1(
        i_data_bus[240]), .B2(n9520), .ZN(n9502) );
  AOI22D1BWP30P140LVT U13880 ( .A1(i_data_bus[144]), .A2(n9522), .B1(
        i_data_bus[208]), .B2(n9521), .ZN(n9501) );
  ND2D1BWP30P140LVT U13881 ( .A1(n9502), .A2(n9501), .ZN(N5145) );
  AOI22D1BWP30P140LVT U13882 ( .A1(i_data_bus[174]), .A2(n9519), .B1(
        i_data_bus[238]), .B2(n9520), .ZN(n9504) );
  AOI22D1BWP30P140LVT U13883 ( .A1(i_data_bus[142]), .A2(n9522), .B1(
        i_data_bus[206]), .B2(n9521), .ZN(n9503) );
  ND2D1BWP30P140LVT U13884 ( .A1(n9504), .A2(n9503), .ZN(N5143) );
  AOI22D1BWP30P140LVT U13885 ( .A1(i_data_bus[140]), .A2(n9522), .B1(
        i_data_bus[172]), .B2(n9519), .ZN(n9506) );
  AOI22D1BWP30P140LVT U13886 ( .A1(i_data_bus[236]), .A2(n9520), .B1(
        i_data_bus[204]), .B2(n9521), .ZN(n9505) );
  ND2D1BWP30P140LVT U13887 ( .A1(n9506), .A2(n9505), .ZN(N5141) );
  AOI22D1BWP30P140LVT U13888 ( .A1(i_data_bus[166]), .A2(n9519), .B1(
        i_data_bus[134]), .B2(n9522), .ZN(n9508) );
  AOI22D1BWP30P140LVT U13889 ( .A1(i_data_bus[230]), .A2(n9520), .B1(
        i_data_bus[198]), .B2(n9521), .ZN(n9507) );
  ND2D1BWP30P140LVT U13890 ( .A1(n9508), .A2(n9507), .ZN(N5135) );
  AOI22D1BWP30P140LVT U13891 ( .A1(i_data_bus[13]), .A2(n9969), .B1(
        i_data_bus[109]), .B2(n9978), .ZN(n9510) );
  AOI22D1BWP30P140LVT U13892 ( .A1(i_data_bus[45]), .A2(n9977), .B1(
        i_data_bus[77]), .B2(n9976), .ZN(n9509) );
  ND2D1BWP30P140LVT U13893 ( .A1(n9510), .A2(n9509), .ZN(N2330) );
  AOI22D1BWP30P140LVT U13894 ( .A1(i_data_bus[52]), .A2(n10118), .B1(
        i_data_bus[116]), .B2(n10117), .ZN(n9512) );
  AOI22D1BWP30P140LVT U13895 ( .A1(i_data_bus[20]), .A2(n10116), .B1(
        i_data_bus[84]), .B2(n10115), .ZN(n9511) );
  ND2D1BWP30P140LVT U13896 ( .A1(n9512), .A2(n9511), .ZN(N7785) );
  AOI22D1BWP30P140LVT U13897 ( .A1(i_data_bus[21]), .A2(n10116), .B1(
        i_data_bus[117]), .B2(n10117), .ZN(n9514) );
  AOI22D1BWP30P140LVT U13898 ( .A1(i_data_bus[53]), .A2(n10118), .B1(
        i_data_bus[85]), .B2(n10115), .ZN(n9513) );
  ND2D1BWP30P140LVT U13899 ( .A1(n9514), .A2(n9513), .ZN(N7786) );
  AOI22D1BWP30P140LVT U13900 ( .A1(i_data_bus[234]), .A2(n9520), .B1(
        i_data_bus[170]), .B2(n9519), .ZN(n9516) );
  AOI22D1BWP30P140LVT U13901 ( .A1(i_data_bus[138]), .A2(n9522), .B1(
        i_data_bus[202]), .B2(n9521), .ZN(n9515) );
  ND2D1BWP30P140LVT U13902 ( .A1(n9516), .A2(n9515), .ZN(N5139) );
  AOI22D1BWP30P140LVT U13903 ( .A1(i_data_bus[25]), .A2(n9969), .B1(
        i_data_bus[57]), .B2(n9977), .ZN(n9518) );
  AOI22D1BWP30P140LVT U13904 ( .A1(i_data_bus[121]), .A2(n9978), .B1(
        i_data_bus[89]), .B2(n9976), .ZN(n9517) );
  ND2D1BWP30P140LVT U13905 ( .A1(n9518), .A2(n9517), .ZN(N2342) );
  AOI22D1BWP30P140LVT U13906 ( .A1(i_data_bus[227]), .A2(n9520), .B1(
        i_data_bus[163]), .B2(n9519), .ZN(n9524) );
  AOI22D1BWP30P140LVT U13907 ( .A1(i_data_bus[131]), .A2(n9522), .B1(
        i_data_bus[195]), .B2(n9521), .ZN(n9523) );
  ND2D1BWP30P140LVT U13908 ( .A1(n9524), .A2(n9523), .ZN(N5132) );
  AOI22D1BWP30P140LVT U13909 ( .A1(i_data_bus[304]), .A2(n10276), .B1(
        i_data_bus[368]), .B2(n10277), .ZN(n9526) );
  AOI22D1BWP30P140LVT U13910 ( .A1(i_data_bus[272]), .A2(n6227), .B1(
        i_data_bus[336]), .B2(n10275), .ZN(n9525) );
  ND2D1BWP30P140LVT U13911 ( .A1(n9526), .A2(n9525), .ZN(N9191) );
  AOI22D1BWP30P140LVT U13912 ( .A1(i_data_bus[896]), .A2(n6226), .B1(
        i_data_bus[992]), .B2(n9543), .ZN(n9528) );
  AOI22D1BWP30P140LVT U13913 ( .A1(i_data_bus[928]), .A2(n9545), .B1(
        i_data_bus[960]), .B2(n9544), .ZN(n9527) );
  ND2D1BWP30P140LVT U13914 ( .A1(n9528), .A2(n9527), .ZN(N2083) );
  AOI22D1BWP30P140LVT U13915 ( .A1(i_data_bus[940]), .A2(n9545), .B1(
        i_data_bus[1004]), .B2(n9543), .ZN(n9530) );
  AOI22D1BWP30P140LVT U13916 ( .A1(i_data_bus[908]), .A2(n6226), .B1(
        i_data_bus[972]), .B2(n9544), .ZN(n9529) );
  ND2D1BWP30P140LVT U13917 ( .A1(n9530), .A2(n9529), .ZN(N2095) );
  AOI22D1BWP30P140LVT U13918 ( .A1(i_data_bus[958]), .A2(n9545), .B1(
        i_data_bus[926]), .B2(n6226), .ZN(n9532) );
  AOI22D1BWP30P140LVT U13919 ( .A1(i_data_bus[1022]), .A2(n9543), .B1(
        i_data_bus[990]), .B2(n9544), .ZN(n9531) );
  ND2D1BWP30P140LVT U13920 ( .A1(n9532), .A2(n9531), .ZN(N2113) );
  AOI22D1BWP30P140LVT U13921 ( .A1(i_data_bus[957]), .A2(n9545), .B1(
        i_data_bus[925]), .B2(n6226), .ZN(n9534) );
  AOI22D1BWP30P140LVT U13922 ( .A1(i_data_bus[1021]), .A2(n9543), .B1(
        i_data_bus[989]), .B2(n9544), .ZN(n9533) );
  ND2D1BWP30P140LVT U13923 ( .A1(n9534), .A2(n9533), .ZN(N2112) );
  AOI22D1BWP30P140LVT U13924 ( .A1(i_data_bus[954]), .A2(n9545), .B1(
        i_data_bus[1018]), .B2(n9543), .ZN(n9536) );
  AOI22D1BWP30P140LVT U13925 ( .A1(i_data_bus[922]), .A2(n6226), .B1(
        i_data_bus[986]), .B2(n9544), .ZN(n9535) );
  ND2D1BWP30P140LVT U13926 ( .A1(n9536), .A2(n9535), .ZN(N2109) );
  AOI22D1BWP30P140LVT U13927 ( .A1(i_data_bus[1012]), .A2(n9543), .B1(
        i_data_bus[916]), .B2(n6226), .ZN(n9538) );
  AOI22D1BWP30P140LVT U13928 ( .A1(i_data_bus[948]), .A2(n9545), .B1(
        i_data_bus[980]), .B2(n9544), .ZN(n9537) );
  ND2D1BWP30P140LVT U13929 ( .A1(n9538), .A2(n9537), .ZN(N2103) );
  AOI22D1BWP30P140LVT U13930 ( .A1(i_data_bus[914]), .A2(n6226), .B1(
        i_data_bus[946]), .B2(n9545), .ZN(n9540) );
  AOI22D1BWP30P140LVT U13931 ( .A1(i_data_bus[1010]), .A2(n9543), .B1(
        i_data_bus[978]), .B2(n9544), .ZN(n9539) );
  ND2D1BWP30P140LVT U13932 ( .A1(n9540), .A2(n9539), .ZN(N2101) );
  AOI22D1BWP30P140LVT U13933 ( .A1(i_data_bus[1005]), .A2(n9543), .B1(
        i_data_bus[941]), .B2(n9545), .ZN(n9542) );
  AOI22D1BWP30P140LVT U13934 ( .A1(i_data_bus[909]), .A2(n6226), .B1(
        i_data_bus[973]), .B2(n9544), .ZN(n9541) );
  ND2D1BWP30P140LVT U13935 ( .A1(n9542), .A2(n9541), .ZN(N2096) );
  AOI22D1BWP30P140LVT U13936 ( .A1(i_data_bus[906]), .A2(n6226), .B1(
        i_data_bus[1002]), .B2(n9543), .ZN(n9547) );
  AOI22D1BWP30P140LVT U13937 ( .A1(i_data_bus[938]), .A2(n9545), .B1(
        i_data_bus[970]), .B2(n9544), .ZN(n9546) );
  ND2D1BWP30P140LVT U13938 ( .A1(n9547), .A2(n9546), .ZN(N2093) );
  AOI22D1BWP30P140LVT U13939 ( .A1(i_data_bus[355]), .A2(n9877), .B1(
        i_data_bus[291]), .B2(n9878), .ZN(n9549) );
  AOI22D1BWP30P140LVT U13940 ( .A1(i_data_bus[259]), .A2(n6217), .B1(
        i_data_bus[323]), .B2(n9879), .ZN(n9548) );
  ND2D1BWP30P140LVT U13941 ( .A1(n9549), .A2(n9548), .ZN(N10668) );
  AOI22D1BWP30P140LVT U13942 ( .A1(i_data_bus[262]), .A2(n6217), .B1(
        i_data_bus[294]), .B2(n9878), .ZN(n9551) );
  AOI22D1BWP30P140LVT U13943 ( .A1(i_data_bus[358]), .A2(n9877), .B1(
        i_data_bus[326]), .B2(n9879), .ZN(n9550) );
  ND2D1BWP30P140LVT U13944 ( .A1(n9551), .A2(n9550), .ZN(N10671) );
  AOI22D1BWP30P140LVT U13945 ( .A1(i_data_bus[318]), .A2(n9843), .B1(
        i_data_bus[382]), .B2(n9845), .ZN(n9553) );
  AOI22D1BWP30P140LVT U13946 ( .A1(i_data_bus[286]), .A2(n9846), .B1(
        i_data_bus[350]), .B2(n9844), .ZN(n9552) );
  ND2D1BWP30P140LVT U13947 ( .A1(n9553), .A2(n9552), .ZN(N7971) );
  AOI22D1BWP30P140LVT U13948 ( .A1(i_data_bus[263]), .A2(n9846), .B1(
        i_data_bus[359]), .B2(n9845), .ZN(n9555) );
  AOI22D1BWP30P140LVT U13949 ( .A1(i_data_bus[295]), .A2(n9843), .B1(
        i_data_bus[327]), .B2(n9844), .ZN(n9554) );
  ND2D1BWP30P140LVT U13950 ( .A1(n9555), .A2(n9554), .ZN(N7948) );
  AOI22D1BWP30P140LVT U13951 ( .A1(i_data_bus[365]), .A2(n10051), .B1(
        i_data_bus[269]), .B2(n10052), .ZN(n9557) );
  AOI22D1BWP30P140LVT U13952 ( .A1(i_data_bus[301]), .A2(n10053), .B1(
        i_data_bus[333]), .B2(n10054), .ZN(n9556) );
  ND2D1BWP30P140LVT U13953 ( .A1(n9557), .A2(n9556), .ZN(N6464) );
  AOI22D1BWP30P140LVT U13954 ( .A1(i_data_bus[266]), .A2(n10052), .B1(
        i_data_bus[362]), .B2(n10051), .ZN(n9559) );
  AOI22D1BWP30P140LVT U13955 ( .A1(i_data_bus[298]), .A2(n10053), .B1(
        i_data_bus[330]), .B2(n10054), .ZN(n9558) );
  ND2D1BWP30P140LVT U13956 ( .A1(n9559), .A2(n9558), .ZN(N6461) );
  AOI22D1BWP30P140LVT U13957 ( .A1(i_data_bus[261]), .A2(n10052), .B1(
        i_data_bus[293]), .B2(n10053), .ZN(n9561) );
  AOI22D1BWP30P140LVT U13958 ( .A1(i_data_bus[357]), .A2(n10051), .B1(
        i_data_bus[325]), .B2(n10054), .ZN(n9560) );
  ND2D1BWP30P140LVT U13959 ( .A1(n9561), .A2(n9560), .ZN(N6456) );
  AOI22D1BWP30P140LVT U13960 ( .A1(i_data_bus[353]), .A2(n10051), .B1(
        i_data_bus[257]), .B2(n10052), .ZN(n9563) );
  AOI22D1BWP30P140LVT U13961 ( .A1(i_data_bus[289]), .A2(n10053), .B1(
        i_data_bus[321]), .B2(n10054), .ZN(n9562) );
  ND2D1BWP30P140LVT U13962 ( .A1(n9563), .A2(n9562), .ZN(N6452) );
  AOI22D1BWP30P140LVT U13963 ( .A1(i_data_bus[279]), .A2(n9846), .B1(
        i_data_bus[311]), .B2(n9843), .ZN(n9565) );
  AOI22D1BWP30P140LVT U13964 ( .A1(i_data_bus[375]), .A2(n9845), .B1(
        i_data_bus[343]), .B2(n9844), .ZN(n9564) );
  ND2D1BWP30P140LVT U13965 ( .A1(n9565), .A2(n9564), .ZN(N7964) );
  AOI22D1BWP30P140LVT U13966 ( .A1(i_data_bus[309]), .A2(n9843), .B1(
        i_data_bus[373]), .B2(n9845), .ZN(n9567) );
  AOI22D1BWP30P140LVT U13967 ( .A1(i_data_bus[277]), .A2(n9846), .B1(
        i_data_bus[341]), .B2(n9844), .ZN(n9566) );
  ND2D1BWP30P140LVT U13968 ( .A1(n9567), .A2(n9566), .ZN(N7962) );
  AOI22D1BWP30P140LVT U13969 ( .A1(i_data_bus[365]), .A2(n9845), .B1(
        i_data_bus[269]), .B2(n9846), .ZN(n9569) );
  AOI22D1BWP30P140LVT U13970 ( .A1(i_data_bus[301]), .A2(n9843), .B1(
        i_data_bus[333]), .B2(n9844), .ZN(n9568) );
  ND2D1BWP30P140LVT U13971 ( .A1(n9569), .A2(n9568), .ZN(N7954) );
  AOI22D1BWP30P140LVT U13972 ( .A1(i_data_bus[361]), .A2(n9845), .B1(
        i_data_bus[265]), .B2(n9846), .ZN(n9571) );
  AOI22D1BWP30P140LVT U13973 ( .A1(i_data_bus[297]), .A2(n9843), .B1(
        i_data_bus[329]), .B2(n9844), .ZN(n9570) );
  ND2D1BWP30P140LVT U13974 ( .A1(n9571), .A2(n9570), .ZN(N7950) );
  AOI22D1BWP30P140LVT U13975 ( .A1(i_data_bus[357]), .A2(n9845), .B1(
        i_data_bus[293]), .B2(n9843), .ZN(n9573) );
  AOI22D1BWP30P140LVT U13976 ( .A1(i_data_bus[261]), .A2(n9846), .B1(
        i_data_bus[325]), .B2(n9844), .ZN(n9572) );
  ND2D1BWP30P140LVT U13977 ( .A1(n9573), .A2(n9572), .ZN(N7946) );
  AOI22D1BWP30P140LVT U13978 ( .A1(i_data_bus[310]), .A2(n9878), .B1(
        i_data_bus[374]), .B2(n9877), .ZN(n9575) );
  AOI22D1BWP30P140LVT U13979 ( .A1(i_data_bus[278]), .A2(n6217), .B1(
        i_data_bus[342]), .B2(n9879), .ZN(n9574) );
  ND2D1BWP30P140LVT U13980 ( .A1(n9575), .A2(n9574), .ZN(N10687) );
  AOI22D1BWP30P140LVT U13981 ( .A1(i_data_bus[309]), .A2(n9878), .B1(
        i_data_bus[277]), .B2(n6217), .ZN(n9577) );
  AOI22D1BWP30P140LVT U13982 ( .A1(i_data_bus[373]), .A2(n9877), .B1(
        i_data_bus[341]), .B2(n9879), .ZN(n9576) );
  ND2D1BWP30P140LVT U13983 ( .A1(n9577), .A2(n9576), .ZN(N10686) );
  AOI22D1BWP30P140LVT U13984 ( .A1(i_data_bus[272]), .A2(n6217), .B1(
        i_data_bus[304]), .B2(n9878), .ZN(n9579) );
  AOI22D1BWP30P140LVT U13985 ( .A1(i_data_bus[368]), .A2(n9877), .B1(
        i_data_bus[336]), .B2(n9879), .ZN(n9578) );
  ND2D1BWP30P140LVT U13986 ( .A1(n9579), .A2(n9578), .ZN(N10681) );
  AOI22D1BWP30P140LVT U13987 ( .A1(i_data_bus[271]), .A2(n10052), .B1(
        i_data_bus[367]), .B2(n10051), .ZN(n9581) );
  AOI22D1BWP30P140LVT U13988 ( .A1(i_data_bus[303]), .A2(n10053), .B1(
        i_data_bus[335]), .B2(n10054), .ZN(n9580) );
  ND2D1BWP30P140LVT U13989 ( .A1(n9581), .A2(n9580), .ZN(N6466) );
  AOI22D1BWP30P140LVT U13990 ( .A1(i_data_bus[284]), .A2(n10052), .B1(
        i_data_bus[316]), .B2(n10053), .ZN(n9583) );
  AOI22D1BWP30P140LVT U13991 ( .A1(i_data_bus[380]), .A2(n10051), .B1(
        i_data_bus[348]), .B2(n10054), .ZN(n9582) );
  ND2D1BWP30P140LVT U13992 ( .A1(n9583), .A2(n9582), .ZN(N6479) );
  AOI22D1BWP30P140LVT U13993 ( .A1(i_data_bus[268]), .A2(n9846), .B1(
        i_data_bus[300]), .B2(n9843), .ZN(n9585) );
  AOI22D1BWP30P140LVT U13994 ( .A1(i_data_bus[364]), .A2(n9845), .B1(
        i_data_bus[332]), .B2(n9844), .ZN(n9584) );
  ND2D1BWP30P140LVT U13995 ( .A1(n9585), .A2(n9584), .ZN(N7953) );
  AOI22D1BWP30P140LVT U13996 ( .A1(i_data_bus[313]), .A2(n9878), .B1(
        i_data_bus[377]), .B2(n9877), .ZN(n9587) );
  AOI22D1BWP30P140LVT U13997 ( .A1(i_data_bus[281]), .A2(n6217), .B1(
        i_data_bus[345]), .B2(n9879), .ZN(n9586) );
  ND2D1BWP30P140LVT U13998 ( .A1(n9587), .A2(n9586), .ZN(N10690) );
  AOI22D1BWP30P140LVT U13999 ( .A1(i_data_bus[376]), .A2(n10051), .B1(
        i_data_bus[312]), .B2(n10053), .ZN(n9589) );
  AOI22D1BWP30P140LVT U14000 ( .A1(i_data_bus[280]), .A2(n10052), .B1(
        i_data_bus[344]), .B2(n10054), .ZN(n9588) );
  ND2D1BWP30P140LVT U14001 ( .A1(n9589), .A2(n9588), .ZN(N6475) );
  AOI22D1BWP30P140LVT U14002 ( .A1(i_data_bus[260]), .A2(n6217), .B1(
        i_data_bus[292]), .B2(n9878), .ZN(n9591) );
  AOI22D1BWP30P140LVT U14003 ( .A1(i_data_bus[356]), .A2(n9877), .B1(
        i_data_bus[324]), .B2(n9879), .ZN(n9590) );
  ND2D1BWP30P140LVT U14004 ( .A1(n9591), .A2(n9590), .ZN(N10669) );
  AOI22D1BWP30P140LVT U14005 ( .A1(i_data_bus[313]), .A2(n10053), .B1(
        i_data_bus[377]), .B2(n10051), .ZN(n9593) );
  AOI22D1BWP30P140LVT U14006 ( .A1(i_data_bus[281]), .A2(n10052), .B1(
        i_data_bus[345]), .B2(n10054), .ZN(n9592) );
  ND2D1BWP30P140LVT U14007 ( .A1(n9593), .A2(n9592), .ZN(N6476) );
  AOI22D1BWP30P140LVT U14008 ( .A1(i_data_bus[316]), .A2(n9732), .B1(
        i_data_bus[380]), .B2(n9730), .ZN(n9595) );
  AOI22D1BWP30P140LVT U14009 ( .A1(i_data_bus[284]), .A2(n6219), .B1(
        i_data_bus[348]), .B2(n9731), .ZN(n9594) );
  ND2D1BWP30P140LVT U14010 ( .A1(n9595), .A2(n9594), .ZN(N3755) );
  AOI22D1BWP30P140LVT U14011 ( .A1(i_data_bus[315]), .A2(n9732), .B1(
        i_data_bus[379]), .B2(n9730), .ZN(n9597) );
  AOI22D1BWP30P140LVT U14012 ( .A1(i_data_bus[283]), .A2(n6219), .B1(
        i_data_bus[347]), .B2(n9731), .ZN(n9596) );
  ND2D1BWP30P140LVT U14013 ( .A1(n9597), .A2(n9596), .ZN(N3754) );
  AOI22D1BWP30P140LVT U14014 ( .A1(i_data_bus[313]), .A2(n9732), .B1(
        i_data_bus[377]), .B2(n9730), .ZN(n9599) );
  AOI22D1BWP30P140LVT U14015 ( .A1(i_data_bus[281]), .A2(n6219), .B1(
        i_data_bus[345]), .B2(n9731), .ZN(n9598) );
  ND2D1BWP30P140LVT U14016 ( .A1(n9599), .A2(n9598), .ZN(N3752) );
  AOI22D1BWP30P140LVT U14017 ( .A1(i_data_bus[271]), .A2(n6219), .B1(
        i_data_bus[367]), .B2(n9730), .ZN(n9601) );
  AOI22D1BWP30P140LVT U14018 ( .A1(i_data_bus[303]), .A2(n9732), .B1(
        i_data_bus[335]), .B2(n9731), .ZN(n9600) );
  ND2D1BWP30P140LVT U14019 ( .A1(n9601), .A2(n9600), .ZN(N3742) );
  AOI22D1BWP30P140LVT U14020 ( .A1(i_data_bus[301]), .A2(n9732), .B1(
        i_data_bus[269]), .B2(n6219), .ZN(n9603) );
  AOI22D1BWP30P140LVT U14021 ( .A1(i_data_bus[365]), .A2(n9730), .B1(
        i_data_bus[333]), .B2(n9731), .ZN(n9602) );
  ND2D1BWP30P140LVT U14022 ( .A1(n9603), .A2(n9602), .ZN(N3740) );
  AOI22D1BWP30P140LVT U14023 ( .A1(i_data_bus[363]), .A2(n9730), .B1(
        i_data_bus[267]), .B2(n6219), .ZN(n9605) );
  AOI22D1BWP30P140LVT U14024 ( .A1(i_data_bus[299]), .A2(n9732), .B1(
        i_data_bus[331]), .B2(n9731), .ZN(n9604) );
  ND2D1BWP30P140LVT U14025 ( .A1(n9605), .A2(n9604), .ZN(N3738) );
  AOI22D1BWP30P140LVT U14026 ( .A1(i_data_bus[261]), .A2(n6219), .B1(
        i_data_bus[293]), .B2(n9732), .ZN(n9607) );
  AOI22D1BWP30P140LVT U14027 ( .A1(i_data_bus[357]), .A2(n9730), .B1(
        i_data_bus[325]), .B2(n9731), .ZN(n9606) );
  ND2D1BWP30P140LVT U14028 ( .A1(n9607), .A2(n9606), .ZN(N3732) );
  AOI22D1BWP30P140LVT U14029 ( .A1(i_data_bus[62]), .A2(n9916), .B1(
        i_data_bus[126]), .B2(n9915), .ZN(n9609) );
  AOI22D1BWP30P140LVT U14030 ( .A1(i_data_bus[30]), .A2(n6218), .B1(
        i_data_bus[94]), .B2(n9914), .ZN(n9608) );
  ND2D1BWP30P140LVT U14031 ( .A1(n9609), .A2(n9608), .ZN(N3325) );
  AOI22D1BWP30P140LVT U14032 ( .A1(i_data_bus[121]), .A2(n9915), .B1(
        i_data_bus[57]), .B2(n9916), .ZN(n9611) );
  AOI22D1BWP30P140LVT U14033 ( .A1(i_data_bus[25]), .A2(n6218), .B1(
        i_data_bus[89]), .B2(n9914), .ZN(n9610) );
  ND2D1BWP30P140LVT U14034 ( .A1(n9611), .A2(n9610), .ZN(N3320) );
  AOI22D1BWP30P140LVT U14035 ( .A1(i_data_bus[45]), .A2(n9916), .B1(
        i_data_bus[109]), .B2(n9915), .ZN(n9613) );
  AOI22D1BWP30P140LVT U14036 ( .A1(i_data_bus[13]), .A2(n6218), .B1(
        i_data_bus[77]), .B2(n9914), .ZN(n9612) );
  ND2D1BWP30P140LVT U14037 ( .A1(n9613), .A2(n9612), .ZN(N3308) );
  AOI22D1BWP30P140LVT U14038 ( .A1(i_data_bus[1]), .A2(n6218), .B1(
        i_data_bus[97]), .B2(n9915), .ZN(n9615) );
  AOI22D1BWP30P140LVT U14039 ( .A1(i_data_bus[33]), .A2(n9916), .B1(
        i_data_bus[65]), .B2(n9914), .ZN(n9614) );
  ND2D1BWP30P140LVT U14040 ( .A1(n9615), .A2(n9614), .ZN(N3296) );
  AOI22D1BWP30P140LVT U14041 ( .A1(i_data_bus[148]), .A2(n10026), .B1(
        i_data_bus[180]), .B2(n10034), .ZN(n9617) );
  AOI22D1BWP30P140LVT U14042 ( .A1(i_data_bus[244]), .A2(n10035), .B1(
        i_data_bus[212]), .B2(n10033), .ZN(n9616) );
  ND2D1BWP30P140LVT U14043 ( .A1(n9617), .A2(n9616), .ZN(N3531) );
  AOI22D1BWP30P140LVT U14044 ( .A1(i_data_bus[242]), .A2(n10035), .B1(
        i_data_bus[178]), .B2(n10034), .ZN(n9619) );
  AOI22D1BWP30P140LVT U14045 ( .A1(i_data_bus[146]), .A2(n10026), .B1(
        i_data_bus[210]), .B2(n10033), .ZN(n9618) );
  ND2D1BWP30P140LVT U14046 ( .A1(n9619), .A2(n9618), .ZN(N3529) );
  AOI22D1BWP30P140LVT U14047 ( .A1(i_data_bus[144]), .A2(n10026), .B1(
        i_data_bus[176]), .B2(n10034), .ZN(n9621) );
  AOI22D1BWP30P140LVT U14048 ( .A1(i_data_bus[240]), .A2(n10035), .B1(
        i_data_bus[208]), .B2(n10033), .ZN(n9620) );
  ND2D1BWP30P140LVT U14049 ( .A1(n9621), .A2(n9620), .ZN(N3527) );
  AOI22D1BWP30P140LVT U14050 ( .A1(i_data_bus[140]), .A2(n10026), .B1(
        i_data_bus[236]), .B2(n10035), .ZN(n9623) );
  AOI22D1BWP30P140LVT U14051 ( .A1(i_data_bus[172]), .A2(n10034), .B1(
        i_data_bus[204]), .B2(n10033), .ZN(n9622) );
  ND2D1BWP30P140LVT U14052 ( .A1(n9623), .A2(n9622), .ZN(N3523) );
  AOI22D1BWP30P140LVT U14053 ( .A1(i_data_bus[234]), .A2(n10035), .B1(
        i_data_bus[170]), .B2(n10034), .ZN(n9625) );
  AOI22D1BWP30P140LVT U14054 ( .A1(i_data_bus[138]), .A2(n10026), .B1(
        i_data_bus[202]), .B2(n10033), .ZN(n9624) );
  ND2D1BWP30P140LVT U14055 ( .A1(n9625), .A2(n9624), .ZN(N3521) );
  AOI22D1BWP30P140LVT U14056 ( .A1(i_data_bus[135]), .A2(n10026), .B1(
        i_data_bus[167]), .B2(n10034), .ZN(n9627) );
  AOI22D1BWP30P140LVT U14057 ( .A1(i_data_bus[231]), .A2(n10035), .B1(
        i_data_bus[199]), .B2(n10033), .ZN(n9626) );
  ND2D1BWP30P140LVT U14058 ( .A1(n9627), .A2(n9626), .ZN(N3518) );
  AOI22D1BWP30P140LVT U14059 ( .A1(i_data_bus[166]), .A2(n10034), .B1(
        i_data_bus[134]), .B2(n10026), .ZN(n9629) );
  AOI22D1BWP30P140LVT U14060 ( .A1(i_data_bus[230]), .A2(n10035), .B1(
        i_data_bus[198]), .B2(n10033), .ZN(n9628) );
  ND2D1BWP30P140LVT U14061 ( .A1(n9629), .A2(n9628), .ZN(N3517) );
  AOI22D1BWP30P140LVT U14062 ( .A1(i_data_bus[188]), .A2(n10034), .B1(
        i_data_bus[252]), .B2(n10035), .ZN(n9631) );
  AOI22D1BWP30P140LVT U14063 ( .A1(i_data_bus[156]), .A2(n10026), .B1(
        i_data_bus[220]), .B2(n10033), .ZN(n9630) );
  ND2D1BWP30P140LVT U14064 ( .A1(n9631), .A2(n9630), .ZN(N3539) );
  AOI22D1BWP30P140LVT U14065 ( .A1(i_data_bus[137]), .A2(n10026), .B1(
        i_data_bus[233]), .B2(n10035), .ZN(n9633) );
  AOI22D1BWP30P140LVT U14066 ( .A1(i_data_bus[169]), .A2(n10034), .B1(
        i_data_bus[201]), .B2(n10033), .ZN(n9632) );
  ND2D1BWP30P140LVT U14067 ( .A1(n9633), .A2(n9632), .ZN(N3520) );
  AOI22D1BWP30P140LVT U14068 ( .A1(i_data_bus[117]), .A2(n9915), .B1(
        i_data_bus[53]), .B2(n9916), .ZN(n9635) );
  AOI22D1BWP30P140LVT U14069 ( .A1(i_data_bus[21]), .A2(n6218), .B1(
        i_data_bus[85]), .B2(n9914), .ZN(n9634) );
  ND2D1BWP30P140LVT U14070 ( .A1(n9635), .A2(n9634), .ZN(N3316) );
  AOI22D1BWP30P140LVT U14071 ( .A1(i_data_bus[113]), .A2(n9915), .B1(
        i_data_bus[49]), .B2(n9916), .ZN(n9637) );
  AOI22D1BWP30P140LVT U14072 ( .A1(i_data_bus[17]), .A2(n6218), .B1(
        i_data_bus[81]), .B2(n9914), .ZN(n9636) );
  ND2D1BWP30P140LVT U14073 ( .A1(n9637), .A2(n9636), .ZN(N3312) );
  AOI22D1BWP30P140LVT U14074 ( .A1(i_data_bus[27]), .A2(n6218), .B1(
        i_data_bus[59]), .B2(n9916), .ZN(n9639) );
  AOI22D1BWP30P140LVT U14075 ( .A1(i_data_bus[123]), .A2(n9915), .B1(
        i_data_bus[91]), .B2(n9914), .ZN(n9638) );
  ND2D1BWP30P140LVT U14076 ( .A1(n9639), .A2(n9638), .ZN(N3322) );
  AOI22D1BWP30P140LVT U14077 ( .A1(i_data_bus[5]), .A2(n6218), .B1(
        i_data_bus[37]), .B2(n9916), .ZN(n9641) );
  AOI22D1BWP30P140LVT U14078 ( .A1(i_data_bus[101]), .A2(n9915), .B1(
        i_data_bus[69]), .B2(n9914), .ZN(n9640) );
  ND2D1BWP30P140LVT U14079 ( .A1(n9641), .A2(n9640), .ZN(N3300) );
  AOI22D1BWP30P140LVT U14080 ( .A1(i_data_bus[1023]), .A2(n9663), .B1(
        i_data_bus[927]), .B2(n9661), .ZN(n9643) );
  AOI22D1BWP30P140LVT U14081 ( .A1(i_data_bus[959]), .A2(n9660), .B1(
        i_data_bus[991]), .B2(n9662), .ZN(n9642) );
  ND2D1BWP30P140LVT U14082 ( .A1(n9643), .A2(n9642), .ZN(N7562) );
  AOI22D1BWP30P140LVT U14083 ( .A1(i_data_bus[955]), .A2(n9660), .B1(
        i_data_bus[1019]), .B2(n9663), .ZN(n9645) );
  AOI22D1BWP30P140LVT U14084 ( .A1(i_data_bus[923]), .A2(n9661), .B1(
        i_data_bus[987]), .B2(n9662), .ZN(n9644) );
  ND2D1BWP30P140LVT U14085 ( .A1(n9645), .A2(n9644), .ZN(N7558) );
  AOI22D1BWP30P140LVT U14086 ( .A1(i_data_bus[951]), .A2(n9660), .B1(
        i_data_bus[1015]), .B2(n9663), .ZN(n9647) );
  AOI22D1BWP30P140LVT U14087 ( .A1(i_data_bus[919]), .A2(n9661), .B1(
        i_data_bus[983]), .B2(n9662), .ZN(n9646) );
  ND2D1BWP30P140LVT U14088 ( .A1(n9647), .A2(n9646), .ZN(N7554) );
  AOI22D1BWP30P140LVT U14089 ( .A1(i_data_bus[1014]), .A2(n9663), .B1(
        i_data_bus[950]), .B2(n9660), .ZN(n9649) );
  AOI22D1BWP30P140LVT U14090 ( .A1(i_data_bus[918]), .A2(n9661), .B1(
        i_data_bus[982]), .B2(n9662), .ZN(n9648) );
  ND2D1BWP30P140LVT U14091 ( .A1(n9649), .A2(n9648), .ZN(N7553) );
  AOI22D1BWP30P140LVT U14092 ( .A1(i_data_bus[914]), .A2(n9661), .B1(
        i_data_bus[946]), .B2(n9660), .ZN(n9651) );
  AOI22D1BWP30P140LVT U14093 ( .A1(i_data_bus[1010]), .A2(n9663), .B1(
        i_data_bus[978]), .B2(n9662), .ZN(n9650) );
  ND2D1BWP30P140LVT U14094 ( .A1(n9651), .A2(n9650), .ZN(N7549) );
  AOI22D1BWP30P140LVT U14095 ( .A1(i_data_bus[906]), .A2(n9661), .B1(
        i_data_bus[1002]), .B2(n9663), .ZN(n9653) );
  AOI22D1BWP30P140LVT U14096 ( .A1(i_data_bus[938]), .A2(n9660), .B1(
        i_data_bus[970]), .B2(n9662), .ZN(n9652) );
  ND2D1BWP30P140LVT U14097 ( .A1(n9653), .A2(n9652), .ZN(N7541) );
  AOI22D1BWP30P140LVT U14098 ( .A1(i_data_bus[902]), .A2(n9661), .B1(
        i_data_bus[998]), .B2(n9663), .ZN(n9655) );
  AOI22D1BWP30P140LVT U14099 ( .A1(i_data_bus[934]), .A2(n9660), .B1(
        i_data_bus[966]), .B2(n9662), .ZN(n9654) );
  ND2D1BWP30P140LVT U14100 ( .A1(n9655), .A2(n9654), .ZN(N7537) );
  AOI22D1BWP30P140LVT U14101 ( .A1(i_data_bus[996]), .A2(n9663), .B1(
        i_data_bus[900]), .B2(n9661), .ZN(n9657) );
  AOI22D1BWP30P140LVT U14102 ( .A1(i_data_bus[932]), .A2(n9660), .B1(
        i_data_bus[964]), .B2(n9662), .ZN(n9656) );
  ND2D1BWP30P140LVT U14103 ( .A1(n9657), .A2(n9656), .ZN(N7535) );
  AOI22D1BWP30P140LVT U14104 ( .A1(i_data_bus[901]), .A2(n9661), .B1(
        i_data_bus[997]), .B2(n9663), .ZN(n9659) );
  AOI22D1BWP30P140LVT U14105 ( .A1(i_data_bus[933]), .A2(n9660), .B1(
        i_data_bus[965]), .B2(n9662), .ZN(n9658) );
  ND2D1BWP30P140LVT U14106 ( .A1(n9659), .A2(n9658), .ZN(N7536) );
  AOI22D1BWP30P140LVT U14107 ( .A1(i_data_bus[910]), .A2(n9661), .B1(
        i_data_bus[942]), .B2(n9660), .ZN(n9665) );
  AOI22D1BWP30P140LVT U14108 ( .A1(i_data_bus[1006]), .A2(n9663), .B1(
        i_data_bus[974]), .B2(n9662), .ZN(n9664) );
  ND2D1BWP30P140LVT U14109 ( .A1(n9665), .A2(n9664), .ZN(N7545) );
  AOI22D1BWP30P140LVT U14110 ( .A1(i_data_bus[301]), .A2(n9758), .B1(
        i_data_bus[269]), .B2(n9756), .ZN(n9667) );
  AOI22D1BWP30P140LVT U14111 ( .A1(i_data_bus[365]), .A2(n9757), .B1(
        i_data_bus[333]), .B2(n9755), .ZN(n9666) );
  ND2D1BWP30P140LVT U14112 ( .A1(n9667), .A2(n9666), .ZN(N5230) );
  AOI22D1BWP30P140LVT U14113 ( .A1(i_data_bus[260]), .A2(n9756), .B1(
        i_data_bus[292]), .B2(n9758), .ZN(n9669) );
  AOI22D1BWP30P140LVT U14114 ( .A1(i_data_bus[356]), .A2(n9757), .B1(
        i_data_bus[324]), .B2(n9755), .ZN(n9668) );
  ND2D1BWP30P140LVT U14115 ( .A1(n9669), .A2(n9668), .ZN(N5221) );
  AOI22D1BWP30P140LVT U14116 ( .A1(i_data_bus[279]), .A2(n9756), .B1(
        i_data_bus[311]), .B2(n9758), .ZN(n9671) );
  AOI22D1BWP30P140LVT U14117 ( .A1(i_data_bus[375]), .A2(n9757), .B1(
        i_data_bus[343]), .B2(n9755), .ZN(n9670) );
  ND2D1BWP30P140LVT U14118 ( .A1(n9671), .A2(n9670), .ZN(N5240) );
  AOI22D1BWP30P140LVT U14119 ( .A1(i_data_bus[315]), .A2(n9758), .B1(
        i_data_bus[379]), .B2(n9757), .ZN(n9673) );
  AOI22D1BWP30P140LVT U14120 ( .A1(i_data_bus[283]), .A2(n9756), .B1(
        i_data_bus[347]), .B2(n9755), .ZN(n9672) );
  ND2D1BWP30P140LVT U14121 ( .A1(n9673), .A2(n9672), .ZN(N5244) );
  AOI22D1BWP30P140LVT U14122 ( .A1(i_data_bus[310]), .A2(n9758), .B1(
        i_data_bus[374]), .B2(n9757), .ZN(n9675) );
  AOI22D1BWP30P140LVT U14123 ( .A1(i_data_bus[278]), .A2(n9756), .B1(
        i_data_bus[342]), .B2(n9755), .ZN(n9674) );
  ND2D1BWP30P140LVT U14124 ( .A1(n9675), .A2(n9674), .ZN(N5239) );
  AOI22D1BWP30P140LVT U14125 ( .A1(i_data_bus[270]), .A2(n9756), .B1(
        i_data_bus[366]), .B2(n9757), .ZN(n9677) );
  AOI22D1BWP30P140LVT U14126 ( .A1(i_data_bus[302]), .A2(n9758), .B1(
        i_data_bus[334]), .B2(n9755), .ZN(n9676) );
  ND2D1BWP30P140LVT U14127 ( .A1(n9677), .A2(n9676), .ZN(N5231) );
  AOI22D1BWP30P140LVT U14128 ( .A1(i_data_bus[361]), .A2(n9757), .B1(
        i_data_bus[265]), .B2(n9756), .ZN(n9679) );
  AOI22D1BWP30P140LVT U14129 ( .A1(i_data_bus[297]), .A2(n9758), .B1(
        i_data_bus[329]), .B2(n9755), .ZN(n9678) );
  ND2D1BWP30P140LVT U14130 ( .A1(n9679), .A2(n9678), .ZN(N5226) );
  AOI22D1BWP30P140LVT U14131 ( .A1(i_data_bus[264]), .A2(n9756), .B1(
        i_data_bus[296]), .B2(n9758), .ZN(n9681) );
  AOI22D1BWP30P140LVT U14132 ( .A1(i_data_bus[360]), .A2(n9757), .B1(
        i_data_bus[328]), .B2(n9755), .ZN(n9680) );
  ND2D1BWP30P140LVT U14133 ( .A1(n9681), .A2(n9680), .ZN(N5225) );
  AOI22D1BWP30P140LVT U14134 ( .A1(i_data_bus[357]), .A2(n9757), .B1(
        i_data_bus[293]), .B2(n9758), .ZN(n9683) );
  AOI22D1BWP30P140LVT U14135 ( .A1(i_data_bus[261]), .A2(n9756), .B1(
        i_data_bus[325]), .B2(n9755), .ZN(n9682) );
  ND2D1BWP30P140LVT U14136 ( .A1(n9683), .A2(n9682), .ZN(N5222) );
  AOI22D1BWP30P140LVT U14137 ( .A1(i_data_bus[363]), .A2(n9757), .B1(
        i_data_bus[267]), .B2(n9756), .ZN(n9685) );
  AOI22D1BWP30P140LVT U14138 ( .A1(i_data_bus[299]), .A2(n9758), .B1(
        i_data_bus[331]), .B2(n9755), .ZN(n9684) );
  ND2D1BWP30P140LVT U14139 ( .A1(n9685), .A2(n9684), .ZN(N5228) );
  AOI22D1BWP30P140LVT U14140 ( .A1(i_data_bus[8]), .A2(n6223), .B1(
        i_data_bus[40]), .B2(n9791), .ZN(n9687) );
  AOI22D1BWP30P140LVT U14141 ( .A1(i_data_bus[104]), .A2(n9792), .B1(
        i_data_bus[72]), .B2(n9790), .ZN(n9686) );
  ND2D1BWP30P140LVT U14142 ( .A1(n9687), .A2(n9686), .ZN(N8751) );
  AOI22D1BWP30P140LVT U14143 ( .A1(i_data_bus[56]), .A2(n9791), .B1(
        i_data_bus[120]), .B2(n9792), .ZN(n9689) );
  AOI22D1BWP30P140LVT U14144 ( .A1(i_data_bus[24]), .A2(n6223), .B1(
        i_data_bus[88]), .B2(n9790), .ZN(n9688) );
  ND2D1BWP30P140LVT U14145 ( .A1(n9689), .A2(n9688), .ZN(N8767) );
  AOI22D1BWP30P140LVT U14146 ( .A1(i_data_bus[103]), .A2(n9792), .B1(
        i_data_bus[39]), .B2(n9791), .ZN(n9691) );
  AOI22D1BWP30P140LVT U14147 ( .A1(i_data_bus[7]), .A2(n6223), .B1(
        i_data_bus[71]), .B2(n9790), .ZN(n9690) );
  ND2D1BWP30P140LVT U14148 ( .A1(n9691), .A2(n9690), .ZN(N8750) );
  AOI22D1BWP30P140LVT U14149 ( .A1(i_data_bus[26]), .A2(n6223), .B1(
        i_data_bus[58]), .B2(n9791), .ZN(n9693) );
  AOI22D1BWP30P140LVT U14150 ( .A1(i_data_bus[122]), .A2(n9792), .B1(
        i_data_bus[90]), .B2(n9790), .ZN(n9692) );
  ND2D1BWP30P140LVT U14151 ( .A1(n9693), .A2(n9692), .ZN(N8769) );
  AOI22D1BWP30P140LVT U14152 ( .A1(i_data_bus[25]), .A2(n6223), .B1(
        i_data_bus[57]), .B2(n9791), .ZN(n9695) );
  AOI22D1BWP30P140LVT U14153 ( .A1(i_data_bus[121]), .A2(n9792), .B1(
        i_data_bus[89]), .B2(n9790), .ZN(n9694) );
  ND2D1BWP30P140LVT U14154 ( .A1(n9695), .A2(n9694), .ZN(N8768) );
  AOI22D1BWP30P140LVT U14155 ( .A1(i_data_bus[36]), .A2(n9791), .B1(
        i_data_bus[4]), .B2(n6223), .ZN(n9697) );
  AOI22D1BWP30P140LVT U14156 ( .A1(i_data_bus[100]), .A2(n9792), .B1(
        i_data_bus[68]), .B2(n9790), .ZN(n9696) );
  ND2D1BWP30P140LVT U14157 ( .A1(n9697), .A2(n9696), .ZN(N8747) );
  AOI22D1BWP30P140LVT U14158 ( .A1(i_data_bus[0]), .A2(n6223), .B1(
        i_data_bus[96]), .B2(n9792), .ZN(n9699) );
  AOI22D1BWP30P140LVT U14159 ( .A1(i_data_bus[32]), .A2(n9791), .B1(
        i_data_bus[64]), .B2(n9790), .ZN(n9698) );
  ND2D1BWP30P140LVT U14160 ( .A1(n9699), .A2(n9698), .ZN(N8743) );
  AOI22D1BWP30P140LVT U14161 ( .A1(i_data_bus[30]), .A2(n6223), .B1(
        i_data_bus[62]), .B2(n9791), .ZN(n9701) );
  AOI22D1BWP30P140LVT U14162 ( .A1(i_data_bus[126]), .A2(n9792), .B1(
        i_data_bus[94]), .B2(n9790), .ZN(n9700) );
  ND2D1BWP30P140LVT U14163 ( .A1(n9701), .A2(n9700), .ZN(N8773) );
  AOI22D1BWP30P140LVT U14164 ( .A1(i_data_bus[28]), .A2(n6223), .B1(
        i_data_bus[124]), .B2(n9792), .ZN(n9703) );
  AOI22D1BWP30P140LVT U14165 ( .A1(i_data_bus[60]), .A2(n9791), .B1(
        i_data_bus[92]), .B2(n9790), .ZN(n9702) );
  ND2D1BWP30P140LVT U14166 ( .A1(n9703), .A2(n9702), .ZN(N8771) );
  AOI22D1BWP30P140LVT U14167 ( .A1(i_data_bus[51]), .A2(n9791), .B1(
        i_data_bus[115]), .B2(n9792), .ZN(n9705) );
  AOI22D1BWP30P140LVT U14168 ( .A1(i_data_bus[19]), .A2(n6223), .B1(
        i_data_bus[83]), .B2(n9790), .ZN(n9704) );
  ND2D1BWP30P140LVT U14169 ( .A1(n9705), .A2(n9704), .ZN(N8762) );
  AOI22D1BWP30P140LVT U14170 ( .A1(i_data_bus[97]), .A2(n9792), .B1(
        i_data_bus[33]), .B2(n9791), .ZN(n9707) );
  AOI22D1BWP30P140LVT U14171 ( .A1(i_data_bus[1]), .A2(n6223), .B1(
        i_data_bus[65]), .B2(n9790), .ZN(n9706) );
  ND2D1BWP30P140LVT U14172 ( .A1(n9707), .A2(n9706), .ZN(N8744) );
  AOI22D1BWP30P140LVT U14173 ( .A1(i_data_bus[16]), .A2(n6223), .B1(
        i_data_bus[112]), .B2(n9792), .ZN(n9709) );
  AOI22D1BWP30P140LVT U14174 ( .A1(i_data_bus[48]), .A2(n9791), .B1(
        i_data_bus[80]), .B2(n9790), .ZN(n9708) );
  ND2D1BWP30P140LVT U14175 ( .A1(n9709), .A2(n9708), .ZN(N8759) );
  AOI22D1BWP30P140LVT U14176 ( .A1(i_data_bus[27]), .A2(n6223), .B1(
        i_data_bus[59]), .B2(n9791), .ZN(n9711) );
  AOI22D1BWP30P140LVT U14177 ( .A1(i_data_bus[123]), .A2(n9792), .B1(
        i_data_bus[91]), .B2(n9790), .ZN(n9710) );
  ND2D1BWP30P140LVT U14178 ( .A1(n9711), .A2(n9710), .ZN(N8770) );
  AOI22D1BWP30P140LVT U14179 ( .A1(i_data_bus[113]), .A2(n9792), .B1(
        i_data_bus[49]), .B2(n9791), .ZN(n9713) );
  AOI22D1BWP30P140LVT U14180 ( .A1(i_data_bus[17]), .A2(n6223), .B1(
        i_data_bus[81]), .B2(n9790), .ZN(n9712) );
  ND2D1BWP30P140LVT U14181 ( .A1(n9713), .A2(n9712), .ZN(N8760) );
  AOI22D1BWP30P140LVT U14182 ( .A1(i_data_bus[346]), .A2(n9731), .B1(
        i_data_bus[378]), .B2(n9730), .ZN(n9715) );
  AOI22D1BWP30P140LVT U14183 ( .A1(i_data_bus[282]), .A2(n6219), .B1(
        i_data_bus[314]), .B2(n9732), .ZN(n9714) );
  ND2D1BWP30P140LVT U14184 ( .A1(n9715), .A2(n9714), .ZN(N3753) );
  AOI22D1BWP30P140LVT U14185 ( .A1(i_data_bus[338]), .A2(n9731), .B1(
        i_data_bus[370]), .B2(n9730), .ZN(n9717) );
  AOI22D1BWP30P140LVT U14186 ( .A1(i_data_bus[274]), .A2(n6219), .B1(
        i_data_bus[306]), .B2(n9732), .ZN(n9716) );
  ND2D1BWP30P140LVT U14187 ( .A1(n9717), .A2(n9716), .ZN(N3745) );
  AOI22D1BWP30P140LVT U14188 ( .A1(i_data_bus[337]), .A2(n9731), .B1(
        i_data_bus[369]), .B2(n9730), .ZN(n9719) );
  AOI22D1BWP30P140LVT U14189 ( .A1(i_data_bus[273]), .A2(n6219), .B1(
        i_data_bus[305]), .B2(n9732), .ZN(n9718) );
  ND2D1BWP30P140LVT U14190 ( .A1(n9719), .A2(n9718), .ZN(N3744) );
  AOI22D1BWP30P140LVT U14191 ( .A1(i_data_bus[268]), .A2(n6219), .B1(
        i_data_bus[332]), .B2(n9731), .ZN(n9721) );
  AOI22D1BWP30P140LVT U14192 ( .A1(i_data_bus[364]), .A2(n9730), .B1(
        i_data_bus[300]), .B2(n9732), .ZN(n9720) );
  ND2D1BWP30P140LVT U14193 ( .A1(n9721), .A2(n9720), .ZN(N3739) );
  AOI22D1BWP30P140LVT U14194 ( .A1(i_data_bus[360]), .A2(n9730), .B1(
        i_data_bus[328]), .B2(n9731), .ZN(n9723) );
  AOI22D1BWP30P140LVT U14195 ( .A1(i_data_bus[264]), .A2(n6219), .B1(
        i_data_bus[296]), .B2(n9732), .ZN(n9722) );
  ND2D1BWP30P140LVT U14196 ( .A1(n9723), .A2(n9722), .ZN(N3735) );
  AOI22D1BWP30P140LVT U14197 ( .A1(i_data_bus[262]), .A2(n6219), .B1(
        i_data_bus[326]), .B2(n9731), .ZN(n9725) );
  AOI22D1BWP30P140LVT U14198 ( .A1(i_data_bus[358]), .A2(n9730), .B1(
        i_data_bus[294]), .B2(n9732), .ZN(n9724) );
  ND2D1BWP30P140LVT U14199 ( .A1(n9725), .A2(n9724), .ZN(N3733) );
  AOI22D1BWP30P140LVT U14200 ( .A1(i_data_bus[259]), .A2(n6219), .B1(
        i_data_bus[323]), .B2(n9731), .ZN(n9727) );
  AOI22D1BWP30P140LVT U14201 ( .A1(i_data_bus[355]), .A2(n9730), .B1(
        i_data_bus[291]), .B2(n9732), .ZN(n9726) );
  ND2D1BWP30P140LVT U14202 ( .A1(n9727), .A2(n9726), .ZN(N3730) );
  AOI22D1BWP30P140LVT U14203 ( .A1(i_data_bus[320]), .A2(n9731), .B1(
        i_data_bus[352]), .B2(n9730), .ZN(n9729) );
  AOI22D1BWP30P140LVT U14204 ( .A1(i_data_bus[256]), .A2(n6219), .B1(
        i_data_bus[288]), .B2(n9732), .ZN(n9728) );
  ND2D1BWP30P140LVT U14205 ( .A1(n9729), .A2(n9728), .ZN(N3727) );
  AOI22D1BWP30P140LVT U14206 ( .A1(i_data_bus[340]), .A2(n9731), .B1(
        i_data_bus[372]), .B2(n9730), .ZN(n9734) );
  AOI22D1BWP30P140LVT U14207 ( .A1(i_data_bus[276]), .A2(n6219), .B1(
        i_data_bus[308]), .B2(n9732), .ZN(n9733) );
  ND2D1BWP30P140LVT U14208 ( .A1(n9734), .A2(n9733), .ZN(N3747) );
  AOI22D1BWP30P140LVT U14209 ( .A1(i_data_bus[317]), .A2(n9758), .B1(
        i_data_bus[285]), .B2(n9756), .ZN(n9736) );
  AOI22D1BWP30P140LVT U14210 ( .A1(i_data_bus[349]), .A2(n9755), .B1(
        i_data_bus[381]), .B2(n9757), .ZN(n9735) );
  ND2D1BWP30P140LVT U14211 ( .A1(n9736), .A2(n9735), .ZN(N5246) );
  AOI22D1BWP30P140LVT U14212 ( .A1(i_data_bus[289]), .A2(n9758), .B1(
        i_data_bus[257]), .B2(n9756), .ZN(n9738) );
  AOI22D1BWP30P140LVT U14213 ( .A1(i_data_bus[321]), .A2(n9755), .B1(
        i_data_bus[353]), .B2(n9757), .ZN(n9737) );
  ND2D1BWP30P140LVT U14214 ( .A1(n9738), .A2(n9737), .ZN(N5218) );
  AOI22D1BWP30P140LVT U14215 ( .A1(i_data_bus[322]), .A2(n9755), .B1(
        i_data_bus[258]), .B2(n9756), .ZN(n9740) );
  AOI22D1BWP30P140LVT U14216 ( .A1(i_data_bus[290]), .A2(n9758), .B1(
        i_data_bus[354]), .B2(n9757), .ZN(n9739) );
  ND2D1BWP30P140LVT U14217 ( .A1(n9740), .A2(n9739), .ZN(N5219) );
  AOI22D1BWP30P140LVT U14218 ( .A1(i_data_bus[304]), .A2(n9758), .B1(
        i_data_bus[336]), .B2(n9755), .ZN(n9742) );
  AOI22D1BWP30P140LVT U14219 ( .A1(i_data_bus[272]), .A2(n9756), .B1(
        i_data_bus[368]), .B2(n9757), .ZN(n9741) );
  ND2D1BWP30P140LVT U14220 ( .A1(n9742), .A2(n9741), .ZN(N5233) );
  AOI22D1BWP30P140LVT U14221 ( .A1(i_data_bus[351]), .A2(n9755), .B1(
        i_data_bus[287]), .B2(n9756), .ZN(n9744) );
  AOI22D1BWP30P140LVT U14222 ( .A1(i_data_bus[319]), .A2(n9758), .B1(
        i_data_bus[383]), .B2(n9757), .ZN(n9743) );
  ND2D1BWP30P140LVT U14223 ( .A1(n9744), .A2(n9743), .ZN(N5248) );
  AOI22D1BWP30P140LVT U14224 ( .A1(i_data_bus[281]), .A2(n9756), .B1(
        i_data_bus[345]), .B2(n9755), .ZN(n9746) );
  AOI22D1BWP30P140LVT U14225 ( .A1(i_data_bus[313]), .A2(n9758), .B1(
        i_data_bus[377]), .B2(n9757), .ZN(n9745) );
  ND2D1BWP30P140LVT U14226 ( .A1(n9746), .A2(n9745), .ZN(N5242) );
  AOI22D1BWP30P140LVT U14227 ( .A1(i_data_bus[277]), .A2(n9756), .B1(
        i_data_bus[341]), .B2(n9755), .ZN(n9748) );
  AOI22D1BWP30P140LVT U14228 ( .A1(i_data_bus[309]), .A2(n9758), .B1(
        i_data_bus[373]), .B2(n9757), .ZN(n9747) );
  ND2D1BWP30P140LVT U14229 ( .A1(n9748), .A2(n9747), .ZN(N5238) );
  AOI22D1BWP30P140LVT U14230 ( .A1(i_data_bus[274]), .A2(n9756), .B1(
        i_data_bus[306]), .B2(n9758), .ZN(n9750) );
  AOI22D1BWP30P140LVT U14231 ( .A1(i_data_bus[338]), .A2(n9755), .B1(
        i_data_bus[370]), .B2(n9757), .ZN(n9749) );
  ND2D1BWP30P140LVT U14232 ( .A1(n9750), .A2(n9749), .ZN(N5235) );
  AOI22D1BWP30P140LVT U14233 ( .A1(i_data_bus[273]), .A2(n9756), .B1(
        i_data_bus[305]), .B2(n9758), .ZN(n9752) );
  AOI22D1BWP30P140LVT U14234 ( .A1(i_data_bus[337]), .A2(n9755), .B1(
        i_data_bus[369]), .B2(n9757), .ZN(n9751) );
  ND2D1BWP30P140LVT U14235 ( .A1(n9752), .A2(n9751), .ZN(N5234) );
  AOI22D1BWP30P140LVT U14236 ( .A1(i_data_bus[298]), .A2(n9758), .B1(
        i_data_bus[330]), .B2(n9755), .ZN(n9754) );
  AOI22D1BWP30P140LVT U14237 ( .A1(i_data_bus[266]), .A2(n9756), .B1(
        i_data_bus[362]), .B2(n9757), .ZN(n9753) );
  ND2D1BWP30P140LVT U14238 ( .A1(n9754), .A2(n9753), .ZN(N5227) );
  AOI22D1BWP30P140LVT U14239 ( .A1(i_data_bus[263]), .A2(n9756), .B1(
        i_data_bus[327]), .B2(n9755), .ZN(n9760) );
  AOI22D1BWP30P140LVT U14240 ( .A1(i_data_bus[295]), .A2(n9758), .B1(
        i_data_bus[359]), .B2(n9757), .ZN(n9759) );
  ND2D1BWP30P140LVT U14241 ( .A1(n9760), .A2(n9759), .ZN(N5224) );
  AOI22D1BWP30P140LVT U14242 ( .A1(i_data_bus[340]), .A2(n9774), .B1(
        i_data_bus[372]), .B2(n9773), .ZN(n9762) );
  AOI22D1BWP30P140LVT U14243 ( .A1(i_data_bus[276]), .A2(n6216), .B1(
        i_data_bus[308]), .B2(n9775), .ZN(n9761) );
  ND2D1BWP30P140LVT U14244 ( .A1(n9762), .A2(n9761), .ZN(N2513) );
  AOI22D1BWP30P140LVT U14245 ( .A1(i_data_bus[275]), .A2(n6216), .B1(
        i_data_bus[339]), .B2(n9774), .ZN(n9764) );
  AOI22D1BWP30P140LVT U14246 ( .A1(i_data_bus[371]), .A2(n9773), .B1(
        i_data_bus[307]), .B2(n9775), .ZN(n9763) );
  ND2D1BWP30P140LVT U14247 ( .A1(n9764), .A2(n9763), .ZN(N2512) );
  AOI22D1BWP30P140LVT U14248 ( .A1(i_data_bus[262]), .A2(n6216), .B1(
        i_data_bus[326]), .B2(n9774), .ZN(n9766) );
  AOI22D1BWP30P140LVT U14249 ( .A1(i_data_bus[358]), .A2(n9773), .B1(
        i_data_bus[294]), .B2(n9775), .ZN(n9765) );
  ND2D1BWP30P140LVT U14250 ( .A1(n9766), .A2(n9765), .ZN(N2499) );
  AOI22D1BWP30P140LVT U14251 ( .A1(i_data_bus[320]), .A2(n9774), .B1(
        i_data_bus[352]), .B2(n9773), .ZN(n9768) );
  AOI22D1BWP30P140LVT U14252 ( .A1(i_data_bus[256]), .A2(n6216), .B1(
        i_data_bus[288]), .B2(n9775), .ZN(n9767) );
  ND2D1BWP30P140LVT U14253 ( .A1(n9768), .A2(n9767), .ZN(N2493) );
  AOI22D1BWP30P140LVT U14254 ( .A1(i_data_bus[334]), .A2(n9774), .B1(
        i_data_bus[366]), .B2(n9773), .ZN(n9770) );
  AOI22D1BWP30P140LVT U14255 ( .A1(i_data_bus[270]), .A2(n6216), .B1(
        i_data_bus[302]), .B2(n9775), .ZN(n9769) );
  ND2D1BWP30P140LVT U14256 ( .A1(n9770), .A2(n9769), .ZN(N2507) );
  AOI22D1BWP30P140LVT U14257 ( .A1(i_data_bus[337]), .A2(n9774), .B1(
        i_data_bus[273]), .B2(n6216), .ZN(n9772) );
  AOI22D1BWP30P140LVT U14258 ( .A1(i_data_bus[369]), .A2(n9773), .B1(
        i_data_bus[305]), .B2(n9775), .ZN(n9771) );
  ND2D1BWP30P140LVT U14259 ( .A1(n9772), .A2(n9771), .ZN(N2510) );
  AOI22D1BWP30P140LVT U14260 ( .A1(i_data_bus[338]), .A2(n9774), .B1(
        i_data_bus[370]), .B2(n9773), .ZN(n9777) );
  AOI22D1BWP30P140LVT U14261 ( .A1(i_data_bus[274]), .A2(n6216), .B1(
        i_data_bus[306]), .B2(n9775), .ZN(n9776) );
  ND2D1BWP30P140LVT U14262 ( .A1(n9777), .A2(n9776), .ZN(N2511) );
  AOI22D1BWP30P140LVT U14263 ( .A1(i_data_bus[70]), .A2(n9790), .B1(
        i_data_bus[38]), .B2(n9791), .ZN(n9779) );
  AOI22D1BWP30P140LVT U14264 ( .A1(i_data_bus[6]), .A2(n6223), .B1(
        i_data_bus[102]), .B2(n9792), .ZN(n9778) );
  ND2D1BWP30P140LVT U14265 ( .A1(n9779), .A2(n9778), .ZN(N8749) );
  AOI22D1BWP30P140LVT U14266 ( .A1(i_data_bus[45]), .A2(n9791), .B1(
        i_data_bus[77]), .B2(n9790), .ZN(n9781) );
  AOI22D1BWP30P140LVT U14267 ( .A1(i_data_bus[13]), .A2(n6223), .B1(
        i_data_bus[109]), .B2(n9792), .ZN(n9780) );
  ND2D1BWP30P140LVT U14268 ( .A1(n9781), .A2(n9780), .ZN(N8756) );
  AOI22D1BWP30P140LVT U14269 ( .A1(i_data_bus[43]), .A2(n9791), .B1(
        i_data_bus[75]), .B2(n9790), .ZN(n9783) );
  AOI22D1BWP30P140LVT U14270 ( .A1(i_data_bus[11]), .A2(n6223), .B1(
        i_data_bus[107]), .B2(n9792), .ZN(n9782) );
  ND2D1BWP30P140LVT U14271 ( .A1(n9783), .A2(n9782), .ZN(N8754) );
  AOI22D1BWP30P140LVT U14272 ( .A1(i_data_bus[50]), .A2(n9791), .B1(
        i_data_bus[82]), .B2(n9790), .ZN(n9785) );
  AOI22D1BWP30P140LVT U14273 ( .A1(i_data_bus[18]), .A2(n6223), .B1(
        i_data_bus[114]), .B2(n9792), .ZN(n9784) );
  ND2D1BWP30P140LVT U14274 ( .A1(n9785), .A2(n9784), .ZN(N8761) );
  AOI22D1BWP30P140LVT U14275 ( .A1(i_data_bus[61]), .A2(n9791), .B1(
        i_data_bus[29]), .B2(n6223), .ZN(n9787) );
  AOI22D1BWP30P140LVT U14276 ( .A1(i_data_bus[93]), .A2(n9790), .B1(
        i_data_bus[125]), .B2(n9792), .ZN(n9786) );
  ND2D1BWP30P140LVT U14277 ( .A1(n9787), .A2(n9786), .ZN(N8772) );
  AOI22D1BWP30P140LVT U14278 ( .A1(i_data_bus[12]), .A2(n6223), .B1(
        i_data_bus[44]), .B2(n9791), .ZN(n9789) );
  AOI22D1BWP30P140LVT U14279 ( .A1(i_data_bus[76]), .A2(n9790), .B1(
        i_data_bus[108]), .B2(n9792), .ZN(n9788) );
  ND2D1BWP30P140LVT U14280 ( .A1(n9789), .A2(n9788), .ZN(N8755) );
  AOI22D1BWP30P140LVT U14281 ( .A1(i_data_bus[53]), .A2(n9791), .B1(
        i_data_bus[85]), .B2(n9790), .ZN(n9794) );
  AOI22D1BWP30P140LVT U14282 ( .A1(i_data_bus[21]), .A2(n6223), .B1(
        i_data_bus[117]), .B2(n9792), .ZN(n9793) );
  ND2D1BWP30P140LVT U14283 ( .A1(n9794), .A2(n9793), .ZN(N8764) );
  AOI22D1BWP30P140LVT U14284 ( .A1(i_data_bus[270]), .A2(n10052), .B1(
        i_data_bus[302]), .B2(n10053), .ZN(n9796) );
  AOI22D1BWP30P140LVT U14285 ( .A1(i_data_bus[334]), .A2(n10054), .B1(
        i_data_bus[366]), .B2(n10051), .ZN(n9795) );
  ND2D1BWP30P140LVT U14286 ( .A1(n9796), .A2(n9795), .ZN(N6465) );
  AOI22D1BWP30P140LVT U14287 ( .A1(i_data_bus[351]), .A2(n9844), .B1(
        i_data_bus[287]), .B2(n9846), .ZN(n9798) );
  AOI22D1BWP30P140LVT U14288 ( .A1(i_data_bus[319]), .A2(n9843), .B1(
        i_data_bus[383]), .B2(n9845), .ZN(n9797) );
  ND2D1BWP30P140LVT U14289 ( .A1(n9798), .A2(n9797), .ZN(N7972) );
  AOI22D1BWP30P140LVT U14290 ( .A1(i_data_bus[292]), .A2(n10053), .B1(
        i_data_bus[324]), .B2(n10054), .ZN(n9800) );
  AOI22D1BWP30P140LVT U14291 ( .A1(i_data_bus[260]), .A2(n10052), .B1(
        i_data_bus[356]), .B2(n10051), .ZN(n9799) );
  ND2D1BWP30P140LVT U14292 ( .A1(n9800), .A2(n9799), .ZN(N6455) );
  AOI22D1BWP30P140LVT U14293 ( .A1(i_data_bus[263]), .A2(n10052), .B1(
        i_data_bus[327]), .B2(n10054), .ZN(n9802) );
  AOI22D1BWP30P140LVT U14294 ( .A1(i_data_bus[295]), .A2(n10053), .B1(
        i_data_bus[359]), .B2(n10051), .ZN(n9801) );
  ND2D1BWP30P140LVT U14295 ( .A1(n9802), .A2(n9801), .ZN(N6458) );
  AOI22D1BWP30P140LVT U14296 ( .A1(i_data_bus[276]), .A2(n10052), .B1(
        i_data_bus[308]), .B2(n10053), .ZN(n9804) );
  AOI22D1BWP30P140LVT U14297 ( .A1(i_data_bus[340]), .A2(n10054), .B1(
        i_data_bus[372]), .B2(n10051), .ZN(n9803) );
  ND2D1BWP30P140LVT U14298 ( .A1(n9804), .A2(n9803), .ZN(N6471) );
  AOI22D1BWP30P140LVT U14299 ( .A1(i_data_bus[326]), .A2(n10054), .B1(
        i_data_bus[294]), .B2(n10053), .ZN(n9806) );
  AOI22D1BWP30P140LVT U14300 ( .A1(i_data_bus[262]), .A2(n10052), .B1(
        i_data_bus[358]), .B2(n10051), .ZN(n9805) );
  ND2D1BWP30P140LVT U14301 ( .A1(n9806), .A2(n9805), .ZN(N6457) );
  AOI22D1BWP30P140LVT U14302 ( .A1(i_data_bus[322]), .A2(n9844), .B1(
        i_data_bus[258]), .B2(n9846), .ZN(n9808) );
  AOI22D1BWP30P140LVT U14303 ( .A1(i_data_bus[290]), .A2(n9843), .B1(
        i_data_bus[354]), .B2(n9845), .ZN(n9807) );
  ND2D1BWP30P140LVT U14304 ( .A1(n9808), .A2(n9807), .ZN(N7943) );
  AOI22D1BWP30P140LVT U14305 ( .A1(i_data_bus[315]), .A2(n9843), .B1(
        i_data_bus[347]), .B2(n9844), .ZN(n9810) );
  AOI22D1BWP30P140LVT U14306 ( .A1(i_data_bus[283]), .A2(n9846), .B1(
        i_data_bus[379]), .B2(n9845), .ZN(n9809) );
  ND2D1BWP30P140LVT U14307 ( .A1(n9810), .A2(n9809), .ZN(N7968) );
  AOI22D1BWP30P140LVT U14308 ( .A1(i_data_bus[278]), .A2(n10052), .B1(
        i_data_bus[310]), .B2(n10053), .ZN(n9812) );
  AOI22D1BWP30P140LVT U14309 ( .A1(i_data_bus[342]), .A2(n10054), .B1(
        i_data_bus[374]), .B2(n10051), .ZN(n9811) );
  ND2D1BWP30P140LVT U14310 ( .A1(n9812), .A2(n9811), .ZN(N6473) );
  AOI22D1BWP30P140LVT U14311 ( .A1(i_data_bus[283]), .A2(n10052), .B1(
        i_data_bus[347]), .B2(n10054), .ZN(n9814) );
  AOI22D1BWP30P140LVT U14312 ( .A1(i_data_bus[315]), .A2(n10053), .B1(
        i_data_bus[379]), .B2(n10051), .ZN(n9813) );
  ND2D1BWP30P140LVT U14313 ( .A1(n9814), .A2(n9813), .ZN(N6478) );
  AOI22D1BWP30P140LVT U14314 ( .A1(i_data_bus[256]), .A2(n10052), .B1(
        i_data_bus[320]), .B2(n10054), .ZN(n9816) );
  AOI22D1BWP30P140LVT U14315 ( .A1(i_data_bus[288]), .A2(n10053), .B1(
        i_data_bus[352]), .B2(n10051), .ZN(n9815) );
  ND2D1BWP30P140LVT U14316 ( .A1(n9816), .A2(n9815), .ZN(N6451) );
  AOI22D1BWP30P140LVT U14317 ( .A1(i_data_bus[319]), .A2(n10053), .B1(
        i_data_bus[287]), .B2(n10052), .ZN(n9818) );
  AOI22D1BWP30P140LVT U14318 ( .A1(i_data_bus[351]), .A2(n10054), .B1(
        i_data_bus[383]), .B2(n10051), .ZN(n9817) );
  ND2D1BWP30P140LVT U14319 ( .A1(n9818), .A2(n9817), .ZN(N6482) );
  AOI22D1BWP30P140LVT U14320 ( .A1(i_data_bus[278]), .A2(n9846), .B1(
        i_data_bus[310]), .B2(n9843), .ZN(n9820) );
  AOI22D1BWP30P140LVT U14321 ( .A1(i_data_bus[342]), .A2(n9844), .B1(
        i_data_bus[374]), .B2(n9845), .ZN(n9819) );
  ND2D1BWP30P140LVT U14322 ( .A1(n9820), .A2(n9819), .ZN(N7963) );
  AOI22D1BWP30P140LVT U14323 ( .A1(i_data_bus[350]), .A2(n10054), .B1(
        i_data_bus[318]), .B2(n10053), .ZN(n9822) );
  AOI22D1BWP30P140LVT U14324 ( .A1(i_data_bus[286]), .A2(n10052), .B1(
        i_data_bus[382]), .B2(n10051), .ZN(n9821) );
  ND2D1BWP30P140LVT U14325 ( .A1(n9822), .A2(n9821), .ZN(N6481) );
  AOI22D1BWP30P140LVT U14326 ( .A1(i_data_bus[322]), .A2(n10054), .B1(
        i_data_bus[290]), .B2(n10053), .ZN(n9824) );
  AOI22D1BWP30P140LVT U14327 ( .A1(i_data_bus[258]), .A2(n10052), .B1(
        i_data_bus[354]), .B2(n10051), .ZN(n9823) );
  ND2D1BWP30P140LVT U14328 ( .A1(n9824), .A2(n9823), .ZN(N6453) );
  AOI22D1BWP30P140LVT U14329 ( .A1(i_data_bus[281]), .A2(n9846), .B1(
        i_data_bus[345]), .B2(n9844), .ZN(n9826) );
  AOI22D1BWP30P140LVT U14330 ( .A1(i_data_bus[313]), .A2(n9843), .B1(
        i_data_bus[377]), .B2(n9845), .ZN(n9825) );
  ND2D1BWP30P140LVT U14331 ( .A1(n9826), .A2(n9825), .ZN(N7966) );
  AOI22D1BWP30P140LVT U14332 ( .A1(i_data_bus[339]), .A2(n9844), .B1(
        i_data_bus[307]), .B2(n9843), .ZN(n9828) );
  AOI22D1BWP30P140LVT U14333 ( .A1(i_data_bus[275]), .A2(n9846), .B1(
        i_data_bus[371]), .B2(n9845), .ZN(n9827) );
  ND2D1BWP30P140LVT U14334 ( .A1(n9828), .A2(n9827), .ZN(N7960) );
  AOI22D1BWP30P140LVT U14335 ( .A1(i_data_bus[303]), .A2(n9843), .B1(
        i_data_bus[335]), .B2(n9844), .ZN(n9830) );
  AOI22D1BWP30P140LVT U14336 ( .A1(i_data_bus[271]), .A2(n9846), .B1(
        i_data_bus[367]), .B2(n9845), .ZN(n9829) );
  ND2D1BWP30P140LVT U14337 ( .A1(n9830), .A2(n9829), .ZN(N7956) );
  AOI22D1BWP30P140LVT U14338 ( .A1(i_data_bus[298]), .A2(n9843), .B1(
        i_data_bus[330]), .B2(n9844), .ZN(n9832) );
  AOI22D1BWP30P140LVT U14339 ( .A1(i_data_bus[266]), .A2(n9846), .B1(
        i_data_bus[362]), .B2(n9845), .ZN(n9831) );
  ND2D1BWP30P140LVT U14340 ( .A1(n9832), .A2(n9831), .ZN(N7951) );
  AOI22D1BWP30P140LVT U14341 ( .A1(i_data_bus[256]), .A2(n9846), .B1(
        i_data_bus[288]), .B2(n9843), .ZN(n9834) );
  AOI22D1BWP30P140LVT U14342 ( .A1(i_data_bus[320]), .A2(n9844), .B1(
        i_data_bus[352]), .B2(n9845), .ZN(n9833) );
  ND2D1BWP30P140LVT U14343 ( .A1(n9834), .A2(n9833), .ZN(N7941) );
  AOI22D1BWP30P140LVT U14344 ( .A1(i_data_bus[302]), .A2(n9843), .B1(
        i_data_bus[334]), .B2(n9844), .ZN(n9836) );
  AOI22D1BWP30P140LVT U14345 ( .A1(i_data_bus[270]), .A2(n9846), .B1(
        i_data_bus[366]), .B2(n9845), .ZN(n9835) );
  ND2D1BWP30P140LVT U14346 ( .A1(n9836), .A2(n9835), .ZN(N7955) );
  AOI22D1BWP30P140LVT U14347 ( .A1(i_data_bus[338]), .A2(n9844), .B1(
        i_data_bus[306]), .B2(n9843), .ZN(n9838) );
  AOI22D1BWP30P140LVT U14348 ( .A1(i_data_bus[274]), .A2(n9846), .B1(
        i_data_bus[370]), .B2(n9845), .ZN(n9837) );
  ND2D1BWP30P140LVT U14349 ( .A1(n9838), .A2(n9837), .ZN(N7959) );
  AOI22D1BWP30P140LVT U14350 ( .A1(i_data_bus[282]), .A2(n10052), .B1(
        i_data_bus[314]), .B2(n10053), .ZN(n9840) );
  AOI22D1BWP30P140LVT U14351 ( .A1(i_data_bus[346]), .A2(n10054), .B1(
        i_data_bus[378]), .B2(n10051), .ZN(n9839) );
  ND2D1BWP30P140LVT U14352 ( .A1(n9840), .A2(n9839), .ZN(N6477) );
  AOI22D1BWP30P140LVT U14353 ( .A1(i_data_bus[274]), .A2(n10052), .B1(
        i_data_bus[338]), .B2(n10054), .ZN(n9842) );
  AOI22D1BWP30P140LVT U14354 ( .A1(i_data_bus[306]), .A2(n10053), .B1(
        i_data_bus[370]), .B2(n10051), .ZN(n9841) );
  ND2D1BWP30P140LVT U14355 ( .A1(n9842), .A2(n9841), .ZN(N6469) );
  AOI22D1BWP30P140LVT U14356 ( .A1(i_data_bus[326]), .A2(n9844), .B1(
        i_data_bus[294]), .B2(n9843), .ZN(n9848) );
  AOI22D1BWP30P140LVT U14357 ( .A1(i_data_bus[262]), .A2(n9846), .B1(
        i_data_bus[358]), .B2(n9845), .ZN(n9847) );
  ND2D1BWP30P140LVT U14358 ( .A1(n9848), .A2(n9847), .ZN(N7947) );
  AOI22D1BWP30P140LVT U14359 ( .A1(i_data_bus[272]), .A2(n10052), .B1(
        i_data_bus[336]), .B2(n10054), .ZN(n9850) );
  AOI22D1BWP30P140LVT U14360 ( .A1(i_data_bus[304]), .A2(n10053), .B1(
        i_data_bus[368]), .B2(n10051), .ZN(n9849) );
  ND2D1BWP30P140LVT U14361 ( .A1(n9850), .A2(n9849), .ZN(N6467) );
  AOI22D1BWP30P140LVT U14362 ( .A1(i_data_bus[357]), .A2(n9877), .B1(
        i_data_bus[325]), .B2(n9879), .ZN(n9852) );
  AOI22D1BWP30P140LVT U14363 ( .A1(i_data_bus[261]), .A2(n6217), .B1(
        i_data_bus[293]), .B2(n9878), .ZN(n9851) );
  ND2D1BWP30P140LVT U14364 ( .A1(n9852), .A2(n9851), .ZN(N10670) );
  AOI22D1BWP30P140LVT U14365 ( .A1(i_data_bus[275]), .A2(n6217), .B1(
        i_data_bus[339]), .B2(n9879), .ZN(n9854) );
  AOI22D1BWP30P140LVT U14366 ( .A1(i_data_bus[371]), .A2(n9877), .B1(
        i_data_bus[307]), .B2(n9878), .ZN(n9853) );
  ND2D1BWP30P140LVT U14367 ( .A1(n9854), .A2(n9853), .ZN(N10684) );
  AOI22D1BWP30P140LVT U14368 ( .A1(i_data_bus[346]), .A2(n10275), .B1(
        i_data_bus[378]), .B2(n10277), .ZN(n9856) );
  AOI22D1BWP30P140LVT U14369 ( .A1(i_data_bus[282]), .A2(n6227), .B1(
        i_data_bus[314]), .B2(n10276), .ZN(n9855) );
  ND2D1BWP30P140LVT U14370 ( .A1(n9856), .A2(n9855), .ZN(N9201) );
  AOI22D1BWP30P140LVT U14371 ( .A1(i_data_bus[259]), .A2(n6227), .B1(
        i_data_bus[355]), .B2(n10277), .ZN(n9858) );
  AOI22D1BWP30P140LVT U14372 ( .A1(i_data_bus[323]), .A2(n10275), .B1(
        i_data_bus[291]), .B2(n10276), .ZN(n9857) );
  ND2D1BWP30P140LVT U14373 ( .A1(n9858), .A2(n9857), .ZN(N9178) );
  AOI22D1BWP30P140LVT U14374 ( .A1(i_data_bus[280]), .A2(n6227), .B1(
        i_data_bus[344]), .B2(n10275), .ZN(n9860) );
  AOI22D1BWP30P140LVT U14375 ( .A1(i_data_bus[376]), .A2(n10277), .B1(
        i_data_bus[312]), .B2(n10276), .ZN(n9859) );
  ND2D1BWP30P140LVT U14376 ( .A1(n9860), .A2(n9859), .ZN(N9199) );
  AOI22D1BWP30P140LVT U14377 ( .A1(i_data_bus[360]), .A2(n10277), .B1(
        i_data_bus[328]), .B2(n10275), .ZN(n9862) );
  AOI22D1BWP30P140LVT U14378 ( .A1(i_data_bus[264]), .A2(n6227), .B1(
        i_data_bus[296]), .B2(n10276), .ZN(n9861) );
  ND2D1BWP30P140LVT U14379 ( .A1(n9862), .A2(n9861), .ZN(N9183) );
  AOI22D1BWP30P140LVT U14380 ( .A1(i_data_bus[356]), .A2(n10277), .B1(
        i_data_bus[324]), .B2(n10275), .ZN(n9864) );
  AOI22D1BWP30P140LVT U14381 ( .A1(i_data_bus[260]), .A2(n6227), .B1(
        i_data_bus[292]), .B2(n10276), .ZN(n9863) );
  ND2D1BWP30P140LVT U14382 ( .A1(n9864), .A2(n9863), .ZN(N9179) );
  AOI22D1BWP30P140LVT U14383 ( .A1(i_data_bus[274]), .A2(n6217), .B1(
        i_data_bus[370]), .B2(n9877), .ZN(n9866) );
  AOI22D1BWP30P140LVT U14384 ( .A1(i_data_bus[338]), .A2(n9879), .B1(
        i_data_bus[306]), .B2(n9878), .ZN(n9865) );
  ND2D1BWP30P140LVT U14385 ( .A1(n9866), .A2(n9865), .ZN(N10683) );
  AOI22D1BWP30P140LVT U14386 ( .A1(i_data_bus[275]), .A2(n6227), .B1(
        i_data_bus[339]), .B2(n10275), .ZN(n9868) );
  AOI22D1BWP30P140LVT U14387 ( .A1(i_data_bus[371]), .A2(n10277), .B1(
        i_data_bus[307]), .B2(n10276), .ZN(n9867) );
  ND2D1BWP30P140LVT U14388 ( .A1(n9868), .A2(n9867), .ZN(N9194) );
  AOI22D1BWP30P140LVT U14389 ( .A1(i_data_bus[331]), .A2(n10275), .B1(
        i_data_bus[267]), .B2(n6227), .ZN(n9870) );
  AOI22D1BWP30P140LVT U14390 ( .A1(i_data_bus[363]), .A2(n10277), .B1(
        i_data_bus[299]), .B2(n10276), .ZN(n9869) );
  ND2D1BWP30P140LVT U14391 ( .A1(n9870), .A2(n9869), .ZN(N9186) );
  AOI22D1BWP30P140LVT U14392 ( .A1(i_data_bus[262]), .A2(n6227), .B1(
        i_data_bus[358]), .B2(n10277), .ZN(n9872) );
  AOI22D1BWP30P140LVT U14393 ( .A1(i_data_bus[326]), .A2(n10275), .B1(
        i_data_bus[294]), .B2(n10276), .ZN(n9871) );
  ND2D1BWP30P140LVT U14394 ( .A1(n9872), .A2(n9871), .ZN(N9181) );
  AOI22D1BWP30P140LVT U14395 ( .A1(i_data_bus[269]), .A2(n6217), .B1(
        i_data_bus[333]), .B2(n9879), .ZN(n9874) );
  AOI22D1BWP30P140LVT U14396 ( .A1(i_data_bus[365]), .A2(n9877), .B1(
        i_data_bus[301]), .B2(n9878), .ZN(n9873) );
  ND2D1BWP30P140LVT U14397 ( .A1(n9874), .A2(n9873), .ZN(N10678) );
  AOI22D1BWP30P140LVT U14398 ( .A1(i_data_bus[328]), .A2(n9879), .B1(
        i_data_bus[264]), .B2(n6217), .ZN(n9876) );
  AOI22D1BWP30P140LVT U14399 ( .A1(i_data_bus[360]), .A2(n9877), .B1(
        i_data_bus[296]), .B2(n9878), .ZN(n9875) );
  ND2D1BWP30P140LVT U14400 ( .A1(n9876), .A2(n9875), .ZN(N10673) );
  AOI22D1BWP30P140LVT U14401 ( .A1(i_data_bus[256]), .A2(n6217), .B1(
        i_data_bus[352]), .B2(n9877), .ZN(n9881) );
  AOI22D1BWP30P140LVT U14402 ( .A1(i_data_bus[320]), .A2(n9879), .B1(
        i_data_bus[288]), .B2(n9878), .ZN(n9880) );
  ND2D1BWP30P140LVT U14403 ( .A1(n9881), .A2(n9880), .ZN(N10665) );
  AOI22D1BWP30P140LVT U14404 ( .A1(i_data_bus[319]), .A2(n10276), .B1(
        i_data_bus[287]), .B2(n6227), .ZN(n9883) );
  AOI22D1BWP30P140LVT U14405 ( .A1(i_data_bus[351]), .A2(n10275), .B1(
        i_data_bus[383]), .B2(n10277), .ZN(n9882) );
  ND2D1BWP30P140LVT U14406 ( .A1(n9883), .A2(n9882), .ZN(N9206) );
  AOI22D1BWP30P140LVT U14407 ( .A1(i_data_bus[309]), .A2(n10276), .B1(
        i_data_bus[277]), .B2(n6227), .ZN(n9885) );
  AOI22D1BWP30P140LVT U14408 ( .A1(i_data_bus[373]), .A2(n10277), .B1(
        i_data_bus[341]), .B2(n10275), .ZN(n9884) );
  ND2D1BWP30P140LVT U14409 ( .A1(n9885), .A2(n9884), .ZN(N9196) );
  AOI22D1BWP30P140LVT U14410 ( .A1(i_data_bus[313]), .A2(n10276), .B1(
        i_data_bus[281]), .B2(n6227), .ZN(n9887) );
  AOI22D1BWP30P140LVT U14411 ( .A1(i_data_bus[377]), .A2(n10277), .B1(
        i_data_bus[345]), .B2(n10275), .ZN(n9886) );
  ND2D1BWP30P140LVT U14412 ( .A1(n9887), .A2(n9886), .ZN(N9200) );
  AOI22D1BWP30P140LVT U14413 ( .A1(i_data_bus[372]), .A2(n10277), .B1(
        i_data_bus[276]), .B2(n6227), .ZN(n9889) );
  AOI22D1BWP30P140LVT U14414 ( .A1(i_data_bus[340]), .A2(n10275), .B1(
        i_data_bus[308]), .B2(n10276), .ZN(n9888) );
  ND2D1BWP30P140LVT U14415 ( .A1(n9889), .A2(n9888), .ZN(N9195) );
  AOI22D1BWP30P140LVT U14416 ( .A1(i_data_bus[361]), .A2(n10277), .B1(
        i_data_bus[265]), .B2(n6227), .ZN(n9891) );
  AOI22D1BWP30P140LVT U14417 ( .A1(i_data_bus[297]), .A2(n10276), .B1(
        i_data_bus[329]), .B2(n10275), .ZN(n9890) );
  ND2D1BWP30P140LVT U14418 ( .A1(n9891), .A2(n9890), .ZN(N9184) );
  AOI22D1BWP30P140LVT U14419 ( .A1(i_data_bus[337]), .A2(n10275), .B1(
        i_data_bus[273]), .B2(n6227), .ZN(n9893) );
  AOI22D1BWP30P140LVT U14420 ( .A1(i_data_bus[369]), .A2(n10277), .B1(
        i_data_bus[305]), .B2(n10276), .ZN(n9892) );
  ND2D1BWP30P140LVT U14421 ( .A1(n9893), .A2(n9892), .ZN(N9192) );
  AOI22D1BWP30P140LVT U14422 ( .A1(i_data_bus[321]), .A2(n10275), .B1(
        i_data_bus[257]), .B2(n6227), .ZN(n9895) );
  AOI22D1BWP30P140LVT U14423 ( .A1(i_data_bus[289]), .A2(n10276), .B1(
        i_data_bus[353]), .B2(n10277), .ZN(n9894) );
  ND2D1BWP30P140LVT U14424 ( .A1(n9895), .A2(n9894), .ZN(N9176) );
  AOI22D1BWP30P140LVT U14425 ( .A1(i_data_bus[84]), .A2(n9914), .B1(
        i_data_bus[116]), .B2(n9915), .ZN(n9897) );
  AOI22D1BWP30P140LVT U14426 ( .A1(i_data_bus[20]), .A2(n6218), .B1(
        i_data_bus[52]), .B2(n9916), .ZN(n9896) );
  ND2D1BWP30P140LVT U14427 ( .A1(n9897), .A2(n9896), .ZN(N3315) );
  AOI22D1BWP30P140LVT U14428 ( .A1(i_data_bus[14]), .A2(n6218), .B1(
        i_data_bus[110]), .B2(n9915), .ZN(n9899) );
  AOI22D1BWP30P140LVT U14429 ( .A1(i_data_bus[78]), .A2(n9914), .B1(
        i_data_bus[46]), .B2(n9916), .ZN(n9898) );
  ND2D1BWP30P140LVT U14430 ( .A1(n9899), .A2(n9898), .ZN(N3309) );
  AOI22D1BWP30P140LVT U14431 ( .A1(i_data_bus[7]), .A2(n6218), .B1(
        i_data_bus[71]), .B2(n9914), .ZN(n9901) );
  AOI22D1BWP30P140LVT U14432 ( .A1(i_data_bus[103]), .A2(n9915), .B1(
        i_data_bus[39]), .B2(n9916), .ZN(n9900) );
  ND2D1BWP30P140LVT U14433 ( .A1(n9901), .A2(n9900), .ZN(N3302) );
  AOI22D1BWP30P140LVT U14434 ( .A1(i_data_bus[6]), .A2(n6218), .B1(
        i_data_bus[102]), .B2(n9915), .ZN(n9903) );
  AOI22D1BWP30P140LVT U14435 ( .A1(i_data_bus[70]), .A2(n9914), .B1(
        i_data_bus[38]), .B2(n9916), .ZN(n9902) );
  ND2D1BWP30P140LVT U14436 ( .A1(n9903), .A2(n9902), .ZN(N3301) );
  AOI22D1BWP30P140LVT U14437 ( .A1(i_data_bus[3]), .A2(n6218), .B1(
        i_data_bus[67]), .B2(n9914), .ZN(n9905) );
  AOI22D1BWP30P140LVT U14438 ( .A1(i_data_bus[99]), .A2(n9915), .B1(
        i_data_bus[35]), .B2(n9916), .ZN(n9904) );
  ND2D1BWP30P140LVT U14439 ( .A1(n9905), .A2(n9904), .ZN(N3298) );
  AOI22D1BWP30P140LVT U14440 ( .A1(i_data_bus[8]), .A2(n6218), .B1(
        i_data_bus[72]), .B2(n9914), .ZN(n9907) );
  AOI22D1BWP30P140LVT U14441 ( .A1(i_data_bus[104]), .A2(n9915), .B1(
        i_data_bus[40]), .B2(n9916), .ZN(n9906) );
  ND2D1BWP30P140LVT U14442 ( .A1(n9907), .A2(n9906), .ZN(N3303) );
  AOI22D1BWP30P140LVT U14443 ( .A1(i_data_bus[19]), .A2(n6218), .B1(
        i_data_bus[115]), .B2(n9915), .ZN(n9909) );
  AOI22D1BWP30P140LVT U14444 ( .A1(i_data_bus[83]), .A2(n9914), .B1(
        i_data_bus[51]), .B2(n9916), .ZN(n9908) );
  ND2D1BWP30P140LVT U14445 ( .A1(n9909), .A2(n9908), .ZN(N3314) );
  AOI22D1BWP30P140LVT U14446 ( .A1(i_data_bus[15]), .A2(n6218), .B1(
        i_data_bus[79]), .B2(n9914), .ZN(n9911) );
  AOI22D1BWP30P140LVT U14447 ( .A1(i_data_bus[111]), .A2(n9915), .B1(
        i_data_bus[47]), .B2(n9916), .ZN(n9910) );
  ND2D1BWP30P140LVT U14448 ( .A1(n9911), .A2(n9910), .ZN(N3310) );
  AOI22D1BWP30P140LVT U14449 ( .A1(i_data_bus[108]), .A2(n9915), .B1(
        i_data_bus[12]), .B2(n6218), .ZN(n9913) );
  AOI22D1BWP30P140LVT U14450 ( .A1(i_data_bus[76]), .A2(n9914), .B1(
        i_data_bus[44]), .B2(n9916), .ZN(n9912) );
  ND2D1BWP30P140LVT U14451 ( .A1(n9913), .A2(n9912), .ZN(N3307) );
  AOI22D1BWP30P140LVT U14452 ( .A1(i_data_bus[122]), .A2(n9915), .B1(
        i_data_bus[90]), .B2(n9914), .ZN(n9918) );
  AOI22D1BWP30P140LVT U14453 ( .A1(i_data_bus[26]), .A2(n6218), .B1(
        i_data_bus[58]), .B2(n9916), .ZN(n9917) );
  ND2D1BWP30P140LVT U14454 ( .A1(n9918), .A2(n9917), .ZN(N3321) );
  AOI22D1BWP30P140LVT U14455 ( .A1(i_data_bus[606]), .A2(n9936), .B1(
        i_data_bus[638]), .B2(n9933), .ZN(n9920) );
  AOI22D1BWP30P140LVT U14456 ( .A1(i_data_bus[542]), .A2(n9934), .B1(
        i_data_bus[574]), .B2(n9935), .ZN(n9919) );
  ND2D1BWP30P140LVT U14457 ( .A1(n9920), .A2(n9919), .ZN(N5423) );
  AOI22D1BWP30P140LVT U14458 ( .A1(i_data_bus[534]), .A2(n9934), .B1(
        i_data_bus[598]), .B2(n9936), .ZN(n9922) );
  AOI22D1BWP30P140LVT U14459 ( .A1(i_data_bus[630]), .A2(n9933), .B1(
        i_data_bus[566]), .B2(n9935), .ZN(n9921) );
  ND2D1BWP30P140LVT U14460 ( .A1(n9922), .A2(n9921), .ZN(N5415) );
  AOI22D1BWP30P140LVT U14461 ( .A1(i_data_bus[628]), .A2(n9933), .B1(
        i_data_bus[596]), .B2(n9936), .ZN(n9924) );
  AOI22D1BWP30P140LVT U14462 ( .A1(i_data_bus[532]), .A2(n9934), .B1(
        i_data_bus[564]), .B2(n9935), .ZN(n9923) );
  ND2D1BWP30P140LVT U14463 ( .A1(n9924), .A2(n9923), .ZN(N5413) );
  AOI22D1BWP30P140LVT U14464 ( .A1(i_data_bus[526]), .A2(n9934), .B1(
        i_data_bus[622]), .B2(n9933), .ZN(n9926) );
  AOI22D1BWP30P140LVT U14465 ( .A1(i_data_bus[590]), .A2(n9936), .B1(
        i_data_bus[558]), .B2(n9935), .ZN(n9925) );
  ND2D1BWP30P140LVT U14466 ( .A1(n9926), .A2(n9925), .ZN(N5407) );
  AOI22D1BWP30P140LVT U14467 ( .A1(i_data_bus[621]), .A2(n9933), .B1(
        i_data_bus[589]), .B2(n9936), .ZN(n9928) );
  AOI22D1BWP30P140LVT U14468 ( .A1(i_data_bus[525]), .A2(n9934), .B1(
        i_data_bus[557]), .B2(n9935), .ZN(n9927) );
  ND2D1BWP30P140LVT U14469 ( .A1(n9928), .A2(n9927), .ZN(N5406) );
  AOI22D1BWP30P140LVT U14470 ( .A1(i_data_bus[586]), .A2(n9936), .B1(
        i_data_bus[522]), .B2(n9934), .ZN(n9930) );
  AOI22D1BWP30P140LVT U14471 ( .A1(i_data_bus[618]), .A2(n9933), .B1(
        i_data_bus[554]), .B2(n9935), .ZN(n9929) );
  ND2D1BWP30P140LVT U14472 ( .A1(n9930), .A2(n9929), .ZN(N5403) );
  AOI22D1BWP30P140LVT U14473 ( .A1(i_data_bus[517]), .A2(n9934), .B1(
        i_data_bus[581]), .B2(n9936), .ZN(n9932) );
  AOI22D1BWP30P140LVT U14474 ( .A1(i_data_bus[613]), .A2(n9933), .B1(
        i_data_bus[549]), .B2(n9935), .ZN(n9931) );
  ND2D1BWP30P140LVT U14475 ( .A1(n9932), .A2(n9931), .ZN(N5398) );
  AOI22D1BWP30P140LVT U14476 ( .A1(i_data_bus[512]), .A2(n9934), .B1(
        i_data_bus[608]), .B2(n9933), .ZN(n9938) );
  AOI22D1BWP30P140LVT U14477 ( .A1(i_data_bus[576]), .A2(n9936), .B1(
        i_data_bus[544]), .B2(n9935), .ZN(n9937) );
  ND2D1BWP30P140LVT U14478 ( .A1(n9938), .A2(n9937), .ZN(N5393) );
  AOI22D1BWP30P140LVT U14479 ( .A1(i_data_bus[31]), .A2(n10096), .B1(
        i_data_bus[63]), .B2(n10097), .ZN(n9940) );
  AOI22D1BWP30P140LVT U14480 ( .A1(i_data_bus[95]), .A2(n10095), .B1(
        i_data_bus[127]), .B2(n10098), .ZN(n9939) );
  ND2D1BWP30P140LVT U14481 ( .A1(n9940), .A2(n9939), .ZN(N6050) );
  AOI22D1BWP30P140LVT U14482 ( .A1(i_data_bus[48]), .A2(n10097), .B1(
        i_data_bus[80]), .B2(n10095), .ZN(n9942) );
  AOI22D1BWP30P140LVT U14483 ( .A1(i_data_bus[16]), .A2(n10096), .B1(
        i_data_bus[112]), .B2(n10098), .ZN(n9941) );
  ND2D1BWP30P140LVT U14484 ( .A1(n9942), .A2(n9941), .ZN(N6035) );
  AOI22D1BWP30P140LVT U14485 ( .A1(i_data_bus[73]), .A2(n10095), .B1(
        i_data_bus[9]), .B2(n10096), .ZN(n9944) );
  AOI22D1BWP30P140LVT U14486 ( .A1(i_data_bus[41]), .A2(n10097), .B1(
        i_data_bus[105]), .B2(n10098), .ZN(n9943) );
  ND2D1BWP30P140LVT U14487 ( .A1(n9944), .A2(n9943), .ZN(N6028) );
  AOI22D1BWP30P140LVT U14488 ( .A1(i_data_bus[43]), .A2(n10097), .B1(
        i_data_bus[75]), .B2(n10095), .ZN(n9946) );
  AOI22D1BWP30P140LVT U14489 ( .A1(i_data_bus[11]), .A2(n10096), .B1(
        i_data_bus[107]), .B2(n10098), .ZN(n9945) );
  ND2D1BWP30P140LVT U14490 ( .A1(n9946), .A2(n9945), .ZN(N6030) );
  AOI22D1BWP30P140LVT U14491 ( .A1(i_data_bus[4]), .A2(n10096), .B1(
        i_data_bus[68]), .B2(n10095), .ZN(n9948) );
  AOI22D1BWP30P140LVT U14492 ( .A1(i_data_bus[36]), .A2(n10097), .B1(
        i_data_bus[100]), .B2(n10098), .ZN(n9947) );
  ND2D1BWP30P140LVT U14493 ( .A1(n9948), .A2(n9947), .ZN(N6023) );
  AOI22D1BWP30P140LVT U14494 ( .A1(i_data_bus[60]), .A2(n10097), .B1(
        i_data_bus[28]), .B2(n10096), .ZN(n9950) );
  AOI22D1BWP30P140LVT U14495 ( .A1(i_data_bus[92]), .A2(n10095), .B1(
        i_data_bus[124]), .B2(n10098), .ZN(n9949) );
  ND2D1BWP30P140LVT U14496 ( .A1(n9950), .A2(n9949), .ZN(N6047) );
  AOI22D1BWP30P140LVT U14497 ( .A1(i_data_bus[24]), .A2(n10096), .B1(
        i_data_bus[88]), .B2(n10095), .ZN(n9952) );
  AOI22D1BWP30P140LVT U14498 ( .A1(i_data_bus[56]), .A2(n10097), .B1(
        i_data_bus[120]), .B2(n10098), .ZN(n9951) );
  ND2D1BWP30P140LVT U14499 ( .A1(n9952), .A2(n9951), .ZN(N6043) );
  AOI22D1BWP30P140LVT U14500 ( .A1(i_data_bus[69]), .A2(n10095), .B1(
        i_data_bus[37]), .B2(n10097), .ZN(n9954) );
  AOI22D1BWP30P140LVT U14501 ( .A1(i_data_bus[5]), .A2(n10096), .B1(
        i_data_bus[101]), .B2(n10098), .ZN(n9953) );
  ND2D1BWP30P140LVT U14502 ( .A1(n9954), .A2(n9953), .ZN(N6024) );
  AOI22D1BWP30P140LVT U14503 ( .A1(i_data_bus[90]), .A2(n10095), .B1(
        i_data_bus[58]), .B2(n10097), .ZN(n9956) );
  AOI22D1BWP30P140LVT U14504 ( .A1(i_data_bus[26]), .A2(n10096), .B1(
        i_data_bus[122]), .B2(n10098), .ZN(n9955) );
  ND2D1BWP30P140LVT U14505 ( .A1(n9956), .A2(n9955), .ZN(N6045) );
  AOI22D1BWP30P140LVT U14506 ( .A1(i_data_bus[17]), .A2(n10096), .B1(
        i_data_bus[49]), .B2(n10097), .ZN(n9958) );
  AOI22D1BWP30P140LVT U14507 ( .A1(i_data_bus[81]), .A2(n10095), .B1(
        i_data_bus[113]), .B2(n10098), .ZN(n9957) );
  ND2D1BWP30P140LVT U14508 ( .A1(n9958), .A2(n9957), .ZN(N6036) );
  AOI22D1BWP30P140LVT U14509 ( .A1(i_data_bus[7]), .A2(n10096), .B1(
        i_data_bus[39]), .B2(n10097), .ZN(n9960) );
  AOI22D1BWP30P140LVT U14510 ( .A1(i_data_bus[71]), .A2(n10095), .B1(
        i_data_bus[103]), .B2(n10098), .ZN(n9959) );
  ND2D1BWP30P140LVT U14511 ( .A1(n9960), .A2(n9959), .ZN(N6026) );
  AOI22D1BWP30P140LVT U14512 ( .A1(i_data_bus[87]), .A2(n10095), .B1(
        i_data_bus[23]), .B2(n10096), .ZN(n9962) );
  AOI22D1BWP30P140LVT U14513 ( .A1(i_data_bus[55]), .A2(n10097), .B1(
        i_data_bus[119]), .B2(n10098), .ZN(n9961) );
  ND2D1BWP30P140LVT U14514 ( .A1(n9962), .A2(n9961), .ZN(N6042) );
  AOI22D1BWP30P140LVT U14515 ( .A1(i_data_bus[13]), .A2(n10096), .B1(
        i_data_bus[45]), .B2(n10097), .ZN(n9964) );
  AOI22D1BWP30P140LVT U14516 ( .A1(i_data_bus[77]), .A2(n10095), .B1(
        i_data_bus[109]), .B2(n10098), .ZN(n9963) );
  ND2D1BWP30P140LVT U14517 ( .A1(n9964), .A2(n9963), .ZN(N6032) );
  AOI22D1BWP30P140LVT U14518 ( .A1(i_data_bus[72]), .A2(n9976), .B1(
        i_data_bus[40]), .B2(n9977), .ZN(n9966) );
  AOI22D1BWP30P140LVT U14519 ( .A1(i_data_bus[8]), .A2(n9969), .B1(
        i_data_bus[104]), .B2(n9978), .ZN(n9965) );
  ND2D1BWP30P140LVT U14520 ( .A1(n9966), .A2(n9965), .ZN(N2325) );
  AOI22D1BWP30P140LVT U14521 ( .A1(i_data_bus[20]), .A2(n9969), .B1(
        i_data_bus[52]), .B2(n9977), .ZN(n9968) );
  AOI22D1BWP30P140LVT U14522 ( .A1(i_data_bus[84]), .A2(n9976), .B1(
        i_data_bus[116]), .B2(n9978), .ZN(n9967) );
  ND2D1BWP30P140LVT U14523 ( .A1(n9968), .A2(n9967), .ZN(N2337) );
  AOI22D1BWP30P140LVT U14524 ( .A1(i_data_bus[11]), .A2(n9969), .B1(
        i_data_bus[75]), .B2(n9976), .ZN(n9971) );
  AOI22D1BWP30P140LVT U14525 ( .A1(i_data_bus[43]), .A2(n9977), .B1(
        i_data_bus[107]), .B2(n9978), .ZN(n9970) );
  ND2D1BWP30P140LVT U14526 ( .A1(n9971), .A2(n9970), .ZN(N2328) );
  AOI22D1BWP30P140LVT U14527 ( .A1(i_data_bus[55]), .A2(n9977), .B1(
        i_data_bus[23]), .B2(n9969), .ZN(n9973) );
  AOI22D1BWP30P140LVT U14528 ( .A1(i_data_bus[87]), .A2(n9976), .B1(
        i_data_bus[119]), .B2(n9978), .ZN(n9972) );
  ND2D1BWP30P140LVT U14529 ( .A1(n9973), .A2(n9972), .ZN(N2340) );
  AOI22D1BWP30P140LVT U14530 ( .A1(i_data_bus[78]), .A2(n9976), .B1(
        i_data_bus[46]), .B2(n9977), .ZN(n9975) );
  AOI22D1BWP30P140LVT U14531 ( .A1(i_data_bus[14]), .A2(n9969), .B1(
        i_data_bus[110]), .B2(n9978), .ZN(n9974) );
  ND2D1BWP30P140LVT U14532 ( .A1(n9975), .A2(n9974), .ZN(N2331) );
  AOI22D1BWP30P140LVT U14533 ( .A1(i_data_bus[60]), .A2(n9977), .B1(
        i_data_bus[92]), .B2(n9976), .ZN(n9980) );
  AOI22D1BWP30P140LVT U14534 ( .A1(i_data_bus[28]), .A2(n9969), .B1(
        i_data_bus[124]), .B2(n9978), .ZN(n9979) );
  ND2D1BWP30P140LVT U14535 ( .A1(n9980), .A2(n9979), .ZN(N2345) );
  AOI22D1BWP30P140LVT U14536 ( .A1(i_data_bus[606]), .A2(n10001), .B1(
        i_data_bus[638]), .B2(n10003), .ZN(n9982) );
  AOI22D1BWP30P140LVT U14537 ( .A1(i_data_bus[542]), .A2(n6222), .B1(
        i_data_bus[574]), .B2(n10002), .ZN(n9981) );
  ND2D1BWP30P140LVT U14538 ( .A1(n9982), .A2(n9981), .ZN(N4189) );
  AOI22D1BWP30P140LVT U14539 ( .A1(i_data_bus[534]), .A2(n10006), .B1(
        i_data_bus[598]), .B2(n10013), .ZN(n9984) );
  AOI22D1BWP30P140LVT U14540 ( .A1(i_data_bus[630]), .A2(n10011), .B1(
        i_data_bus[566]), .B2(n10012), .ZN(n9983) );
  ND2D1BWP30P140LVT U14541 ( .A1(n9984), .A2(n9983), .ZN(N2691) );
  AOI22D1BWP30P140LVT U14542 ( .A1(i_data_bus[630]), .A2(n10003), .B1(
        i_data_bus[598]), .B2(n10001), .ZN(n9986) );
  AOI22D1BWP30P140LVT U14543 ( .A1(i_data_bus[534]), .A2(n6222), .B1(
        i_data_bus[566]), .B2(n10002), .ZN(n9985) );
  ND2D1BWP30P140LVT U14544 ( .A1(n9986), .A2(n9985), .ZN(N4181) );
  AOI22D1BWP30P140LVT U14545 ( .A1(i_data_bus[629]), .A2(n10003), .B1(
        i_data_bus[597]), .B2(n10001), .ZN(n9988) );
  AOI22D1BWP30P140LVT U14546 ( .A1(i_data_bus[533]), .A2(n6222), .B1(
        i_data_bus[565]), .B2(n10002), .ZN(n9987) );
  ND2D1BWP30P140LVT U14547 ( .A1(n9988), .A2(n9987), .ZN(N4180) );
  AOI22D1BWP30P140LVT U14548 ( .A1(i_data_bus[584]), .A2(n10013), .B1(
        i_data_bus[616]), .B2(n10011), .ZN(n9990) );
  AOI22D1BWP30P140LVT U14549 ( .A1(i_data_bus[520]), .A2(n10006), .B1(
        i_data_bus[552]), .B2(n10012), .ZN(n9989) );
  ND2D1BWP30P140LVT U14550 ( .A1(n9990), .A2(n9989), .ZN(N2677) );
  AOI22D1BWP30P140LVT U14551 ( .A1(i_data_bus[525]), .A2(n6222), .B1(
        i_data_bus[589]), .B2(n10001), .ZN(n9992) );
  AOI22D1BWP30P140LVT U14552 ( .A1(i_data_bus[621]), .A2(n10003), .B1(
        i_data_bus[557]), .B2(n10002), .ZN(n9991) );
  ND2D1BWP30P140LVT U14553 ( .A1(n9992), .A2(n9991), .ZN(N4172) );
  AOI22D1BWP30P140LVT U14554 ( .A1(i_data_bus[634]), .A2(n10011), .B1(
        i_data_bus[602]), .B2(n10013), .ZN(n9994) );
  AOI22D1BWP30P140LVT U14555 ( .A1(i_data_bus[538]), .A2(n10006), .B1(
        i_data_bus[570]), .B2(n10012), .ZN(n9993) );
  ND2D1BWP30P140LVT U14556 ( .A1(n9994), .A2(n9993), .ZN(N2695) );
  AOI22D1BWP30P140LVT U14557 ( .A1(i_data_bus[619]), .A2(n10011), .B1(
        i_data_bus[523]), .B2(n10006), .ZN(n9996) );
  AOI22D1BWP30P140LVT U14558 ( .A1(i_data_bus[587]), .A2(n10013), .B1(
        i_data_bus[555]), .B2(n10012), .ZN(n9995) );
  ND2D1BWP30P140LVT U14559 ( .A1(n9996), .A2(n9995), .ZN(N2680) );
  AOI22D1BWP30P140LVT U14560 ( .A1(i_data_bus[517]), .A2(n6222), .B1(
        i_data_bus[581]), .B2(n10001), .ZN(n9998) );
  AOI22D1BWP30P140LVT U14561 ( .A1(i_data_bus[613]), .A2(n10003), .B1(
        i_data_bus[549]), .B2(n10002), .ZN(n9997) );
  ND2D1BWP30P140LVT U14562 ( .A1(n9998), .A2(n9997), .ZN(N4164) );
  AOI22D1BWP30P140LVT U14563 ( .A1(i_data_bus[578]), .A2(n10001), .B1(
        i_data_bus[514]), .B2(n6222), .ZN(n10000) );
  AOI22D1BWP30P140LVT U14564 ( .A1(i_data_bus[610]), .A2(n10003), .B1(
        i_data_bus[546]), .B2(n10002), .ZN(n9999) );
  ND2D1BWP30P140LVT U14565 ( .A1(n10000), .A2(n9999), .ZN(N4161) );
  AOI22D1BWP30P140LVT U14566 ( .A1(i_data_bus[541]), .A2(n6222), .B1(
        i_data_bus[605]), .B2(n10001), .ZN(n10005) );
  AOI22D1BWP30P140LVT U14567 ( .A1(i_data_bus[637]), .A2(n10003), .B1(
        i_data_bus[573]), .B2(n10002), .ZN(n10004) );
  ND2D1BWP30P140LVT U14568 ( .A1(n10005), .A2(n10004), .ZN(N4188) );
  AOI22D1BWP30P140LVT U14569 ( .A1(i_data_bus[512]), .A2(n10006), .B1(
        i_data_bus[576]), .B2(n10013), .ZN(n10008) );
  AOI22D1BWP30P140LVT U14570 ( .A1(i_data_bus[608]), .A2(n10011), .B1(
        i_data_bus[544]), .B2(n10012), .ZN(n10007) );
  ND2D1BWP30P140LVT U14571 ( .A1(n10008), .A2(n10007), .ZN(N2669) );
  AOI22D1BWP30P140LVT U14572 ( .A1(i_data_bus[606]), .A2(n10013), .B1(
        i_data_bus[542]), .B2(n10006), .ZN(n10010) );
  AOI22D1BWP30P140LVT U14573 ( .A1(i_data_bus[638]), .A2(n10011), .B1(
        i_data_bus[574]), .B2(n10012), .ZN(n10009) );
  ND2D1BWP30P140LVT U14574 ( .A1(n10010), .A2(n10009), .ZN(N2699) );
  AOI22D1BWP30P140LVT U14575 ( .A1(i_data_bus[533]), .A2(n10006), .B1(
        i_data_bus[629]), .B2(n10011), .ZN(n10015) );
  AOI22D1BWP30P140LVT U14576 ( .A1(i_data_bus[597]), .A2(n10013), .B1(
        i_data_bus[565]), .B2(n10012), .ZN(n10014) );
  ND2D1BWP30P140LVT U14577 ( .A1(n10015), .A2(n10014), .ZN(N2690) );
  AOI22D1BWP30P140LVT U14578 ( .A1(i_data_bus[249]), .A2(n10035), .B1(
        i_data_bus[217]), .B2(n10033), .ZN(n10017) );
  AOI22D1BWP30P140LVT U14579 ( .A1(i_data_bus[153]), .A2(n10026), .B1(
        i_data_bus[185]), .B2(n10034), .ZN(n10016) );
  ND2D1BWP30P140LVT U14580 ( .A1(n10017), .A2(n10016), .ZN(N3536) );
  AOI22D1BWP30P140LVT U14581 ( .A1(i_data_bus[245]), .A2(n10035), .B1(
        i_data_bus[149]), .B2(n10026), .ZN(n10019) );
  AOI22D1BWP30P140LVT U14582 ( .A1(i_data_bus[213]), .A2(n10033), .B1(
        i_data_bus[181]), .B2(n10034), .ZN(n10018) );
  ND2D1BWP30P140LVT U14583 ( .A1(n10019), .A2(n10018), .ZN(N3532) );
  AOI22D1BWP30P140LVT U14584 ( .A1(i_data_bus[235]), .A2(n10035), .B1(
        i_data_bus[203]), .B2(n10033), .ZN(n10021) );
  AOI22D1BWP30P140LVT U14585 ( .A1(i_data_bus[139]), .A2(n10026), .B1(
        i_data_bus[171]), .B2(n10034), .ZN(n10020) );
  ND2D1BWP30P140LVT U14586 ( .A1(n10021), .A2(n10020), .ZN(N3522) );
  AOI22D1BWP30P140LVT U14587 ( .A1(i_data_bus[232]), .A2(n10035), .B1(
        i_data_bus[200]), .B2(n10033), .ZN(n10023) );
  AOI22D1BWP30P140LVT U14588 ( .A1(i_data_bus[136]), .A2(n10026), .B1(
        i_data_bus[168]), .B2(n10034), .ZN(n10022) );
  ND2D1BWP30P140LVT U14589 ( .A1(n10023), .A2(n10022), .ZN(N3519) );
  AOI22D1BWP30P140LVT U14590 ( .A1(i_data_bus[231]), .A2(n10038), .B1(
        i_data_bus[135]), .B2(n9318), .ZN(n10025) );
  AOI22D1BWP30P140LVT U14591 ( .A1(i_data_bus[199]), .A2(n10039), .B1(
        i_data_bus[167]), .B2(n10040), .ZN(n10024) );
  ND2D1BWP30P140LVT U14592 ( .A1(n10025), .A2(n10024), .ZN(N8966) );
  AOI22D1BWP30P140LVT U14593 ( .A1(i_data_bus[128]), .A2(n10026), .B1(
        i_data_bus[192]), .B2(n10033), .ZN(n10028) );
  AOI22D1BWP30P140LVT U14594 ( .A1(i_data_bus[224]), .A2(n10035), .B1(
        i_data_bus[160]), .B2(n10034), .ZN(n10027) );
  ND2D1BWP30P140LVT U14595 ( .A1(n10028), .A2(n10027), .ZN(N3511) );
  AOI22D1BWP30P140LVT U14596 ( .A1(i_data_bus[213]), .A2(n10039), .B1(
        i_data_bus[149]), .B2(n9318), .ZN(n10030) );
  AOI22D1BWP30P140LVT U14597 ( .A1(i_data_bus[245]), .A2(n10038), .B1(
        i_data_bus[181]), .B2(n10040), .ZN(n10029) );
  ND2D1BWP30P140LVT U14598 ( .A1(n10030), .A2(n10029), .ZN(N8980) );
  AOI22D1BWP30P140LVT U14599 ( .A1(i_data_bus[138]), .A2(n9318), .B1(
        i_data_bus[202]), .B2(n10039), .ZN(n10032) );
  AOI22D1BWP30P140LVT U14600 ( .A1(i_data_bus[234]), .A2(n10038), .B1(
        i_data_bus[170]), .B2(n10040), .ZN(n10031) );
  ND2D1BWP30P140LVT U14601 ( .A1(n10032), .A2(n10031), .ZN(N8969) );
  AOI22D1BWP30P140LVT U14602 ( .A1(i_data_bus[131]), .A2(n10026), .B1(
        i_data_bus[195]), .B2(n10033), .ZN(n10037) );
  AOI22D1BWP30P140LVT U14603 ( .A1(i_data_bus[227]), .A2(n10035), .B1(
        i_data_bus[163]), .B2(n10034), .ZN(n10036) );
  ND2D1BWP30P140LVT U14604 ( .A1(n10037), .A2(n10036), .ZN(N3514) );
  AOI22D1BWP30P140LVT U14605 ( .A1(i_data_bus[215]), .A2(n10039), .B1(
        i_data_bus[247]), .B2(n10038), .ZN(n10042) );
  AOI22D1BWP30P140LVT U14606 ( .A1(i_data_bus[151]), .A2(n9318), .B1(
        i_data_bus[183]), .B2(n10040), .ZN(n10041) );
  ND2D1BWP30P140LVT U14607 ( .A1(n10042), .A2(n10041), .ZN(N8982) );
  AOI22D1BWP30P140LVT U14608 ( .A1(i_data_bus[375]), .A2(n10051), .B1(
        i_data_bus[343]), .B2(n10054), .ZN(n10044) );
  AOI22D1BWP30P140LVT U14609 ( .A1(i_data_bus[279]), .A2(n10052), .B1(
        i_data_bus[311]), .B2(n10053), .ZN(n10043) );
  ND2D1BWP30P140LVT U14610 ( .A1(n10044), .A2(n10043), .ZN(N6474) );
  AOI22D1BWP30P140LVT U14611 ( .A1(i_data_bus[355]), .A2(n10051), .B1(
        i_data_bus[323]), .B2(n10054), .ZN(n10046) );
  AOI22D1BWP30P140LVT U14612 ( .A1(i_data_bus[259]), .A2(n10052), .B1(
        i_data_bus[291]), .B2(n10053), .ZN(n10045) );
  ND2D1BWP30P140LVT U14613 ( .A1(n10046), .A2(n10045), .ZN(N6454) );
  AOI22D1BWP30P140LVT U14614 ( .A1(i_data_bus[268]), .A2(n10052), .B1(
        i_data_bus[332]), .B2(n10054), .ZN(n10048) );
  AOI22D1BWP30P140LVT U14615 ( .A1(i_data_bus[364]), .A2(n10051), .B1(
        i_data_bus[300]), .B2(n10053), .ZN(n10047) );
  ND2D1BWP30P140LVT U14616 ( .A1(n10048), .A2(n10047), .ZN(N6463) );
  AOI22D1BWP30P140LVT U14617 ( .A1(i_data_bus[360]), .A2(n10051), .B1(
        i_data_bus[264]), .B2(n10052), .ZN(n10050) );
  AOI22D1BWP30P140LVT U14618 ( .A1(i_data_bus[328]), .A2(n10054), .B1(
        i_data_bus[296]), .B2(n10053), .ZN(n10049) );
  ND2D1BWP30P140LVT U14619 ( .A1(n10050), .A2(n10049), .ZN(N6459) );
  AOI22D1BWP30P140LVT U14620 ( .A1(i_data_bus[275]), .A2(n10052), .B1(
        i_data_bus[371]), .B2(n10051), .ZN(n10056) );
  AOI22D1BWP30P140LVT U14621 ( .A1(i_data_bus[339]), .A2(n10054), .B1(
        i_data_bus[307]), .B2(n10053), .ZN(n10055) );
  ND2D1BWP30P140LVT U14622 ( .A1(n10056), .A2(n10055), .ZN(N6470) );
  AOI22D1BWP30P140LVT U14623 ( .A1(i_data_bus[25]), .A2(n10096), .B1(
        i_data_bus[89]), .B2(n10095), .ZN(n10058) );
  AOI22D1BWP30P140LVT U14624 ( .A1(i_data_bus[121]), .A2(n10098), .B1(
        i_data_bus[57]), .B2(n10097), .ZN(n10057) );
  ND2D1BWP30P140LVT U14625 ( .A1(n10058), .A2(n10057), .ZN(N6044) );
  AOI22D1BWP30P140LVT U14626 ( .A1(i_data_bus[76]), .A2(n10086), .B1(
        i_data_bus[108]), .B2(n10085), .ZN(n10060) );
  AOI22D1BWP30P140LVT U14627 ( .A1(i_data_bus[12]), .A2(n10088), .B1(
        i_data_bus[44]), .B2(n10087), .ZN(n10059) );
  ND2D1BWP30P140LVT U14628 ( .A1(n10060), .A2(n10059), .ZN(N5053) );
  AOI22D1BWP30P140LVT U14629 ( .A1(i_data_bus[101]), .A2(n10085), .B1(
        i_data_bus[69]), .B2(n10086), .ZN(n10062) );
  AOI22D1BWP30P140LVT U14630 ( .A1(i_data_bus[5]), .A2(n10088), .B1(
        i_data_bus[37]), .B2(n10087), .ZN(n10061) );
  ND2D1BWP30P140LVT U14631 ( .A1(n10062), .A2(n10061), .ZN(N5046) );
  AOI22D1BWP30P140LVT U14632 ( .A1(i_data_bus[15]), .A2(n10088), .B1(
        i_data_bus[79]), .B2(n10086), .ZN(n10064) );
  AOI22D1BWP30P140LVT U14633 ( .A1(i_data_bus[111]), .A2(n10085), .B1(
        i_data_bus[47]), .B2(n10087), .ZN(n10063) );
  ND2D1BWP30P140LVT U14634 ( .A1(n10064), .A2(n10063), .ZN(N5056) );
  AOI22D1BWP30P140LVT U14635 ( .A1(i_data_bus[125]), .A2(n10098), .B1(
        i_data_bus[29]), .B2(n10096), .ZN(n10066) );
  AOI22D1BWP30P140LVT U14636 ( .A1(i_data_bus[93]), .A2(n10095), .B1(
        i_data_bus[61]), .B2(n10097), .ZN(n10065) );
  ND2D1BWP30P140LVT U14637 ( .A1(n10066), .A2(n10065), .ZN(N6048) );
  AOI22D1BWP30P140LVT U14638 ( .A1(i_data_bus[102]), .A2(n10098), .B1(
        i_data_bus[70]), .B2(n10095), .ZN(n10068) );
  AOI22D1BWP30P140LVT U14639 ( .A1(i_data_bus[6]), .A2(n10096), .B1(
        i_data_bus[38]), .B2(n10097), .ZN(n10067) );
  ND2D1BWP30P140LVT U14640 ( .A1(n10068), .A2(n10067), .ZN(N6025) );
  AOI22D1BWP30P140LVT U14641 ( .A1(i_data_bus[14]), .A2(n10088), .B1(
        i_data_bus[110]), .B2(n10085), .ZN(n10070) );
  AOI22D1BWP30P140LVT U14642 ( .A1(i_data_bus[78]), .A2(n10086), .B1(
        i_data_bus[46]), .B2(n10087), .ZN(n10069) );
  ND2D1BWP30P140LVT U14643 ( .A1(n10070), .A2(n10069), .ZN(N5055) );
  AOI22D1BWP30P140LVT U14644 ( .A1(i_data_bus[81]), .A2(n10086), .B1(
        i_data_bus[113]), .B2(n10085), .ZN(n10072) );
  AOI22D1BWP30P140LVT U14645 ( .A1(i_data_bus[17]), .A2(n10088), .B1(
        i_data_bus[49]), .B2(n10087), .ZN(n10071) );
  ND2D1BWP30P140LVT U14646 ( .A1(n10072), .A2(n10071), .ZN(N5058) );
  AOI22D1BWP30P140LVT U14647 ( .A1(i_data_bus[84]), .A2(n10095), .B1(
        i_data_bus[116]), .B2(n10098), .ZN(n10074) );
  AOI22D1BWP30P140LVT U14648 ( .A1(i_data_bus[20]), .A2(n10096), .B1(
        i_data_bus[52]), .B2(n10097), .ZN(n10073) );
  ND2D1BWP30P140LVT U14649 ( .A1(n10074), .A2(n10073), .ZN(N6039) );
  AOI22D1BWP30P140LVT U14650 ( .A1(i_data_bus[19]), .A2(n10088), .B1(
        i_data_bus[115]), .B2(n10085), .ZN(n10076) );
  AOI22D1BWP30P140LVT U14651 ( .A1(i_data_bus[83]), .A2(n10086), .B1(
        i_data_bus[51]), .B2(n10087), .ZN(n10075) );
  ND2D1BWP30P140LVT U14652 ( .A1(n10076), .A2(n10075), .ZN(N5060) );
  AOI22D1BWP30P140LVT U14653 ( .A1(i_data_bus[97]), .A2(n10085), .B1(
        i_data_bus[65]), .B2(n10086), .ZN(n10078) );
  AOI22D1BWP30P140LVT U14654 ( .A1(i_data_bus[1]), .A2(n10088), .B1(
        i_data_bus[33]), .B2(n10087), .ZN(n10077) );
  ND2D1BWP30P140LVT U14655 ( .A1(n10078), .A2(n10077), .ZN(N5042) );
  AOI22D1BWP30P140LVT U14656 ( .A1(i_data_bus[26]), .A2(n10088), .B1(
        i_data_bus[90]), .B2(n10086), .ZN(n10080) );
  AOI22D1BWP30P140LVT U14657 ( .A1(i_data_bus[122]), .A2(n10085), .B1(
        i_data_bus[58]), .B2(n10087), .ZN(n10079) );
  ND2D1BWP30P140LVT U14658 ( .A1(n10080), .A2(n10079), .ZN(N5067) );
  AOI22D1BWP30P140LVT U14659 ( .A1(i_data_bus[88]), .A2(n10086), .B1(
        i_data_bus[120]), .B2(n10085), .ZN(n10082) );
  AOI22D1BWP30P140LVT U14660 ( .A1(i_data_bus[24]), .A2(n10088), .B1(
        i_data_bus[56]), .B2(n10087), .ZN(n10081) );
  ND2D1BWP30P140LVT U14661 ( .A1(n10082), .A2(n10081), .ZN(N5065) );
  AOI22D1BWP30P140LVT U14662 ( .A1(i_data_bus[8]), .A2(n10088), .B1(
        i_data_bus[72]), .B2(n10086), .ZN(n10084) );
  AOI22D1BWP30P140LVT U14663 ( .A1(i_data_bus[104]), .A2(n10085), .B1(
        i_data_bus[40]), .B2(n10087), .ZN(n10083) );
  ND2D1BWP30P140LVT U14664 ( .A1(n10084), .A2(n10083), .ZN(N5049) );
  AOI22D1BWP30P140LVT U14665 ( .A1(i_data_bus[64]), .A2(n10086), .B1(
        i_data_bus[96]), .B2(n10085), .ZN(n10090) );
  AOI22D1BWP30P140LVT U14666 ( .A1(i_data_bus[0]), .A2(n10088), .B1(
        i_data_bus[32]), .B2(n10087), .ZN(n10089) );
  ND2D1BWP30P140LVT U14667 ( .A1(n10090), .A2(n10089), .ZN(N5041) );
  AOI22D1BWP30P140LVT U14668 ( .A1(i_data_bus[123]), .A2(n10098), .B1(
        i_data_bus[91]), .B2(n10095), .ZN(n10092) );
  AOI22D1BWP30P140LVT U14669 ( .A1(i_data_bus[27]), .A2(n10096), .B1(
        i_data_bus[59]), .B2(n10097), .ZN(n10091) );
  ND2D1BWP30P140LVT U14670 ( .A1(n10092), .A2(n10091), .ZN(N6046) );
  AOI22D1BWP30P140LVT U14671 ( .A1(i_data_bus[14]), .A2(n10096), .B1(
        i_data_bus[78]), .B2(n10095), .ZN(n10094) );
  AOI22D1BWP30P140LVT U14672 ( .A1(i_data_bus[110]), .A2(n10098), .B1(
        i_data_bus[46]), .B2(n10097), .ZN(n10093) );
  ND2D1BWP30P140LVT U14673 ( .A1(n10094), .A2(n10093), .ZN(N6033) );
  AOI22D1BWP30P140LVT U14674 ( .A1(i_data_bus[15]), .A2(n10096), .B1(
        i_data_bus[79]), .B2(n10095), .ZN(n10100) );
  AOI22D1BWP30P140LVT U14675 ( .A1(i_data_bus[111]), .A2(n10098), .B1(
        i_data_bus[47]), .B2(n10097), .ZN(n10099) );
  ND2D1BWP30P140LVT U14676 ( .A1(n10100), .A2(n10099), .ZN(N6034) );
  AOI22D1BWP30P140LVT U14677 ( .A1(i_data_bus[41]), .A2(n10118), .B1(
        i_data_bus[9]), .B2(n10116), .ZN(n10102) );
  AOI22D1BWP30P140LVT U14678 ( .A1(i_data_bus[73]), .A2(n10115), .B1(
        i_data_bus[105]), .B2(n10117), .ZN(n10101) );
  ND2D1BWP30P140LVT U14679 ( .A1(n10102), .A2(n10101), .ZN(N7774) );
  AOI22D1BWP30P140LVT U14680 ( .A1(i_data_bus[72]), .A2(n10115), .B1(
        i_data_bus[40]), .B2(n10118), .ZN(n10104) );
  AOI22D1BWP30P140LVT U14681 ( .A1(i_data_bus[8]), .A2(n10116), .B1(
        i_data_bus[104]), .B2(n10117), .ZN(n10103) );
  ND2D1BWP30P140LVT U14682 ( .A1(n10104), .A2(n10103), .ZN(N7773) );
  AOI22D1BWP30P140LVT U14683 ( .A1(i_data_bus[32]), .A2(n10118), .B1(
        i_data_bus[64]), .B2(n10115), .ZN(n10106) );
  AOI22D1BWP30P140LVT U14684 ( .A1(i_data_bus[0]), .A2(n10116), .B1(
        i_data_bus[96]), .B2(n10117), .ZN(n10105) );
  ND2D1BWP30P140LVT U14685 ( .A1(n10106), .A2(n10105), .ZN(N7765) );
  AOI22D1BWP30P140LVT U14686 ( .A1(i_data_bus[19]), .A2(n10116), .B1(
        i_data_bus[83]), .B2(n10115), .ZN(n10108) );
  AOI22D1BWP30P140LVT U14687 ( .A1(i_data_bus[51]), .A2(n10118), .B1(
        i_data_bus[115]), .B2(n10117), .ZN(n10107) );
  ND2D1BWP30P140LVT U14688 ( .A1(n10108), .A2(n10107), .ZN(N7784) );
  AOI22D1BWP30P140LVT U14689 ( .A1(i_data_bus[78]), .A2(n10115), .B1(
        i_data_bus[46]), .B2(n10118), .ZN(n10110) );
  AOI22D1BWP30P140LVT U14690 ( .A1(i_data_bus[14]), .A2(n10116), .B1(
        i_data_bus[110]), .B2(n10117), .ZN(n10109) );
  ND2D1BWP30P140LVT U14691 ( .A1(n10110), .A2(n10109), .ZN(N7779) );
  AOI22D1BWP30P140LVT U14692 ( .A1(i_data_bus[50]), .A2(n10118), .B1(
        i_data_bus[82]), .B2(n10115), .ZN(n10112) );
  AOI22D1BWP30P140LVT U14693 ( .A1(i_data_bus[18]), .A2(n10116), .B1(
        i_data_bus[114]), .B2(n10117), .ZN(n10111) );
  ND2D1BWP30P140LVT U14694 ( .A1(n10112), .A2(n10111), .ZN(N7783) );
  AOI22D1BWP30P140LVT U14695 ( .A1(i_data_bus[90]), .A2(n10115), .B1(
        i_data_bus[58]), .B2(n10118), .ZN(n10114) );
  AOI22D1BWP30P140LVT U14696 ( .A1(i_data_bus[26]), .A2(n10116), .B1(
        i_data_bus[122]), .B2(n10117), .ZN(n10113) );
  ND2D1BWP30P140LVT U14697 ( .A1(n10114), .A2(n10113), .ZN(N7791) );
  AOI22D1BWP30P140LVT U14698 ( .A1(i_data_bus[30]), .A2(n10116), .B1(
        i_data_bus[94]), .B2(n10115), .ZN(n10120) );
  AOI22D1BWP30P140LVT U14699 ( .A1(i_data_bus[62]), .A2(n10118), .B1(
        i_data_bus[126]), .B2(n10117), .ZN(n10119) );
  ND2D1BWP30P140LVT U14700 ( .A1(n10120), .A2(n10119), .ZN(N7795) );
  AOI22D1BWP30P140LVT U14701 ( .A1(i_data_bus[213]), .A2(n10132), .B1(
        i_data_bus[245]), .B2(n10131), .ZN(n10122) );
  AOI22D1BWP30P140LVT U14702 ( .A1(i_data_bus[149]), .A2(n10134), .B1(
        i_data_bus[181]), .B2(n10133), .ZN(n10121) );
  ND2D1BWP30P140LVT U14703 ( .A1(n10122), .A2(n10121), .ZN(N7874) );
  AOI22D1BWP30P140LVT U14704 ( .A1(i_data_bus[206]), .A2(n10132), .B1(
        i_data_bus[238]), .B2(n10131), .ZN(n10124) );
  AOI22D1BWP30P140LVT U14705 ( .A1(i_data_bus[142]), .A2(n10134), .B1(
        i_data_bus[174]), .B2(n10133), .ZN(n10123) );
  ND2D1BWP30P140LVT U14706 ( .A1(n10124), .A2(n10123), .ZN(N7867) );
  AOI22D1BWP30P140LVT U14707 ( .A1(i_data_bus[138]), .A2(n10134), .B1(
        i_data_bus[202]), .B2(n10132), .ZN(n10126) );
  AOI22D1BWP30P140LVT U14708 ( .A1(i_data_bus[234]), .A2(n10131), .B1(
        i_data_bus[170]), .B2(n10133), .ZN(n10125) );
  ND2D1BWP30P140LVT U14709 ( .A1(n10126), .A2(n10125), .ZN(N7863) );
  AOI22D1BWP30P140LVT U14710 ( .A1(i_data_bus[136]), .A2(n10134), .B1(
        i_data_bus[200]), .B2(n10132), .ZN(n10128) );
  AOI22D1BWP30P140LVT U14711 ( .A1(i_data_bus[232]), .A2(n10131), .B1(
        i_data_bus[168]), .B2(n10133), .ZN(n10127) );
  ND2D1BWP30P140LVT U14712 ( .A1(n10128), .A2(n10127), .ZN(N7861) );
  AOI22D1BWP30P140LVT U14713 ( .A1(i_data_bus[231]), .A2(n10131), .B1(
        i_data_bus[135]), .B2(n10134), .ZN(n10130) );
  AOI22D1BWP30P140LVT U14714 ( .A1(i_data_bus[199]), .A2(n10132), .B1(
        i_data_bus[167]), .B2(n10133), .ZN(n10129) );
  ND2D1BWP30P140LVT U14715 ( .A1(n10130), .A2(n10129), .ZN(N7860) );
  AOI22D1BWP30P140LVT U14716 ( .A1(i_data_bus[218]), .A2(n10132), .B1(
        i_data_bus[250]), .B2(n10131), .ZN(n10136) );
  AOI22D1BWP30P140LVT U14717 ( .A1(i_data_bus[154]), .A2(n10134), .B1(
        i_data_bus[186]), .B2(n10133), .ZN(n10135) );
  ND2D1BWP30P140LVT U14718 ( .A1(n10136), .A2(n10135), .ZN(N7879) );
  NR4D1BWP30P140LVT U14719 ( .A1(i_cmd[56]), .A2(n11180), .A3(n10137), .A4(
        n10664), .ZN(n10368) );
  INR4D1BWP30P140LVT U14720 ( .A1(i_cmd[48]), .B1(i_cmd[32]), .B2(n11177), 
        .B3(n10667), .ZN(n10367) );
  AOI22D1BWP30P140LVT U14721 ( .A1(n10368), .A2(i_data_bus[163]), .B1(n10367), 
        .B2(i_data_bus[195]), .ZN(n10139) );
  NR4D1BWP30P140LVT U14722 ( .A1(i_cmd[40]), .A2(n10670), .A3(n11179), .A4(
        n10137), .ZN(n10369) );
  NR3D0P7BWP30P140LVT U14723 ( .A1(i_cmd[40]), .A2(i_cmd[56]), .A3(i_cmd[48]), 
        .ZN(n11176) );
  AOI22D1BWP30P140LVT U14724 ( .A1(n10369), .A2(i_data_bus[227]), .B1(n10360), 
        .B2(i_data_bus[131]), .ZN(n10138) );
  ND2D1BWP30P140LVT U14725 ( .A1(n10139), .A2(n10138), .ZN(N766) );
  AOI22D1BWP30P140LVT U14726 ( .A1(n10368), .A2(i_data_bus[189]), .B1(n10367), 
        .B2(i_data_bus[221]), .ZN(n10141) );
  AOI22D1BWP30P140LVT U14727 ( .A1(n10369), .A2(i_data_bus[253]), .B1(n10360), 
        .B2(i_data_bus[157]), .ZN(n10140) );
  ND2D1BWP30P140LVT U14728 ( .A1(n10141), .A2(n10140), .ZN(N792) );
  AOI22D1BWP30P140LVT U14729 ( .A1(n10368), .A2(i_data_bus[170]), .B1(n10367), 
        .B2(i_data_bus[202]), .ZN(n10143) );
  AOI22D1BWP30P140LVT U14730 ( .A1(n10369), .A2(i_data_bus[234]), .B1(n10360), 
        .B2(i_data_bus[138]), .ZN(n10142) );
  ND2D1BWP30P140LVT U14731 ( .A1(n10143), .A2(n10142), .ZN(N773) );
  AOI22D1BWP30P140LVT U14732 ( .A1(n10368), .A2(i_data_bus[168]), .B1(n10367), 
        .B2(i_data_bus[200]), .ZN(n10145) );
  AOI22D1BWP30P140LVT U14733 ( .A1(n10369), .A2(i_data_bus[232]), .B1(n10360), 
        .B2(i_data_bus[136]), .ZN(n10144) );
  ND2D1BWP30P140LVT U14734 ( .A1(n10145), .A2(n10144), .ZN(N771) );
  AOI22D1BWP30P140LVT U14735 ( .A1(n10369), .A2(i_data_bus[235]), .B1(n10367), 
        .B2(i_data_bus[203]), .ZN(n10147) );
  AOI22D1BWP30P140LVT U14736 ( .A1(n10368), .A2(i_data_bus[171]), .B1(n10360), 
        .B2(i_data_bus[139]), .ZN(n10146) );
  ND2D1BWP30P140LVT U14737 ( .A1(n10147), .A2(n10146), .ZN(N774) );
  AOI22D1BWP30P140LVT U14738 ( .A1(n10369), .A2(i_data_bus[236]), .B1(n10367), 
        .B2(i_data_bus[204]), .ZN(n10149) );
  AOI22D1BWP30P140LVT U14739 ( .A1(n10368), .A2(i_data_bus[172]), .B1(n10360), 
        .B2(i_data_bus[140]), .ZN(n10148) );
  ND2D1BWP30P140LVT U14740 ( .A1(n10149), .A2(n10148), .ZN(N775) );
  AOI22D1BWP30P140LVT U14741 ( .A1(n10369), .A2(i_data_bus[240]), .B1(n10367), 
        .B2(i_data_bus[208]), .ZN(n10151) );
  AOI22D1BWP30P140LVT U14742 ( .A1(n10368), .A2(i_data_bus[176]), .B1(n10360), 
        .B2(i_data_bus[144]), .ZN(n10150) );
  ND2D1BWP30P140LVT U14743 ( .A1(n10151), .A2(n10150), .ZN(N779) );
  AOI22D1BWP30P140LVT U14744 ( .A1(n10369), .A2(i_data_bus[239]), .B1(n10367), 
        .B2(i_data_bus[207]), .ZN(n10153) );
  AOI22D1BWP30P140LVT U14745 ( .A1(n10368), .A2(i_data_bus[175]), .B1(n10360), 
        .B2(i_data_bus[143]), .ZN(n10152) );
  ND2D1BWP30P140LVT U14746 ( .A1(n10153), .A2(n10152), .ZN(N778) );
  AOI22D1BWP30P140LVT U14747 ( .A1(n10369), .A2(i_data_bus[251]), .B1(n10367), 
        .B2(i_data_bus[219]), .ZN(n10155) );
  AOI22D1BWP30P140LVT U14748 ( .A1(n10368), .A2(i_data_bus[187]), .B1(n10360), 
        .B2(i_data_bus[155]), .ZN(n10154) );
  ND2D1BWP30P140LVT U14749 ( .A1(n10155), .A2(n10154), .ZN(N790) );
  AOI22D1BWP30P140LVT U14750 ( .A1(n10369), .A2(i_data_bus[233]), .B1(n10367), 
        .B2(i_data_bus[201]), .ZN(n10157) );
  AOI22D1BWP30P140LVT U14751 ( .A1(n10368), .A2(i_data_bus[169]), .B1(n10360), 
        .B2(i_data_bus[137]), .ZN(n10156) );
  ND2D1BWP30P140LVT U14752 ( .A1(n10157), .A2(n10156), .ZN(N772) );
  AOI22D1BWP30P140LVT U14753 ( .A1(i_data_bus[607]), .A2(n10183), .B1(
        i_data_bus[543]), .B2(n10182), .ZN(n10159) );
  AOI22D1BWP30P140LVT U14754 ( .A1(i_data_bus[639]), .A2(n10185), .B1(
        i_data_bus[575]), .B2(n10184), .ZN(n10158) );
  ND2D1BWP30P140LVT U14755 ( .A1(n10159), .A2(n10158), .ZN(N6914) );
  AOI22D1BWP30P140LVT U14756 ( .A1(i_data_bus[630]), .A2(n10185), .B1(
        i_data_bus[598]), .B2(n10183), .ZN(n10161) );
  AOI22D1BWP30P140LVT U14757 ( .A1(i_data_bus[534]), .A2(n10182), .B1(
        i_data_bus[566]), .B2(n10184), .ZN(n10160) );
  ND2D1BWP30P140LVT U14758 ( .A1(n10161), .A2(n10160), .ZN(N6905) );
  AOI22D1BWP30P140LVT U14759 ( .A1(i_data_bus[526]), .A2(n10182), .B1(
        i_data_bus[622]), .B2(n10185), .ZN(n10163) );
  AOI22D1BWP30P140LVT U14760 ( .A1(i_data_bus[590]), .A2(n10183), .B1(
        i_data_bus[558]), .B2(n10184), .ZN(n10162) );
  ND2D1BWP30P140LVT U14761 ( .A1(n10163), .A2(n10162), .ZN(N6897) );
  AOI22D1BWP30P140LVT U14762 ( .A1(i_data_bus[584]), .A2(n10183), .B1(
        i_data_bus[616]), .B2(n10185), .ZN(n10165) );
  AOI22D1BWP30P140LVT U14763 ( .A1(i_data_bus[520]), .A2(n10182), .B1(
        i_data_bus[552]), .B2(n10184), .ZN(n10164) );
  ND2D1BWP30P140LVT U14764 ( .A1(n10165), .A2(n10164), .ZN(N6891) );
  AOI22D1BWP30P140LVT U14765 ( .A1(i_data_bus[581]), .A2(n10183), .B1(
        i_data_bus[613]), .B2(n10185), .ZN(n10167) );
  AOI22D1BWP30P140LVT U14766 ( .A1(i_data_bus[517]), .A2(n10182), .B1(
        i_data_bus[549]), .B2(n10184), .ZN(n10166) );
  ND2D1BWP30P140LVT U14767 ( .A1(n10167), .A2(n10166), .ZN(N6888) );
  AOI22D1BWP30P140LVT U14768 ( .A1(i_data_bus[537]), .A2(n10182), .B1(
        i_data_bus[601]), .B2(n10183), .ZN(n10169) );
  AOI22D1BWP30P140LVT U14769 ( .A1(i_data_bus[633]), .A2(n10185), .B1(
        i_data_bus[569]), .B2(n10184), .ZN(n10168) );
  ND2D1BWP30P140LVT U14770 ( .A1(n10169), .A2(n10168), .ZN(N6908) );
  AOI22D1BWP30P140LVT U14771 ( .A1(i_data_bus[525]), .A2(n10182), .B1(
        i_data_bus[589]), .B2(n10183), .ZN(n10171) );
  AOI22D1BWP30P140LVT U14772 ( .A1(i_data_bus[621]), .A2(n10185), .B1(
        i_data_bus[557]), .B2(n10184), .ZN(n10170) );
  ND2D1BWP30P140LVT U14773 ( .A1(n10171), .A2(n10170), .ZN(N6896) );
  AOI22D1BWP30P140LVT U14774 ( .A1(i_data_bus[578]), .A2(n10183), .B1(
        i_data_bus[514]), .B2(n10182), .ZN(n10173) );
  AOI22D1BWP30P140LVT U14775 ( .A1(i_data_bus[610]), .A2(n10185), .B1(
        i_data_bus[546]), .B2(n10184), .ZN(n10172) );
  ND2D1BWP30P140LVT U14776 ( .A1(n10173), .A2(n10172), .ZN(N6885) );
  AOI22D1BWP30P140LVT U14777 ( .A1(i_data_bus[627]), .A2(n10185), .B1(
        i_data_bus[595]), .B2(n10183), .ZN(n10175) );
  AOI22D1BWP30P140LVT U14778 ( .A1(i_data_bus[531]), .A2(n10182), .B1(
        i_data_bus[563]), .B2(n10184), .ZN(n10174) );
  ND2D1BWP30P140LVT U14779 ( .A1(n10175), .A2(n10174), .ZN(N6902) );
  AOI22D1BWP30P140LVT U14780 ( .A1(i_data_bus[512]), .A2(n10182), .B1(
        i_data_bus[608]), .B2(n10185), .ZN(n10177) );
  AOI22D1BWP30P140LVT U14781 ( .A1(i_data_bus[576]), .A2(n10183), .B1(
        i_data_bus[544]), .B2(n10184), .ZN(n10176) );
  ND2D1BWP30P140LVT U14782 ( .A1(n10177), .A2(n10176), .ZN(N6883) );
  AOI22D1BWP30P140LVT U14783 ( .A1(i_data_bus[634]), .A2(n10185), .B1(
        i_data_bus[602]), .B2(n10183), .ZN(n10179) );
  AOI22D1BWP30P140LVT U14784 ( .A1(i_data_bus[538]), .A2(n10182), .B1(
        i_data_bus[570]), .B2(n10184), .ZN(n10178) );
  ND2D1BWP30P140LVT U14785 ( .A1(n10179), .A2(n10178), .ZN(N6909) );
  AOI22D1BWP30P140LVT U14786 ( .A1(i_data_bus[533]), .A2(n10182), .B1(
        i_data_bus[597]), .B2(n10183), .ZN(n10181) );
  AOI22D1BWP30P140LVT U14787 ( .A1(i_data_bus[629]), .A2(n10185), .B1(
        i_data_bus[565]), .B2(n10184), .ZN(n10180) );
  ND2D1BWP30P140LVT U14788 ( .A1(n10181), .A2(n10180), .ZN(N6904) );
  AOI22D1BWP30P140LVT U14789 ( .A1(i_data_bus[596]), .A2(n10183), .B1(
        i_data_bus[532]), .B2(n10182), .ZN(n10187) );
  AOI22D1BWP30P140LVT U14790 ( .A1(i_data_bus[628]), .A2(n10185), .B1(
        i_data_bus[564]), .B2(n10184), .ZN(n10186) );
  ND2D1BWP30P140LVT U14791 ( .A1(n10187), .A2(n10186), .ZN(N6903) );
  AOI22D1BWP30P140LVT U14792 ( .A1(i_data_bus[206]), .A2(n10223), .B1(
        i_data_bus[238]), .B2(n10226), .ZN(n10189) );
  AOI22D1BWP30P140LVT U14793 ( .A1(i_data_bus[142]), .A2(n10224), .B1(
        i_data_bus[174]), .B2(n10225), .ZN(n10188) );
  ND2D1BWP30P140LVT U14794 ( .A1(n10189), .A2(n10188), .ZN(N6249) );
  AOI22D1BWP30P140LVT U14795 ( .A1(i_data_bus[249]), .A2(n10226), .B1(
        i_data_bus[217]), .B2(n10223), .ZN(n10191) );
  AOI22D1BWP30P140LVT U14796 ( .A1(i_data_bus[153]), .A2(n10224), .B1(
        i_data_bus[185]), .B2(n10225), .ZN(n10190) );
  ND2D1BWP30P140LVT U14797 ( .A1(n10191), .A2(n10190), .ZN(N6260) );
  AOI22D1BWP30P140LVT U14798 ( .A1(i_data_bus[131]), .A2(n10224), .B1(
        i_data_bus[227]), .B2(n10226), .ZN(n10193) );
  AOI22D1BWP30P140LVT U14799 ( .A1(i_data_bus[195]), .A2(n10223), .B1(
        i_data_bus[163]), .B2(n10225), .ZN(n10192) );
  ND2D1BWP30P140LVT U14800 ( .A1(n10193), .A2(n10192), .ZN(N6238) );
  AOI22D1BWP30P140LVT U14801 ( .A1(i_data_bus[236]), .A2(n10226), .B1(
        i_data_bus[204]), .B2(n10223), .ZN(n10195) );
  AOI22D1BWP30P140LVT U14802 ( .A1(i_data_bus[140]), .A2(n10224), .B1(
        i_data_bus[172]), .B2(n10225), .ZN(n10194) );
  ND2D1BWP30P140LVT U14803 ( .A1(n10195), .A2(n10194), .ZN(N6247) );
  AOI22D1BWP30P140LVT U14804 ( .A1(i_data_bus[215]), .A2(n10218), .B1(
        i_data_bus[247]), .B2(n10220), .ZN(n10197) );
  AOI22D1BWP30P140LVT U14805 ( .A1(i_data_bus[151]), .A2(n6213), .B1(
        i_data_bus[183]), .B2(n10219), .ZN(n10196) );
  ND2D1BWP30P140LVT U14806 ( .A1(n10197), .A2(n10196), .ZN(N2428) );
  AOI22D1BWP30P140LVT U14807 ( .A1(i_data_bus[212]), .A2(n10218), .B1(
        i_data_bus[148]), .B2(n6213), .ZN(n10199) );
  AOI22D1BWP30P140LVT U14808 ( .A1(i_data_bus[244]), .A2(n10220), .B1(
        i_data_bus[180]), .B2(n10219), .ZN(n10198) );
  ND2D1BWP30P140LVT U14809 ( .A1(n10199), .A2(n10198), .ZN(N2425) );
  AOI22D1BWP30P140LVT U14810 ( .A1(i_data_bus[146]), .A2(n6213), .B1(
        i_data_bus[242]), .B2(n10220), .ZN(n10201) );
  AOI22D1BWP30P140LVT U14811 ( .A1(i_data_bus[210]), .A2(n10218), .B1(
        i_data_bus[178]), .B2(n10219), .ZN(n10200) );
  ND2D1BWP30P140LVT U14812 ( .A1(n10201), .A2(n10200), .ZN(N2423) );
  AOI22D1BWP30P140LVT U14813 ( .A1(i_data_bus[236]), .A2(n10220), .B1(
        i_data_bus[204]), .B2(n10218), .ZN(n10203) );
  AOI22D1BWP30P140LVT U14814 ( .A1(i_data_bus[140]), .A2(n6213), .B1(
        i_data_bus[172]), .B2(n10219), .ZN(n10202) );
  ND2D1BWP30P140LVT U14815 ( .A1(n10203), .A2(n10202), .ZN(N2417) );
  AOI22D1BWP30P140LVT U14816 ( .A1(i_data_bus[136]), .A2(n6213), .B1(
        i_data_bus[200]), .B2(n10218), .ZN(n10205) );
  AOI22D1BWP30P140LVT U14817 ( .A1(i_data_bus[232]), .A2(n10220), .B1(
        i_data_bus[168]), .B2(n10219), .ZN(n10204) );
  ND2D1BWP30P140LVT U14818 ( .A1(n10205), .A2(n10204), .ZN(N2413) );
  AOI22D1BWP30P140LVT U14819 ( .A1(i_data_bus[240]), .A2(n10220), .B1(
        i_data_bus[208]), .B2(n10218), .ZN(n10207) );
  AOI22D1BWP30P140LVT U14820 ( .A1(i_data_bus[144]), .A2(n6213), .B1(
        i_data_bus[176]), .B2(n10219), .ZN(n10206) );
  ND2D1BWP30P140LVT U14821 ( .A1(n10207), .A2(n10206), .ZN(N2421) );
  AOI22D1BWP30P140LVT U14822 ( .A1(i_data_bus[244]), .A2(n10226), .B1(
        i_data_bus[148]), .B2(n10224), .ZN(n10209) );
  AOI22D1BWP30P140LVT U14823 ( .A1(i_data_bus[212]), .A2(n10223), .B1(
        i_data_bus[180]), .B2(n10225), .ZN(n10208) );
  ND2D1BWP30P140LVT U14824 ( .A1(n10209), .A2(n10208), .ZN(N6255) );
  AOI22D1BWP30P140LVT U14825 ( .A1(i_data_bus[253]), .A2(n10226), .B1(
        i_data_bus[221]), .B2(n10223), .ZN(n10211) );
  AOI22D1BWP30P140LVT U14826 ( .A1(i_data_bus[157]), .A2(n10224), .B1(
        i_data_bus[189]), .B2(n10225), .ZN(n10210) );
  ND2D1BWP30P140LVT U14827 ( .A1(n10211), .A2(n10210), .ZN(N6264) );
  AOI22D1BWP30P140LVT U14828 ( .A1(i_data_bus[222]), .A2(n10223), .B1(
        i_data_bus[158]), .B2(n10224), .ZN(n10213) );
  AOI22D1BWP30P140LVT U14829 ( .A1(i_data_bus[254]), .A2(n10226), .B1(
        i_data_bus[190]), .B2(n10225), .ZN(n10212) );
  ND2D1BWP30P140LVT U14830 ( .A1(n10213), .A2(n10212), .ZN(N6265) );
  AOI22D1BWP30P140LVT U14831 ( .A1(i_data_bus[251]), .A2(n10226), .B1(
        i_data_bus[219]), .B2(n10223), .ZN(n10215) );
  AOI22D1BWP30P140LVT U14832 ( .A1(i_data_bus[155]), .A2(n10224), .B1(
        i_data_bus[187]), .B2(n10225), .ZN(n10214) );
  ND2D1BWP30P140LVT U14833 ( .A1(n10215), .A2(n10214), .ZN(N6262) );
  AOI22D1BWP30P140LVT U14834 ( .A1(i_data_bus[231]), .A2(n10220), .B1(
        i_data_bus[135]), .B2(n6213), .ZN(n10217) );
  AOI22D1BWP30P140LVT U14835 ( .A1(i_data_bus[199]), .A2(n10218), .B1(
        i_data_bus[167]), .B2(n10219), .ZN(n10216) );
  ND2D1BWP30P140LVT U14836 ( .A1(n10217), .A2(n10216), .ZN(N2412) );
  AOI22D1BWP30P140LVT U14837 ( .A1(i_data_bus[223]), .A2(n10218), .B1(
        i_data_bus[159]), .B2(n6213), .ZN(n10222) );
  AOI22D1BWP30P140LVT U14838 ( .A1(i_data_bus[255]), .A2(n10220), .B1(
        i_data_bus[191]), .B2(n10219), .ZN(n10221) );
  ND2D1BWP30P140LVT U14839 ( .A1(n10222), .A2(n10221), .ZN(N2436) );
  AOI22D1BWP30P140LVT U14840 ( .A1(i_data_bus[134]), .A2(n10224), .B1(
        i_data_bus[198]), .B2(n10223), .ZN(n10228) );
  AOI22D1BWP30P140LVT U14841 ( .A1(i_data_bus[230]), .A2(n10226), .B1(
        i_data_bus[166]), .B2(n10225), .ZN(n10227) );
  ND2D1BWP30P140LVT U14842 ( .A1(n10228), .A2(n10227), .ZN(N6241) );
  AOI22D1BWP30P140LVT U14843 ( .A1(i_data_bus[606]), .A2(n10252), .B1(
        i_data_bus[542]), .B2(n10245), .ZN(n10230) );
  AOI22D1BWP30P140LVT U14844 ( .A1(i_data_bus[638]), .A2(n10254), .B1(
        i_data_bus[574]), .B2(n10253), .ZN(n10229) );
  ND2D1BWP30P140LVT U14845 ( .A1(n10230), .A2(n10229), .ZN(N9637) );
  AOI22D1BWP30P140LVT U14846 ( .A1(i_data_bus[586]), .A2(n10252), .B1(
        i_data_bus[522]), .B2(n10245), .ZN(n10232) );
  AOI22D1BWP30P140LVT U14847 ( .A1(i_data_bus[618]), .A2(n10254), .B1(
        i_data_bus[554]), .B2(n10253), .ZN(n10231) );
  ND2D1BWP30P140LVT U14848 ( .A1(n10232), .A2(n10231), .ZN(N9617) );
  AOI22D1BWP30P140LVT U14849 ( .A1(i_data_bus[580]), .A2(n10252), .B1(
        i_data_bus[612]), .B2(n10254), .ZN(n10234) );
  AOI22D1BWP30P140LVT U14850 ( .A1(i_data_bus[516]), .A2(n10245), .B1(
        i_data_bus[548]), .B2(n10253), .ZN(n10233) );
  ND2D1BWP30P140LVT U14851 ( .A1(n10234), .A2(n10233), .ZN(N9611) );
  AOI22D1BWP30P140LVT U14852 ( .A1(i_data_bus[526]), .A2(n10245), .B1(
        i_data_bus[622]), .B2(n10254), .ZN(n10236) );
  AOI22D1BWP30P140LVT U14853 ( .A1(i_data_bus[590]), .A2(n10252), .B1(
        i_data_bus[558]), .B2(n10253), .ZN(n10235) );
  ND2D1BWP30P140LVT U14854 ( .A1(n10236), .A2(n10235), .ZN(N9621) );
  AOI22D1BWP30P140LVT U14855 ( .A1(i_data_bus[614]), .A2(n10254), .B1(
        i_data_bus[582]), .B2(n10252), .ZN(n10238) );
  AOI22D1BWP30P140LVT U14856 ( .A1(i_data_bus[518]), .A2(n10245), .B1(
        i_data_bus[550]), .B2(n10253), .ZN(n10237) );
  ND2D1BWP30P140LVT U14857 ( .A1(n10238), .A2(n10237), .ZN(N9613) );
  AOI22D1BWP30P140LVT U14858 ( .A1(i_data_bus[521]), .A2(n10245), .B1(
        i_data_bus[617]), .B2(n10254), .ZN(n10240) );
  AOI22D1BWP30P140LVT U14859 ( .A1(i_data_bus[585]), .A2(n10252), .B1(
        i_data_bus[553]), .B2(n10253), .ZN(n10239) );
  ND2D1BWP30P140LVT U14860 ( .A1(n10240), .A2(n10239), .ZN(N9616) );
  AOI22D1BWP30P140LVT U14861 ( .A1(i_data_bus[611]), .A2(n10254), .B1(
        i_data_bus[515]), .B2(n10245), .ZN(n10242) );
  AOI22D1BWP30P140LVT U14862 ( .A1(i_data_bus[579]), .A2(n10252), .B1(
        i_data_bus[547]), .B2(n10253), .ZN(n10241) );
  ND2D1BWP30P140LVT U14863 ( .A1(n10242), .A2(n10241), .ZN(N9610) );
  AOI22D1BWP30P140LVT U14864 ( .A1(i_data_bus[584]), .A2(n10252), .B1(
        i_data_bus[616]), .B2(n10254), .ZN(n10244) );
  AOI22D1BWP30P140LVT U14865 ( .A1(i_data_bus[520]), .A2(n10245), .B1(
        i_data_bus[552]), .B2(n10253), .ZN(n10243) );
  ND2D1BWP30P140LVT U14866 ( .A1(n10244), .A2(n10243), .ZN(N9615) );
  AOI22D1BWP30P140LVT U14867 ( .A1(i_data_bus[533]), .A2(n10245), .B1(
        i_data_bus[597]), .B2(n10252), .ZN(n10247) );
  AOI22D1BWP30P140LVT U14868 ( .A1(i_data_bus[629]), .A2(n10254), .B1(
        i_data_bus[565]), .B2(n10253), .ZN(n10246) );
  ND2D1BWP30P140LVT U14869 ( .A1(n10247), .A2(n10246), .ZN(N9628) );
  AOI22D1BWP30P140LVT U14870 ( .A1(i_data_bus[512]), .A2(n10245), .B1(
        i_data_bus[576]), .B2(n10252), .ZN(n10249) );
  AOI22D1BWP30P140LVT U14871 ( .A1(i_data_bus[608]), .A2(n10254), .B1(
        i_data_bus[544]), .B2(n10253), .ZN(n10248) );
  ND2D1BWP30P140LVT U14872 ( .A1(n10249), .A2(n10248), .ZN(N9607) );
  AOI22D1BWP30P140LVT U14873 ( .A1(i_data_bus[538]), .A2(n10245), .B1(
        i_data_bus[602]), .B2(n10252), .ZN(n10251) );
  AOI22D1BWP30P140LVT U14874 ( .A1(i_data_bus[634]), .A2(n10254), .B1(
        i_data_bus[570]), .B2(n10253), .ZN(n10250) );
  ND2D1BWP30P140LVT U14875 ( .A1(n10251), .A2(n10250), .ZN(N9633) );
  AOI22D1BWP30P140LVT U14876 ( .A1(i_data_bus[578]), .A2(n10252), .B1(
        i_data_bus[514]), .B2(n10245), .ZN(n10256) );
  AOI22D1BWP30P140LVT U14877 ( .A1(i_data_bus[610]), .A2(n10254), .B1(
        i_data_bus[546]), .B2(n10253), .ZN(n10255) );
  ND2D1BWP30P140LVT U14878 ( .A1(n10256), .A2(n10255), .ZN(N9609) );
  AOI22D1BWP30P140LVT U14879 ( .A1(i_data_bus[531]), .A2(n10272), .B1(
        i_data_bus[595]), .B2(n10269), .ZN(n10258) );
  AOI22D1BWP30P140LVT U14880 ( .A1(i_data_bus[627]), .A2(n10270), .B1(
        i_data_bus[563]), .B2(n10271), .ZN(n10257) );
  ND2D1BWP30P140LVT U14881 ( .A1(n10258), .A2(n10257), .ZN(N8136) );
  AOI22D1BWP30P140LVT U14882 ( .A1(i_data_bus[578]), .A2(n10269), .B1(
        i_data_bus[514]), .B2(n10272), .ZN(n10260) );
  AOI22D1BWP30P140LVT U14883 ( .A1(i_data_bus[610]), .A2(n10270), .B1(
        i_data_bus[546]), .B2(n10271), .ZN(n10259) );
  ND2D1BWP30P140LVT U14884 ( .A1(n10260), .A2(n10259), .ZN(N8119) );
  AOI22D1BWP30P140LVT U14885 ( .A1(i_data_bus[586]), .A2(n10269), .B1(
        i_data_bus[522]), .B2(n10272), .ZN(n10262) );
  AOI22D1BWP30P140LVT U14886 ( .A1(i_data_bus[618]), .A2(n10270), .B1(
        i_data_bus[554]), .B2(n10271), .ZN(n10261) );
  ND2D1BWP30P140LVT U14887 ( .A1(n10262), .A2(n10261), .ZN(N8127) );
  AOI22D1BWP30P140LVT U14888 ( .A1(i_data_bus[585]), .A2(n10269), .B1(
        i_data_bus[617]), .B2(n10270), .ZN(n10264) );
  AOI22D1BWP30P140LVT U14889 ( .A1(i_data_bus[521]), .A2(n10272), .B1(
        i_data_bus[553]), .B2(n10271), .ZN(n10263) );
  ND2D1BWP30P140LVT U14890 ( .A1(n10264), .A2(n10263), .ZN(N8126) );
  AOI22D1BWP30P140LVT U14891 ( .A1(i_data_bus[517]), .A2(n10272), .B1(
        i_data_bus[581]), .B2(n10269), .ZN(n10266) );
  AOI22D1BWP30P140LVT U14892 ( .A1(i_data_bus[613]), .A2(n10270), .B1(
        i_data_bus[549]), .B2(n10271), .ZN(n10265) );
  ND2D1BWP30P140LVT U14893 ( .A1(n10266), .A2(n10265), .ZN(N8122) );
  AOI22D1BWP30P140LVT U14894 ( .A1(i_data_bus[512]), .A2(n10272), .B1(
        i_data_bus[576]), .B2(n10269), .ZN(n10268) );
  AOI22D1BWP30P140LVT U14895 ( .A1(i_data_bus[608]), .A2(n10270), .B1(
        i_data_bus[544]), .B2(n10271), .ZN(n10267) );
  ND2D1BWP30P140LVT U14896 ( .A1(n10268), .A2(n10267), .ZN(N8117) );
  AOI22D1BWP30P140LVT U14897 ( .A1(i_data_bus[628]), .A2(n10270), .B1(
        i_data_bus[596]), .B2(n10269), .ZN(n10274) );
  AOI22D1BWP30P140LVT U14898 ( .A1(i_data_bus[532]), .A2(n10272), .B1(
        i_data_bus[564]), .B2(n10271), .ZN(n10273) );
  ND2D1BWP30P140LVT U14899 ( .A1(n10274), .A2(n10273), .ZN(N8137) );
  AOI22D1BWP30P140LVT U14900 ( .A1(i_data_bus[301]), .A2(n10276), .B1(
        i_data_bus[333]), .B2(n10275), .ZN(n10279) );
  AOI22D1BWP30P140LVT U14901 ( .A1(i_data_bus[365]), .A2(n10277), .B1(
        i_data_bus[269]), .B2(n6227), .ZN(n10278) );
  ND2D1BWP30P140LVT U14902 ( .A1(n10279), .A2(n10278), .ZN(N9188) );
  AOI22D1BWP30P140LVT U14903 ( .A1(n10368), .A2(i_data_bus[190]), .B1(n10360), 
        .B2(i_data_bus[158]), .ZN(n10281) );
  AOI22D1BWP30P140LVT U14904 ( .A1(n10369), .A2(i_data_bus[254]), .B1(n10367), 
        .B2(i_data_bus[222]), .ZN(n10280) );
  ND2D1BWP30P140LVT U14905 ( .A1(n10281), .A2(n10280), .ZN(N793) );
  AOI22D1BWP30P140LVT U14906 ( .A1(n10369), .A2(i_data_bus[237]), .B1(n10360), 
        .B2(i_data_bus[141]), .ZN(n10283) );
  AOI22D1BWP30P140LVT U14907 ( .A1(n10368), .A2(i_data_bus[173]), .B1(n10367), 
        .B2(i_data_bus[205]), .ZN(n10282) );
  ND2D1BWP30P140LVT U14908 ( .A1(n10283), .A2(n10282), .ZN(N776) );
  AOI22D1BWP30P140LVT U14909 ( .A1(n10368), .A2(i_data_bus[167]), .B1(n10360), 
        .B2(i_data_bus[135]), .ZN(n10285) );
  AOI22D1BWP30P140LVT U14910 ( .A1(n10369), .A2(i_data_bus[231]), .B1(n10367), 
        .B2(i_data_bus[199]), .ZN(n10284) );
  ND2D1BWP30P140LVT U14911 ( .A1(n10285), .A2(n10284), .ZN(N770) );
  AOI22D1BWP30P140LVT U14912 ( .A1(n10369), .A2(i_data_bus[241]), .B1(n10360), 
        .B2(i_data_bus[145]), .ZN(n10287) );
  AOI22D1BWP30P140LVT U14913 ( .A1(n10368), .A2(i_data_bus[177]), .B1(n10367), 
        .B2(i_data_bus[209]), .ZN(n10286) );
  ND2D1BWP30P140LVT U14914 ( .A1(n10287), .A2(n10286), .ZN(N780) );
  AOI22D1BWP30P140LVT U14915 ( .A1(n10368), .A2(i_data_bus[185]), .B1(n10360), 
        .B2(i_data_bus[153]), .ZN(n10289) );
  AOI22D1BWP30P140LVT U14916 ( .A1(n10369), .A2(i_data_bus[249]), .B1(n10367), 
        .B2(i_data_bus[217]), .ZN(n10288) );
  ND2D1BWP30P140LVT U14917 ( .A1(n10289), .A2(n10288), .ZN(N788) );
  AOI22D1BWP30P140LVT U14918 ( .A1(n10368), .A2(i_data_bus[181]), .B1(n10360), 
        .B2(i_data_bus[149]), .ZN(n10291) );
  AOI22D1BWP30P140LVT U14919 ( .A1(n10369), .A2(i_data_bus[245]), .B1(n10367), 
        .B2(i_data_bus[213]), .ZN(n10290) );
  ND2D1BWP30P140LVT U14920 ( .A1(n10291), .A2(n10290), .ZN(N784) );
  AOI22D1BWP30P140LVT U14921 ( .A1(n10369), .A2(i_data_bus[246]), .B1(n10360), 
        .B2(i_data_bus[150]), .ZN(n10293) );
  AOI22D1BWP30P140LVT U14922 ( .A1(n10368), .A2(i_data_bus[182]), .B1(n10367), 
        .B2(i_data_bus[214]), .ZN(n10292) );
  ND2D1BWP30P140LVT U14923 ( .A1(n10293), .A2(n10292), .ZN(N785) );
  AOI22D1BWP30P140LVT U14924 ( .A1(n10368), .A2(i_data_bus[180]), .B1(n10360), 
        .B2(i_data_bus[148]), .ZN(n10295) );
  AOI22D1BWP30P140LVT U14925 ( .A1(n10369), .A2(i_data_bus[244]), .B1(n10367), 
        .B2(i_data_bus[212]), .ZN(n10294) );
  ND2D1BWP30P140LVT U14926 ( .A1(n10295), .A2(n10294), .ZN(N783) );
  AOI22D1BWP30P140LVT U14927 ( .A1(n10368), .A2(i_data_bus[191]), .B1(n10360), 
        .B2(i_data_bus[159]), .ZN(n10297) );
  AOI22D1BWP30P140LVT U14928 ( .A1(n10369), .A2(i_data_bus[255]), .B1(n10367), 
        .B2(i_data_bus[223]), .ZN(n10296) );
  ND2D1BWP30P140LVT U14929 ( .A1(n10297), .A2(n10296), .ZN(N794) );
  AOI22D1BWP30P140LVT U14930 ( .A1(n10369), .A2(i_data_bus[226]), .B1(n10360), 
        .B2(i_data_bus[130]), .ZN(n10299) );
  AOI22D1BWP30P140LVT U14931 ( .A1(n10368), .A2(i_data_bus[162]), .B1(n10367), 
        .B2(i_data_bus[194]), .ZN(n10298) );
  ND2D1BWP30P140LVT U14932 ( .A1(n10299), .A2(n10298), .ZN(N765) );
  AOI22D1BWP30P140LVT U14933 ( .A1(n10368), .A2(i_data_bus[165]), .B1(n10360), 
        .B2(i_data_bus[133]), .ZN(n10301) );
  AOI22D1BWP30P140LVT U14934 ( .A1(n10369), .A2(i_data_bus[229]), .B1(n10367), 
        .B2(i_data_bus[197]), .ZN(n10300) );
  ND2D1BWP30P140LVT U14935 ( .A1(n10301), .A2(n10300), .ZN(N768) );
  AOI22D1BWP30P140LVT U14936 ( .A1(n10369), .A2(i_data_bus[228]), .B1(n10360), 
        .B2(i_data_bus[132]), .ZN(n10303) );
  AOI22D1BWP30P140LVT U14937 ( .A1(n10368), .A2(i_data_bus[164]), .B1(n10367), 
        .B2(i_data_bus[196]), .ZN(n10302) );
  ND2D1BWP30P140LVT U14938 ( .A1(n10303), .A2(n10302), .ZN(N767) );
  AOI22D1BWP30P140LVT U14939 ( .A1(n10369), .A2(i_data_bus[248]), .B1(n10368), 
        .B2(i_data_bus[184]), .ZN(n10305) );
  AOI22D1BWP30P140LVT U14940 ( .A1(n10360), .A2(i_data_bus[152]), .B1(n10367), 
        .B2(i_data_bus[216]), .ZN(n10304) );
  AOI22D1BWP30P140LVT U14941 ( .A1(n10369), .A2(i_data_bus[238]), .B1(n10368), 
        .B2(i_data_bus[174]), .ZN(n10307) );
  AOI22D1BWP30P140LVT U14942 ( .A1(n10360), .A2(i_data_bus[142]), .B1(n10367), 
        .B2(i_data_bus[206]), .ZN(n10306) );
  AOI22D1BWP30P140LVT U14943 ( .A1(n10369), .A2(i_data_bus[242]), .B1(n10368), 
        .B2(i_data_bus[178]), .ZN(n10309) );
  AOI22D1BWP30P140LVT U14944 ( .A1(n10360), .A2(i_data_bus[146]), .B1(n10367), 
        .B2(i_data_bus[210]), .ZN(n10308) );
  AOI22D1BWP30P140LVT U14945 ( .A1(n10369), .A2(i_data_bus[247]), .B1(n10368), 
        .B2(i_data_bus[183]), .ZN(n10311) );
  AOI22D1BWP30P140LVT U14946 ( .A1(n10360), .A2(i_data_bus[151]), .B1(n10367), 
        .B2(i_data_bus[215]), .ZN(n10310) );
  AOI22D1BWP30P140LVT U14947 ( .A1(n10369), .A2(i_data_bus[250]), .B1(n10368), 
        .B2(i_data_bus[186]), .ZN(n10313) );
  AOI22D1BWP30P140LVT U14948 ( .A1(n10360), .A2(i_data_bus[154]), .B1(n10367), 
        .B2(i_data_bus[218]), .ZN(n10312) );
  AOI22D1BWP30P140LVT U14949 ( .A1(i_data_bus[498]), .A2(n10385), .B1(
        i_data_bus[402]), .B2(n10387), .ZN(n10315) );
  AOI22D1BWP30P140LVT U14950 ( .A1(i_data_bus[434]), .A2(n10386), .B1(
        i_data_bus[466]), .B2(n10388), .ZN(n10314) );
  ND2D1BWP30P140LVT U14951 ( .A1(n10315), .A2(n10314), .ZN(N10771) );
  AOI22D1BWP30P140LVT U14952 ( .A1(i_data_bus[438]), .A2(n10386), .B1(
        i_data_bus[406]), .B2(n10387), .ZN(n10317) );
  AOI22D1BWP30P140LVT U14953 ( .A1(i_data_bus[502]), .A2(n10385), .B1(
        i_data_bus[470]), .B2(n10388), .ZN(n10316) );
  ND2D1BWP30P140LVT U14954 ( .A1(n10317), .A2(n10316), .ZN(N10775) );
  AOI22D1BWP30P140LVT U14955 ( .A1(i_data_bus[506]), .A2(n10385), .B1(
        i_data_bus[410]), .B2(n10387), .ZN(n10319) );
  AOI22D1BWP30P140LVT U14956 ( .A1(i_data_bus[474]), .A2(n10388), .B1(
        i_data_bus[442]), .B2(n10386), .ZN(n10318) );
  ND2D1BWP30P140LVT U14957 ( .A1(n10319), .A2(n10318), .ZN(N10779) );
  AOI22D1BWP30P140LVT U14958 ( .A1(i_data_bus[507]), .A2(n10385), .B1(
        i_data_bus[411]), .B2(n10387), .ZN(n10321) );
  AOI22D1BWP30P140LVT U14959 ( .A1(i_data_bus[475]), .A2(n10388), .B1(
        i_data_bus[443]), .B2(n10386), .ZN(n10320) );
  ND2D1BWP30P140LVT U14960 ( .A1(n10321), .A2(n10320), .ZN(N10780) );
  AOI22D1BWP30P140LVT U14961 ( .A1(i_data_bus[469]), .A2(n10388), .B1(
        i_data_bus[405]), .B2(n10387), .ZN(n10323) );
  AOI22D1BWP30P140LVT U14962 ( .A1(i_data_bus[501]), .A2(n10385), .B1(
        i_data_bus[437]), .B2(n10386), .ZN(n10322) );
  ND2D1BWP30P140LVT U14963 ( .A1(n10323), .A2(n10322), .ZN(N10774) );
  AOI22D1BWP30P140LVT U14964 ( .A1(i_data_bus[511]), .A2(n10385), .B1(
        i_data_bus[415]), .B2(n10387), .ZN(n10325) );
  AOI22D1BWP30P140LVT U14965 ( .A1(i_data_bus[479]), .A2(n10388), .B1(
        i_data_bus[447]), .B2(n10386), .ZN(n10324) );
  ND2D1BWP30P140LVT U14966 ( .A1(n10325), .A2(n10324), .ZN(N10784) );
  AOI22D1BWP30P140LVT U14967 ( .A1(i_data_bus[425]), .A2(n10386), .B1(
        i_data_bus[393]), .B2(n10387), .ZN(n10327) );
  AOI22D1BWP30P140LVT U14968 ( .A1(i_data_bus[457]), .A2(n10388), .B1(
        i_data_bus[489]), .B2(n10385), .ZN(n10326) );
  ND2D1BWP30P140LVT U14969 ( .A1(n10327), .A2(n10326), .ZN(N10762) );
  AOI22D1BWP30P140LVT U14970 ( .A1(i_data_bus[417]), .A2(n10405), .B1(
        i_data_bus[385]), .B2(n10407), .ZN(n10329) );
  AOI22D1BWP30P140LVT U14971 ( .A1(i_data_bus[449]), .A2(n10408), .B1(
        i_data_bus[481]), .B2(n10406), .ZN(n10328) );
  ND2D1BWP30P140LVT U14972 ( .A1(n10329), .A2(n10328), .ZN(N9392) );
  AOI22D1BWP30P140LVT U14973 ( .A1(i_data_bus[457]), .A2(n10408), .B1(
        i_data_bus[393]), .B2(n10407), .ZN(n10331) );
  AOI22D1BWP30P140LVT U14974 ( .A1(i_data_bus[425]), .A2(n10405), .B1(
        i_data_bus[489]), .B2(n10406), .ZN(n10330) );
  ND2D1BWP30P140LVT U14975 ( .A1(n10331), .A2(n10330), .ZN(N9400) );
  AOI22D1BWP30P140LVT U14976 ( .A1(i_data_bus[419]), .A2(n10405), .B1(
        i_data_bus[387]), .B2(n10407), .ZN(n10333) );
  AOI22D1BWP30P140LVT U14977 ( .A1(i_data_bus[451]), .A2(n10408), .B1(
        i_data_bus[483]), .B2(n10406), .ZN(n10332) );
  ND2D1BWP30P140LVT U14978 ( .A1(n10333), .A2(n10332), .ZN(N9394) );
  AOI22D1BWP30P140LVT U14979 ( .A1(i_data_bus[420]), .A2(n10405), .B1(
        i_data_bus[388]), .B2(n10407), .ZN(n10335) );
  AOI22D1BWP30P140LVT U14980 ( .A1(i_data_bus[452]), .A2(n10408), .B1(
        i_data_bus[484]), .B2(n10406), .ZN(n10334) );
  ND2D1BWP30P140LVT U14981 ( .A1(n10335), .A2(n10334), .ZN(N9395) );
  AOI22D1BWP30P140LVT U14982 ( .A1(i_data_bus[511]), .A2(n10406), .B1(
        i_data_bus[415]), .B2(n10407), .ZN(n10337) );
  AOI22D1BWP30P140LVT U14983 ( .A1(i_data_bus[479]), .A2(n10408), .B1(
        i_data_bus[447]), .B2(n10405), .ZN(n10336) );
  ND2D1BWP30P140LVT U14984 ( .A1(n10337), .A2(n10336), .ZN(N9422) );
  AOI22D1BWP30P140LVT U14985 ( .A1(i_data_bus[444]), .A2(n10405), .B1(
        i_data_bus[412]), .B2(n10407), .ZN(n10339) );
  AOI22D1BWP30P140LVT U14986 ( .A1(i_data_bus[508]), .A2(n10406), .B1(
        i_data_bus[476]), .B2(n10408), .ZN(n10338) );
  ND2D1BWP30P140LVT U14987 ( .A1(n10339), .A2(n10338), .ZN(N9419) );
  AOI22D1BWP30P140LVT U14988 ( .A1(i_data_bus[428]), .A2(n10405), .B1(
        i_data_bus[396]), .B2(n10407), .ZN(n10341) );
  AOI22D1BWP30P140LVT U14989 ( .A1(i_data_bus[492]), .A2(n10406), .B1(
        i_data_bus[460]), .B2(n10408), .ZN(n10340) );
  ND2D1BWP30P140LVT U14990 ( .A1(n10341), .A2(n10340), .ZN(N9403) );
  AOI22D1BWP30P140LVT U14991 ( .A1(i_data_bus[421]), .A2(n10405), .B1(
        i_data_bus[389]), .B2(n10407), .ZN(n10343) );
  AOI22D1BWP30P140LVT U14992 ( .A1(i_data_bus[485]), .A2(n10406), .B1(
        i_data_bus[453]), .B2(n10408), .ZN(n10342) );
  ND2D1BWP30P140LVT U14993 ( .A1(n10343), .A2(n10342), .ZN(N9396) );
  AOI22D1BWP30P140LVT U14994 ( .A1(i_data_bus[480]), .A2(n10406), .B1(
        i_data_bus[384]), .B2(n10407), .ZN(n10345) );
  AOI22D1BWP30P140LVT U14995 ( .A1(i_data_bus[416]), .A2(n10405), .B1(
        i_data_bus[448]), .B2(n10408), .ZN(n10344) );
  ND2D1BWP30P140LVT U14996 ( .A1(n10345), .A2(n10344), .ZN(N9391) );
  AOI22D1BWP30P140LVT U14997 ( .A1(i_data_bus[434]), .A2(n10405), .B1(
        i_data_bus[402]), .B2(n10407), .ZN(n10347) );
  AOI22D1BWP30P140LVT U14998 ( .A1(i_data_bus[498]), .A2(n10406), .B1(
        i_data_bus[466]), .B2(n10408), .ZN(n10346) );
  ND2D1BWP30P140LVT U14999 ( .A1(n10347), .A2(n10346), .ZN(N9409) );
  AOI22D1BWP30P140LVT U15000 ( .A1(i_data_bus[440]), .A2(n10427), .B1(
        i_data_bus[408]), .B2(n10429), .ZN(n10349) );
  AOI22D1BWP30P140LVT U15001 ( .A1(i_data_bus[504]), .A2(n10428), .B1(
        i_data_bus[472]), .B2(n10430), .ZN(n10348) );
  ND2D1BWP30P140LVT U15002 ( .A1(n10349), .A2(n10348), .ZN(N6691) );
  AOI22D1BWP30P140LVT U15003 ( .A1(i_data_bus[488]), .A2(n10428), .B1(
        i_data_bus[392]), .B2(n10429), .ZN(n10351) );
  AOI22D1BWP30P140LVT U15004 ( .A1(i_data_bus[456]), .A2(n10430), .B1(
        i_data_bus[424]), .B2(n10427), .ZN(n10350) );
  ND2D1BWP30P140LVT U15005 ( .A1(n10351), .A2(n10350), .ZN(N6675) );
  AOI22D1BWP30P140LVT U15006 ( .A1(i_data_bus[495]), .A2(n10428), .B1(
        i_data_bus[399]), .B2(n10429), .ZN(n10353) );
  AOI22D1BWP30P140LVT U15007 ( .A1(i_data_bus[463]), .A2(n10430), .B1(
        i_data_bus[431]), .B2(n10427), .ZN(n10352) );
  ND2D1BWP30P140LVT U15008 ( .A1(n10353), .A2(n10352), .ZN(N6682) );
  AOI22D1BWP30P140LVT U15009 ( .A1(i_data_bus[419]), .A2(n10427), .B1(
        i_data_bus[387]), .B2(n10429), .ZN(n10355) );
  AOI22D1BWP30P140LVT U15010 ( .A1(i_data_bus[451]), .A2(n10430), .B1(
        i_data_bus[483]), .B2(n10428), .ZN(n10354) );
  ND2D1BWP30P140LVT U15011 ( .A1(n10355), .A2(n10354), .ZN(N6670) );
  AOI22D1BWP30P140LVT U15012 ( .A1(i_data_bus[416]), .A2(n10427), .B1(
        i_data_bus[384]), .B2(n10429), .ZN(n10357) );
  AOI22D1BWP30P140LVT U15013 ( .A1(i_data_bus[448]), .A2(n10430), .B1(
        i_data_bus[480]), .B2(n10428), .ZN(n10356) );
  ND2D1BWP30P140LVT U15014 ( .A1(n10357), .A2(n10356), .ZN(N6667) );
  AOI22D1BWP30P140LVT U15015 ( .A1(i_data_bus[128]), .A2(n10360), .B1(
        i_data_bus[192]), .B2(n10367), .ZN(n10359) );
  AOI22D1BWP30P140LVT U15016 ( .A1(i_data_bus[224]), .A2(n10369), .B1(
        i_data_bus[160]), .B2(n10368), .ZN(n10358) );
  AOI22D1BWP30P140LVT U15017 ( .A1(n10360), .A2(i_data_bus[129]), .B1(n10367), 
        .B2(i_data_bus[193]), .ZN(n10362) );
  AOI22D1BWP30P140LVT U15018 ( .A1(n10369), .A2(i_data_bus[225]), .B1(n10368), 
        .B2(i_data_bus[161]), .ZN(n10361) );
  AOI22D1BWP30P140LVT U15019 ( .A1(n10360), .A2(i_data_bus[147]), .B1(n10367), 
        .B2(i_data_bus[211]), .ZN(n10364) );
  AOI22D1BWP30P140LVT U15020 ( .A1(n10369), .A2(i_data_bus[243]), .B1(n10368), 
        .B2(i_data_bus[179]), .ZN(n10363) );
  AOI22D1BWP30P140LVT U15021 ( .A1(n10360), .A2(i_data_bus[156]), .B1(n10367), 
        .B2(i_data_bus[220]), .ZN(n10366) );
  AOI22D1BWP30P140LVT U15022 ( .A1(n10369), .A2(i_data_bus[252]), .B1(n10368), 
        .B2(i_data_bus[188]), .ZN(n10365) );
  AOI22D1BWP30P140LVT U15023 ( .A1(n10360), .A2(i_data_bus[134]), .B1(n10367), 
        .B2(i_data_bus[198]), .ZN(n10371) );
  AOI22D1BWP30P140LVT U15024 ( .A1(n10369), .A2(i_data_bus[230]), .B1(n10368), 
        .B2(i_data_bus[166]), .ZN(n10370) );
  INR4D1BWP30P140LVT U15025 ( .A1(i_cmd[16]), .B1(i_cmd[0]), .B2(n10372), .B3(
        n10632), .ZN(n10589) );
  NR4D1BWP30P140LVT U15026 ( .A1(i_cmd[8]), .A2(n10373), .A3(n10375), .A4(
        n10630), .ZN(n10588) );
  AOI22D1BWP30P140LVT U15027 ( .A1(i_data_bus[64]), .A2(n10589), .B1(
        i_data_bus[96]), .B2(n10588), .ZN(n10378) );
  NR4D1BWP30P140LVT U15028 ( .A1(i_cmd[24]), .A2(n10376), .A3(n10634), .A4(
        n10375), .ZN(n10587) );
  AOI22D1BWP30P140LVT U15029 ( .A1(i_data_bus[0]), .A2(n6221), .B1(
        i_data_bus[32]), .B2(n10587), .ZN(n10377) );
  AOI22D1BWP30P140LVT U15030 ( .A1(i_data_bus[416]), .A2(n10386), .B1(
        i_data_bus[480]), .B2(n10385), .ZN(n10380) );
  AOI22D1BWP30P140LVT U15031 ( .A1(i_data_bus[448]), .A2(n10388), .B1(
        i_data_bus[384]), .B2(n10387), .ZN(n10379) );
  ND2D1BWP30P140LVT U15032 ( .A1(n10380), .A2(n10379), .ZN(N10753) );
  AOI22D1BWP30P140LVT U15033 ( .A1(i_data_bus[449]), .A2(n10388), .B1(
        i_data_bus[417]), .B2(n10386), .ZN(n10382) );
  AOI22D1BWP30P140LVT U15034 ( .A1(i_data_bus[481]), .A2(n10385), .B1(
        i_data_bus[385]), .B2(n10387), .ZN(n10381) );
  ND2D1BWP30P140LVT U15035 ( .A1(n10382), .A2(n10381), .ZN(N10754) );
  AOI22D1BWP30P140LVT U15036 ( .A1(i_data_bus[488]), .A2(n10385), .B1(
        i_data_bus[424]), .B2(n10386), .ZN(n10384) );
  AOI22D1BWP30P140LVT U15037 ( .A1(i_data_bus[456]), .A2(n10388), .B1(
        i_data_bus[392]), .B2(n10387), .ZN(n10383) );
  ND2D1BWP30P140LVT U15038 ( .A1(n10384), .A2(n10383), .ZN(N10761) );
  AOI22D1BWP30P140LVT U15039 ( .A1(i_data_bus[419]), .A2(n10386), .B1(
        i_data_bus[483]), .B2(n10385), .ZN(n10390) );
  AOI22D1BWP30P140LVT U15040 ( .A1(i_data_bus[451]), .A2(n10388), .B1(
        i_data_bus[387]), .B2(n10387), .ZN(n10389) );
  ND2D1BWP30P140LVT U15041 ( .A1(n10390), .A2(n10389), .ZN(N10756) );
  NR4D1BWP30P140LVT U15042 ( .A1(i_cmd[88]), .A2(n11172), .A3(n10391), .A4(
        n10393), .ZN(n10554) );
  NR4D1BWP30P140LVT U15043 ( .A1(i_cmd[72]), .A2(n11171), .A3(n10393), .A4(
        n10392), .ZN(n10553) );
  AOI22D1BWP30P140LVT U15044 ( .A1(n10554), .A2(i_data_bus[318]), .B1(n10553), 
        .B2(i_data_bus[382]), .ZN(n10397) );
  NR3D0P7BWP30P140LVT U15045 ( .A1(i_cmd[80]), .A2(i_cmd[72]), .A3(i_cmd[88]), 
        .ZN(n11168) );
  INR4D1BWP30P140LVT U15046 ( .A1(i_cmd[80]), .B1(i_cmd[64]), .B2(n11169), 
        .B3(n10395), .ZN(n10551) );
  AOI22D1BWP30P140LVT U15047 ( .A1(n10552), .A2(i_data_bus[286]), .B1(n10551), 
        .B2(i_data_bus[350]), .ZN(n10396) );
  NR4D1BWP30P140LVT U15048 ( .A1(i_cmd[136]), .A2(n11164), .A3(n10694), .A4(
        n10398), .ZN(n10624) );
  NR4D1BWP30P140LVT U15049 ( .A1(i_cmd[152]), .A2(n11165), .A3(n10398), .A4(
        n10696), .ZN(n10626) );
  AOI22D1BWP30P140LVT U15050 ( .A1(i_data_bus[608]), .A2(n10624), .B1(
        i_data_bus[544]), .B2(n10626), .ZN(n10400) );
  NR3D0P7BWP30P140LVT U15051 ( .A1(i_cmd[136]), .A2(i_cmd[152]), .A3(
        i_cmd[144]), .ZN(n11161) );
  INR4D1BWP30P140LVT U15052 ( .A1(i_cmd[144]), .B1(i_cmd[128]), .B2(n11162), 
        .B3(n10692), .ZN(n10625) );
  AOI22D1BWP30P140LVT U15053 ( .A1(i_data_bus[512]), .A2(n6220), .B1(
        i_data_bus[576]), .B2(n10625), .ZN(n10399) );
  AOI22D1BWP30P140LVT U15054 ( .A1(i_data_bus[504]), .A2(n10406), .B1(
        i_data_bus[472]), .B2(n10408), .ZN(n10402) );
  AOI22D1BWP30P140LVT U15055 ( .A1(i_data_bus[440]), .A2(n10405), .B1(
        i_data_bus[408]), .B2(n10407), .ZN(n10401) );
  ND2D1BWP30P140LVT U15056 ( .A1(n10402), .A2(n10401), .ZN(N9415) );
  AOI22D1BWP30P140LVT U15057 ( .A1(i_data_bus[475]), .A2(n10408), .B1(
        i_data_bus[443]), .B2(n10405), .ZN(n10404) );
  AOI22D1BWP30P140LVT U15058 ( .A1(i_data_bus[507]), .A2(n10406), .B1(
        i_data_bus[411]), .B2(n10407), .ZN(n10403) );
  ND2D1BWP30P140LVT U15059 ( .A1(n10404), .A2(n10403), .ZN(N9418) );
  AOI22D1BWP30P140LVT U15060 ( .A1(i_data_bus[488]), .A2(n10406), .B1(
        i_data_bus[424]), .B2(n10405), .ZN(n10410) );
  AOI22D1BWP30P140LVT U15061 ( .A1(i_data_bus[456]), .A2(n10408), .B1(
        i_data_bus[392]), .B2(n10407), .ZN(n10409) );
  ND2D1BWP30P140LVT U15062 ( .A1(n10410), .A2(n10409), .ZN(N9399) );
  AOI22D1BWP30P140LVT U15063 ( .A1(i_data_bus[425]), .A2(n10427), .B1(
        i_data_bus[489]), .B2(n10428), .ZN(n10412) );
  AOI22D1BWP30P140LVT U15064 ( .A1(i_data_bus[457]), .A2(n10430), .B1(
        i_data_bus[393]), .B2(n10429), .ZN(n10411) );
  ND2D1BWP30P140LVT U15065 ( .A1(n10412), .A2(n10411), .ZN(N6676) );
  AOI22D1BWP30P140LVT U15066 ( .A1(i_data_bus[511]), .A2(n10428), .B1(
        i_data_bus[447]), .B2(n10427), .ZN(n10414) );
  AOI22D1BWP30P140LVT U15067 ( .A1(i_data_bus[479]), .A2(n10430), .B1(
        i_data_bus[415]), .B2(n10429), .ZN(n10413) );
  ND2D1BWP30P140LVT U15068 ( .A1(n10414), .A2(n10413), .ZN(N6698) );
  AOI22D1BWP30P140LVT U15069 ( .A1(i_data_bus[508]), .A2(n10428), .B1(
        i_data_bus[476]), .B2(n10430), .ZN(n10416) );
  AOI22D1BWP30P140LVT U15070 ( .A1(i_data_bus[444]), .A2(n10427), .B1(
        i_data_bus[412]), .B2(n10429), .ZN(n10415) );
  ND2D1BWP30P140LVT U15071 ( .A1(n10416), .A2(n10415), .ZN(N6695) );
  AOI22D1BWP30P140LVT U15072 ( .A1(i_data_bus[506]), .A2(n10428), .B1(
        i_data_bus[442]), .B2(n10427), .ZN(n10418) );
  AOI22D1BWP30P140LVT U15073 ( .A1(i_data_bus[474]), .A2(n10430), .B1(
        i_data_bus[410]), .B2(n10429), .ZN(n10417) );
  ND2D1BWP30P140LVT U15074 ( .A1(n10418), .A2(n10417), .ZN(N6693) );
  AOI22D1BWP30P140LVT U15075 ( .A1(i_data_bus[502]), .A2(n10428), .B1(
        i_data_bus[470]), .B2(n10430), .ZN(n10420) );
  AOI22D1BWP30P140LVT U15076 ( .A1(i_data_bus[438]), .A2(n10427), .B1(
        i_data_bus[406]), .B2(n10429), .ZN(n10419) );
  ND2D1BWP30P140LVT U15077 ( .A1(n10420), .A2(n10419), .ZN(N6689) );
  AOI22D1BWP30P140LVT U15078 ( .A1(i_data_bus[449]), .A2(n10430), .B1(
        i_data_bus[481]), .B2(n10428), .ZN(n10422) );
  AOI22D1BWP30P140LVT U15079 ( .A1(i_data_bus[417]), .A2(n10427), .B1(
        i_data_bus[385]), .B2(n10429), .ZN(n10421) );
  ND2D1BWP30P140LVT U15080 ( .A1(n10422), .A2(n10421), .ZN(N6668) );
  AOI22D1BWP30P140LVT U15081 ( .A1(i_data_bus[498]), .A2(n10428), .B1(
        i_data_bus[466]), .B2(n10430), .ZN(n10424) );
  AOI22D1BWP30P140LVT U15082 ( .A1(i_data_bus[434]), .A2(n10427), .B1(
        i_data_bus[402]), .B2(n10429), .ZN(n10423) );
  ND2D1BWP30P140LVT U15083 ( .A1(n10424), .A2(n10423), .ZN(N6685) );
  AOI22D1BWP30P140LVT U15084 ( .A1(i_data_bus[475]), .A2(n10430), .B1(
        i_data_bus[443]), .B2(n10427), .ZN(n10426) );
  AOI22D1BWP30P140LVT U15085 ( .A1(i_data_bus[507]), .A2(n10428), .B1(
        i_data_bus[411]), .B2(n10429), .ZN(n10425) );
  ND2D1BWP30P140LVT U15086 ( .A1(n10426), .A2(n10425), .ZN(N6694) );
  AOI22D1BWP30P140LVT U15087 ( .A1(i_data_bus[501]), .A2(n10428), .B1(
        i_data_bus[437]), .B2(n10427), .ZN(n10432) );
  AOI22D1BWP30P140LVT U15088 ( .A1(i_data_bus[469]), .A2(n10430), .B1(
        i_data_bus[405]), .B2(n10429), .ZN(n10431) );
  ND2D1BWP30P140LVT U15089 ( .A1(n10432), .A2(n10431), .ZN(N6688) );
  AOI22D1BWP30P140LVT U15090 ( .A1(n10589), .A2(i_data_bus[75]), .B1(n10588), 
        .B2(i_data_bus[107]), .ZN(n10434) );
  AOI22D1BWP30P140LVT U15091 ( .A1(n6221), .A2(i_data_bus[11]), .B1(n10587), 
        .B2(i_data_bus[43]), .ZN(n10433) );
  AOI22D1BWP30P140LVT U15092 ( .A1(n10589), .A2(i_data_bus[80]), .B1(n10588), 
        .B2(i_data_bus[112]), .ZN(n10436) );
  AOI22D1BWP30P140LVT U15093 ( .A1(n6221), .A2(i_data_bus[16]), .B1(n10587), 
        .B2(i_data_bus[48]), .ZN(n10435) );
  AOI22D1BWP30P140LVT U15094 ( .A1(n10589), .A2(i_data_bus[77]), .B1(n10588), 
        .B2(i_data_bus[109]), .ZN(n10438) );
  AOI22D1BWP30P140LVT U15095 ( .A1(n6221), .A2(i_data_bus[13]), .B1(n10587), 
        .B2(i_data_bus[45]), .ZN(n10437) );
  AOI22D1BWP30P140LVT U15096 ( .A1(n10589), .A2(i_data_bus[94]), .B1(n10588), 
        .B2(i_data_bus[126]), .ZN(n10440) );
  AOI22D1BWP30P140LVT U15097 ( .A1(n6221), .A2(i_data_bus[30]), .B1(n10587), 
        .B2(i_data_bus[62]), .ZN(n10439) );
  AOI22D1BWP30P140LVT U15098 ( .A1(n10587), .A2(i_data_bus[46]), .B1(n10588), 
        .B2(i_data_bus[110]), .ZN(n10442) );
  AOI22D1BWP30P140LVT U15099 ( .A1(n6221), .A2(i_data_bus[14]), .B1(n10589), 
        .B2(i_data_bus[78]), .ZN(n10441) );
  AOI22D1BWP30P140LVT U15100 ( .A1(n10587), .A2(i_data_bus[49]), .B1(n10588), 
        .B2(i_data_bus[113]), .ZN(n10444) );
  AOI22D1BWP30P140LVT U15101 ( .A1(n6221), .A2(i_data_bus[17]), .B1(n10589), 
        .B2(i_data_bus[81]), .ZN(n10443) );
  AOI22D1BWP30P140LVT U15102 ( .A1(n6221), .A2(i_data_bus[28]), .B1(n10588), 
        .B2(i_data_bus[124]), .ZN(n10446) );
  AOI22D1BWP30P140LVT U15103 ( .A1(n10587), .A2(i_data_bus[60]), .B1(n10589), 
        .B2(i_data_bus[92]), .ZN(n10445) );
  AOI22D1BWP30P140LVT U15104 ( .A1(n10587), .A2(i_data_bus[39]), .B1(n10588), 
        .B2(i_data_bus[103]), .ZN(n10448) );
  AOI22D1BWP30P140LVT U15105 ( .A1(n6221), .A2(i_data_bus[7]), .B1(n10589), 
        .B2(i_data_bus[71]), .ZN(n10447) );
  AOI22D1BWP30P140LVT U15106 ( .A1(n6221), .A2(i_data_bus[9]), .B1(n10588), 
        .B2(i_data_bus[105]), .ZN(n10450) );
  AOI22D1BWP30P140LVT U15107 ( .A1(n10587), .A2(i_data_bus[41]), .B1(n10589), 
        .B2(i_data_bus[73]), .ZN(n10449) );
  AOI22D1BWP30P140LVT U15108 ( .A1(n6221), .A2(i_data_bus[23]), .B1(n10588), 
        .B2(i_data_bus[119]), .ZN(n10452) );
  AOI22D1BWP30P140LVT U15109 ( .A1(n10587), .A2(i_data_bus[55]), .B1(n10589), 
        .B2(i_data_bus[87]), .ZN(n10451) );
  AOI22D1BWP30P140LVT U15110 ( .A1(n10587), .A2(i_data_bus[56]), .B1(n10588), 
        .B2(i_data_bus[120]), .ZN(n10454) );
  AOI22D1BWP30P140LVT U15111 ( .A1(n6221), .A2(i_data_bus[24]), .B1(n10589), 
        .B2(i_data_bus[88]), .ZN(n10453) );
  AOI22D1BWP30P140LVT U15112 ( .A1(n6221), .A2(i_data_bus[18]), .B1(n10588), 
        .B2(i_data_bus[114]), .ZN(n10456) );
  AOI22D1BWP30P140LVT U15113 ( .A1(n10587), .A2(i_data_bus[50]), .B1(n10589), 
        .B2(i_data_bus[82]), .ZN(n10455) );
  AOI22D1BWP30P140LVT U15114 ( .A1(n10587), .A2(i_data_bus[51]), .B1(n10588), 
        .B2(i_data_bus[115]), .ZN(n10458) );
  AOI22D1BWP30P140LVT U15115 ( .A1(n6221), .A2(i_data_bus[19]), .B1(n10589), 
        .B2(i_data_bus[83]), .ZN(n10457) );
  AOI22D1BWP30P140LVT U15116 ( .A1(n6221), .A2(i_data_bus[29]), .B1(n10588), 
        .B2(i_data_bus[125]), .ZN(n10460) );
  AOI22D1BWP30P140LVT U15117 ( .A1(n10587), .A2(i_data_bus[61]), .B1(n10589), 
        .B2(i_data_bus[93]), .ZN(n10459) );
  AOI22D1BWP30P140LVT U15118 ( .A1(n10587), .A2(i_data_bus[52]), .B1(n10588), 
        .B2(i_data_bus[116]), .ZN(n10462) );
  AOI22D1BWP30P140LVT U15119 ( .A1(n6221), .A2(i_data_bus[20]), .B1(n10589), 
        .B2(i_data_bus[84]), .ZN(n10461) );
  AOI22D1BWP30P140LVT U15120 ( .A1(n6220), .A2(i_data_bus[532]), .B1(n10626), 
        .B2(i_data_bus[564]), .ZN(n10464) );
  AOI22D1BWP30P140LVT U15121 ( .A1(n10625), .A2(i_data_bus[596]), .B1(n10624), 
        .B2(i_data_bus[628]), .ZN(n10463) );
  AOI22D1BWP30P140LVT U15122 ( .A1(n6220), .A2(i_data_bus[514]), .B1(n10626), 
        .B2(i_data_bus[546]), .ZN(n10466) );
  AOI22D1BWP30P140LVT U15123 ( .A1(n10625), .A2(i_data_bus[578]), .B1(n10624), 
        .B2(i_data_bus[610]), .ZN(n10465) );
  AOI22D1BWP30P140LVT U15124 ( .A1(n6220), .A2(i_data_bus[522]), .B1(n10626), 
        .B2(i_data_bus[554]), .ZN(n10468) );
  AOI22D1BWP30P140LVT U15125 ( .A1(n10625), .A2(i_data_bus[586]), .B1(n10624), 
        .B2(i_data_bus[618]), .ZN(n10467) );
  AOI22D1BWP30P140LVT U15126 ( .A1(n10625), .A2(i_data_bus[597]), .B1(n10626), 
        .B2(i_data_bus[565]), .ZN(n10470) );
  AOI22D1BWP30P140LVT U15127 ( .A1(n6220), .A2(i_data_bus[533]), .B1(n10624), 
        .B2(i_data_bus[629]), .ZN(n10469) );
  AOI22D1BWP30P140LVT U15128 ( .A1(n10625), .A2(i_data_bus[598]), .B1(n10626), 
        .B2(i_data_bus[566]), .ZN(n10472) );
  AOI22D1BWP30P140LVT U15129 ( .A1(n6220), .A2(i_data_bus[534]), .B1(n10624), 
        .B2(i_data_bus[630]), .ZN(n10471) );
  AOI22D1BWP30P140LVT U15130 ( .A1(n10625), .A2(i_data_bus[595]), .B1(n10626), 
        .B2(i_data_bus[563]), .ZN(n10474) );
  AOI22D1BWP30P140LVT U15131 ( .A1(n6220), .A2(i_data_bus[531]), .B1(n10624), 
        .B2(i_data_bus[627]), .ZN(n10473) );
  AOI22D1BWP30P140LVT U15132 ( .A1(n10625), .A2(i_data_bus[589]), .B1(n10626), 
        .B2(i_data_bus[557]), .ZN(n10476) );
  AOI22D1BWP30P140LVT U15133 ( .A1(n6220), .A2(i_data_bus[525]), .B1(n10624), 
        .B2(i_data_bus[621]), .ZN(n10475) );
  AOI22D1BWP30P140LVT U15134 ( .A1(n6220), .A2(i_data_bus[543]), .B1(n10626), 
        .B2(i_data_bus[575]), .ZN(n10478) );
  AOI22D1BWP30P140LVT U15135 ( .A1(n10625), .A2(i_data_bus[607]), .B1(n10624), 
        .B2(i_data_bus[639]), .ZN(n10477) );
  AOI22D1BWP30P140LVT U15136 ( .A1(n6220), .A2(i_data_bus[520]), .B1(n10626), 
        .B2(i_data_bus[552]), .ZN(n10480) );
  AOI22D1BWP30P140LVT U15137 ( .A1(n10625), .A2(i_data_bus[584]), .B1(n10624), 
        .B2(i_data_bus[616]), .ZN(n10479) );
  AOI22D1BWP30P140LVT U15138 ( .A1(n6220), .A2(i_data_bus[523]), .B1(n10626), 
        .B2(i_data_bus[555]), .ZN(n10482) );
  AOI22D1BWP30P140LVT U15139 ( .A1(n10625), .A2(i_data_bus[587]), .B1(n10624), 
        .B2(i_data_bus[619]), .ZN(n10481) );
  AOI22D1BWP30P140LVT U15140 ( .A1(n10625), .A2(i_data_bus[602]), .B1(n10626), 
        .B2(i_data_bus[570]), .ZN(n10484) );
  AOI22D1BWP30P140LVT U15141 ( .A1(n6220), .A2(i_data_bus[538]), .B1(n10624), 
        .B2(i_data_bus[634]), .ZN(n10483) );
  AOI22D1BWP30P140LVT U15142 ( .A1(n6220), .A2(i_data_bus[542]), .B1(n10626), 
        .B2(i_data_bus[574]), .ZN(n10486) );
  AOI22D1BWP30P140LVT U15143 ( .A1(n10625), .A2(i_data_bus[606]), .B1(n10624), 
        .B2(i_data_bus[638]), .ZN(n10485) );
  AOI22D1BWP30P140LVT U15144 ( .A1(n10624), .A2(i_data_bus[617]), .B1(n10626), 
        .B2(i_data_bus[553]), .ZN(n10488) );
  AOI22D1BWP30P140LVT U15145 ( .A1(n6220), .A2(i_data_bus[521]), .B1(n10625), 
        .B2(i_data_bus[585]), .ZN(n10487) );
  AOI22D1BWP30P140LVT U15146 ( .A1(n10624), .A2(i_data_bus[613]), .B1(n10626), 
        .B2(i_data_bus[549]), .ZN(n10490) );
  AOI22D1BWP30P140LVT U15147 ( .A1(n6220), .A2(i_data_bus[517]), .B1(n10625), 
        .B2(i_data_bus[581]), .ZN(n10489) );
  AOI22D1BWP30P140LVT U15148 ( .A1(n10552), .A2(i_data_bus[257]), .B1(n10553), 
        .B2(i_data_bus[353]), .ZN(n10492) );
  AOI22D1BWP30P140LVT U15149 ( .A1(n10551), .A2(i_data_bus[321]), .B1(n10554), 
        .B2(i_data_bus[289]), .ZN(n10491) );
  AOI22D1BWP30P140LVT U15150 ( .A1(n10551), .A2(i_data_bus[348]), .B1(n10553), 
        .B2(i_data_bus[380]), .ZN(n10494) );
  AOI22D1BWP30P140LVT U15151 ( .A1(n10552), .A2(i_data_bus[284]), .B1(n10554), 
        .B2(i_data_bus[316]), .ZN(n10493) );
  AOI22D1BWP30P140LVT U15152 ( .A1(n10552), .A2(i_data_bus[271]), .B1(n10553), 
        .B2(i_data_bus[367]), .ZN(n10496) );
  AOI22D1BWP30P140LVT U15153 ( .A1(n10551), .A2(i_data_bus[335]), .B1(n10554), 
        .B2(i_data_bus[303]), .ZN(n10495) );
  AOI22D1BWP30P140LVT U15154 ( .A1(n10552), .A2(i_data_bus[258]), .B1(n10553), 
        .B2(i_data_bus[354]), .ZN(n10498) );
  AOI22D1BWP30P140LVT U15155 ( .A1(n10551), .A2(i_data_bus[322]), .B1(n10554), 
        .B2(i_data_bus[290]), .ZN(n10497) );
  AOI22D1BWP30P140LVT U15156 ( .A1(n10552), .A2(i_data_bus[287]), .B1(n10553), 
        .B2(i_data_bus[383]), .ZN(n10500) );
  AOI22D1BWP30P140LVT U15157 ( .A1(n10551), .A2(i_data_bus[351]), .B1(n10554), 
        .B2(i_data_bus[319]), .ZN(n10499) );
  AOI22D1BWP30P140LVT U15158 ( .A1(n10552), .A2(i_data_bus[285]), .B1(n10553), 
        .B2(i_data_bus[381]), .ZN(n10502) );
  AOI22D1BWP30P140LVT U15159 ( .A1(n10551), .A2(i_data_bus[349]), .B1(n10554), 
        .B2(i_data_bus[317]), .ZN(n10501) );
  AOI22D1BWP30P140LVT U15160 ( .A1(n10551), .A2(i_data_bus[330]), .B1(n10553), 
        .B2(i_data_bus[362]), .ZN(n10504) );
  AOI22D1BWP30P140LVT U15161 ( .A1(n10552), .A2(i_data_bus[266]), .B1(n10554), 
        .B2(i_data_bus[298]), .ZN(n10503) );
  AOI22D1BWP30P140LVT U15162 ( .A1(i_data_bus[288]), .A2(n10554), .B1(
        i_data_bus[352]), .B2(n10553), .ZN(n10506) );
  AOI22D1BWP30P140LVT U15163 ( .A1(i_data_bus[256]), .A2(n10552), .B1(
        i_data_bus[320]), .B2(n10551), .ZN(n10505) );
  AOI22D1BWP30P140LVT U15164 ( .A1(n10551), .A2(i_data_bus[324]), .B1(n10553), 
        .B2(i_data_bus[356]), .ZN(n10508) );
  AOI22D1BWP30P140LVT U15165 ( .A1(n10552), .A2(i_data_bus[260]), .B1(n10554), 
        .B2(i_data_bus[292]), .ZN(n10507) );
  AOI22D1BWP30P140LVT U15166 ( .A1(n10551), .A2(i_data_bus[347]), .B1(n10553), 
        .B2(i_data_bus[379]), .ZN(n10510) );
  AOI22D1BWP30P140LVT U15167 ( .A1(n10552), .A2(i_data_bus[283]), .B1(n10554), 
        .B2(i_data_bus[315]), .ZN(n10509) );
  AOI22D1BWP30P140LVT U15168 ( .A1(n10551), .A2(i_data_bus[343]), .B1(n10553), 
        .B2(i_data_bus[375]), .ZN(n10512) );
  AOI22D1BWP30P140LVT U15169 ( .A1(n10552), .A2(i_data_bus[279]), .B1(n10554), 
        .B2(i_data_bus[311]), .ZN(n10511) );
  AOI22D1BWP30P140LVT U15170 ( .A1(n10551), .A2(i_data_bus[342]), .B1(n10553), 
        .B2(i_data_bus[374]), .ZN(n10514) );
  AOI22D1BWP30P140LVT U15171 ( .A1(n10552), .A2(i_data_bus[278]), .B1(n10554), 
        .B2(i_data_bus[310]), .ZN(n10513) );
  AOI22D1BWP30P140LVT U15172 ( .A1(n10551), .A2(i_data_bus[334]), .B1(n10553), 
        .B2(i_data_bus[366]), .ZN(n10516) );
  AOI22D1BWP30P140LVT U15173 ( .A1(n10552), .A2(i_data_bus[270]), .B1(n10554), 
        .B2(i_data_bus[302]), .ZN(n10515) );
  AOI22D1BWP30P140LVT U15174 ( .A1(n10551), .A2(i_data_bus[327]), .B1(n10553), 
        .B2(i_data_bus[359]), .ZN(n10518) );
  AOI22D1BWP30P140LVT U15175 ( .A1(n10552), .A2(i_data_bus[263]), .B1(n10554), 
        .B2(i_data_bus[295]), .ZN(n10517) );
  AOI22D1BWP30P140LVT U15176 ( .A1(n10551), .A2(i_data_bus[336]), .B1(n10553), 
        .B2(i_data_bus[368]), .ZN(n10520) );
  AOI22D1BWP30P140LVT U15177 ( .A1(n10552), .A2(i_data_bus[272]), .B1(n10554), 
        .B2(i_data_bus[304]), .ZN(n10519) );
  AOI22D1BWP30P140LVT U15178 ( .A1(n10554), .A2(i_data_bus[306]), .B1(n10553), 
        .B2(i_data_bus[370]), .ZN(n10522) );
  AOI22D1BWP30P140LVT U15179 ( .A1(n10552), .A2(i_data_bus[274]), .B1(n10551), 
        .B2(i_data_bus[338]), .ZN(n10521) );
  AOI22D1BWP30P140LVT U15180 ( .A1(n10551), .A2(i_data_bus[332]), .B1(n10554), 
        .B2(i_data_bus[300]), .ZN(n10524) );
  AOI22D1BWP30P140LVT U15181 ( .A1(n10552), .A2(i_data_bus[268]), .B1(n10553), 
        .B2(i_data_bus[364]), .ZN(n10523) );
  AOI22D1BWP30P140LVT U15182 ( .A1(n10552), .A2(i_data_bus[276]), .B1(n10554), 
        .B2(i_data_bus[308]), .ZN(n10526) );
  AOI22D1BWP30P140LVT U15183 ( .A1(n10551), .A2(i_data_bus[340]), .B1(n10553), 
        .B2(i_data_bus[372]), .ZN(n10525) );
  AOI22D1BWP30P140LVT U15184 ( .A1(n10552), .A2(i_data_bus[281]), .B1(n10551), 
        .B2(i_data_bus[345]), .ZN(n10528) );
  AOI22D1BWP30P140LVT U15185 ( .A1(n10554), .A2(i_data_bus[313]), .B1(n10553), 
        .B2(i_data_bus[377]), .ZN(n10527) );
  AOI22D1BWP30P140LVT U15186 ( .A1(n10552), .A2(i_data_bus[280]), .B1(n10551), 
        .B2(i_data_bus[344]), .ZN(n10530) );
  AOI22D1BWP30P140LVT U15187 ( .A1(n10554), .A2(i_data_bus[312]), .B1(n10553), 
        .B2(i_data_bus[376]), .ZN(n10529) );
  AOI22D1BWP30P140LVT U15188 ( .A1(n10552), .A2(i_data_bus[282]), .B1(n10554), 
        .B2(i_data_bus[314]), .ZN(n10532) );
  AOI22D1BWP30P140LVT U15189 ( .A1(n10551), .A2(i_data_bus[346]), .B1(n10553), 
        .B2(i_data_bus[378]), .ZN(n10531) );
  AOI22D1BWP30P140LVT U15190 ( .A1(n10552), .A2(i_data_bus[267]), .B1(n10551), 
        .B2(i_data_bus[331]), .ZN(n10534) );
  AOI22D1BWP30P140LVT U15191 ( .A1(n10554), .A2(i_data_bus[299]), .B1(n10553), 
        .B2(i_data_bus[363]), .ZN(n10533) );
  AOI22D1BWP30P140LVT U15192 ( .A1(n10552), .A2(i_data_bus[269]), .B1(n10551), 
        .B2(i_data_bus[333]), .ZN(n10536) );
  AOI22D1BWP30P140LVT U15193 ( .A1(n10554), .A2(i_data_bus[301]), .B1(n10553), 
        .B2(i_data_bus[365]), .ZN(n10535) );
  AOI22D1BWP30P140LVT U15194 ( .A1(n10552), .A2(i_data_bus[264]), .B1(n10554), 
        .B2(i_data_bus[296]), .ZN(n10538) );
  AOI22D1BWP30P140LVT U15195 ( .A1(n10551), .A2(i_data_bus[328]), .B1(n10553), 
        .B2(i_data_bus[360]), .ZN(n10537) );
  AOI22D1BWP30P140LVT U15196 ( .A1(n10551), .A2(i_data_bus[339]), .B1(n10554), 
        .B2(i_data_bus[307]), .ZN(n10540) );
  AOI22D1BWP30P140LVT U15197 ( .A1(n10552), .A2(i_data_bus[275]), .B1(n10553), 
        .B2(i_data_bus[371]), .ZN(n10539) );
  AOI22D1BWP30P140LVT U15198 ( .A1(n10551), .A2(i_data_bus[325]), .B1(n10554), 
        .B2(i_data_bus[293]), .ZN(n10542) );
  AOI22D1BWP30P140LVT U15199 ( .A1(n10552), .A2(i_data_bus[261]), .B1(n10553), 
        .B2(i_data_bus[357]), .ZN(n10541) );
  AOI22D1BWP30P140LVT U15200 ( .A1(n10551), .A2(i_data_bus[326]), .B1(n10554), 
        .B2(i_data_bus[294]), .ZN(n10544) );
  AOI22D1BWP30P140LVT U15201 ( .A1(n10552), .A2(i_data_bus[262]), .B1(n10553), 
        .B2(i_data_bus[358]), .ZN(n10543) );
  AOI22D1BWP30P140LVT U15202 ( .A1(n10552), .A2(i_data_bus[265]), .B1(n10551), 
        .B2(i_data_bus[329]), .ZN(n10546) );
  AOI22D1BWP30P140LVT U15203 ( .A1(n10554), .A2(i_data_bus[297]), .B1(n10553), 
        .B2(i_data_bus[361]), .ZN(n10545) );
  AOI22D1BWP30P140LVT U15204 ( .A1(n10551), .A2(i_data_bus[323]), .B1(n10554), 
        .B2(i_data_bus[291]), .ZN(n10548) );
  AOI22D1BWP30P140LVT U15205 ( .A1(n10552), .A2(i_data_bus[259]), .B1(n10553), 
        .B2(i_data_bus[355]), .ZN(n10547) );
  AOI22D1BWP30P140LVT U15206 ( .A1(n10552), .A2(i_data_bus[273]), .B1(n10554), 
        .B2(i_data_bus[305]), .ZN(n10550) );
  AOI22D1BWP30P140LVT U15207 ( .A1(n10551), .A2(i_data_bus[337]), .B1(n10553), 
        .B2(i_data_bus[369]), .ZN(n10549) );
  AOI22D1BWP30P140LVT U15208 ( .A1(n10552), .A2(i_data_bus[277]), .B1(n10551), 
        .B2(i_data_bus[341]), .ZN(n10556) );
  AOI22D1BWP30P140LVT U15209 ( .A1(n10554), .A2(i_data_bus[309]), .B1(n10553), 
        .B2(i_data_bus[373]), .ZN(n10555) );
  AOI22D1BWP30P140LVT U15210 ( .A1(n10587), .A2(i_data_bus[38]), .B1(n10589), 
        .B2(i_data_bus[70]), .ZN(n10558) );
  AOI22D1BWP30P140LVT U15211 ( .A1(n6221), .A2(i_data_bus[6]), .B1(n10588), 
        .B2(i_data_bus[102]), .ZN(n10557) );
  AOI22D1BWP30P140LVT U15212 ( .A1(n6221), .A2(i_data_bus[3]), .B1(n10589), 
        .B2(i_data_bus[67]), .ZN(n10560) );
  AOI22D1BWP30P140LVT U15213 ( .A1(n10587), .A2(i_data_bus[35]), .B1(n10588), 
        .B2(i_data_bus[99]), .ZN(n10559) );
  AOI22D1BWP30P140LVT U15214 ( .A1(n10587), .A2(i_data_bus[37]), .B1(n10589), 
        .B2(i_data_bus[69]), .ZN(n10562) );
  AOI22D1BWP30P140LVT U15215 ( .A1(n6221), .A2(i_data_bus[5]), .B1(n10588), 
        .B2(i_data_bus[101]), .ZN(n10561) );
  AOI22D1BWP30P140LVT U15216 ( .A1(n6221), .A2(i_data_bus[22]), .B1(n10587), 
        .B2(i_data_bus[54]), .ZN(n10564) );
  AOI22D1BWP30P140LVT U15217 ( .A1(n10589), .A2(i_data_bus[86]), .B1(n10588), 
        .B2(i_data_bus[118]), .ZN(n10563) );
  AOI22D1BWP30P140LVT U15218 ( .A1(n6221), .A2(i_data_bus[4]), .B1(n10589), 
        .B2(i_data_bus[68]), .ZN(n10566) );
  AOI22D1BWP30P140LVT U15219 ( .A1(n10587), .A2(i_data_bus[36]), .B1(n10588), 
        .B2(i_data_bus[100]), .ZN(n10565) );
  AOI22D1BWP30P140LVT U15220 ( .A1(n10587), .A2(i_data_bus[47]), .B1(n10589), 
        .B2(i_data_bus[79]), .ZN(n10568) );
  AOI22D1BWP30P140LVT U15221 ( .A1(n6221), .A2(i_data_bus[15]), .B1(n10588), 
        .B2(i_data_bus[111]), .ZN(n10567) );
  AOI22D1BWP30P140LVT U15222 ( .A1(n10587), .A2(i_data_bus[33]), .B1(n10589), 
        .B2(i_data_bus[65]), .ZN(n10570) );
  AOI22D1BWP30P140LVT U15223 ( .A1(n6221), .A2(i_data_bus[1]), .B1(n10588), 
        .B2(i_data_bus[97]), .ZN(n10569) );
  AOI22D1BWP30P140LVT U15224 ( .A1(n10587), .A2(i_data_bus[57]), .B1(n10589), 
        .B2(i_data_bus[89]), .ZN(n10572) );
  AOI22D1BWP30P140LVT U15225 ( .A1(n6221), .A2(i_data_bus[25]), .B1(n10588), 
        .B2(i_data_bus[121]), .ZN(n10571) );
  AOI22D1BWP30P140LVT U15226 ( .A1(n6221), .A2(i_data_bus[2]), .B1(n10589), 
        .B2(i_data_bus[66]), .ZN(n10574) );
  AOI22D1BWP30P140LVT U15227 ( .A1(n10587), .A2(i_data_bus[34]), .B1(n10588), 
        .B2(i_data_bus[98]), .ZN(n10573) );
  AOI22D1BWP30P140LVT U15228 ( .A1(n10587), .A2(i_data_bus[58]), .B1(n10589), 
        .B2(i_data_bus[90]), .ZN(n10576) );
  AOI22D1BWP30P140LVT U15229 ( .A1(n6221), .A2(i_data_bus[26]), .B1(n10588), 
        .B2(i_data_bus[122]), .ZN(n10575) );
  AOI22D1BWP30P140LVT U15230 ( .A1(n6221), .A2(i_data_bus[10]), .B1(n10587), 
        .B2(i_data_bus[42]), .ZN(n10578) );
  AOI22D1BWP30P140LVT U15231 ( .A1(n10589), .A2(i_data_bus[74]), .B1(n10588), 
        .B2(i_data_bus[106]), .ZN(n10577) );
  AOI22D1BWP30P140LVT U15232 ( .A1(n6221), .A2(i_data_bus[12]), .B1(n10587), 
        .B2(i_data_bus[44]), .ZN(n10580) );
  AOI22D1BWP30P140LVT U15233 ( .A1(n10589), .A2(i_data_bus[76]), .B1(n10588), 
        .B2(i_data_bus[108]), .ZN(n10579) );
  AOI22D1BWP30P140LVT U15234 ( .A1(n10587), .A2(i_data_bus[40]), .B1(n10589), 
        .B2(i_data_bus[72]), .ZN(n10582) );
  AOI22D1BWP30P140LVT U15235 ( .A1(n6221), .A2(i_data_bus[8]), .B1(n10588), 
        .B2(i_data_bus[104]), .ZN(n10581) );
  AOI22D1BWP30P140LVT U15236 ( .A1(n10587), .A2(i_data_bus[53]), .B1(n10589), 
        .B2(i_data_bus[85]), .ZN(n10584) );
  AOI22D1BWP30P140LVT U15237 ( .A1(n6221), .A2(i_data_bus[21]), .B1(n10588), 
        .B2(i_data_bus[117]), .ZN(n10583) );
  AOI22D1BWP30P140LVT U15238 ( .A1(n10587), .A2(i_data_bus[59]), .B1(n10589), 
        .B2(i_data_bus[91]), .ZN(n10586) );
  AOI22D1BWP30P140LVT U15239 ( .A1(n6221), .A2(i_data_bus[27]), .B1(n10588), 
        .B2(i_data_bus[123]), .ZN(n10585) );
  AOI22D1BWP30P140LVT U15240 ( .A1(n6221), .A2(i_data_bus[31]), .B1(n10587), 
        .B2(i_data_bus[63]), .ZN(n10591) );
  AOI22D1BWP30P140LVT U15241 ( .A1(n10589), .A2(i_data_bus[95]), .B1(n10588), 
        .B2(i_data_bus[127]), .ZN(n10590) );
  AOI22D1BWP30P140LVT U15242 ( .A1(n6220), .A2(i_data_bus[536]), .B1(n10624), 
        .B2(i_data_bus[632]), .ZN(n10593) );
  AOI22D1BWP30P140LVT U15243 ( .A1(n10625), .A2(i_data_bus[600]), .B1(n10626), 
        .B2(i_data_bus[568]), .ZN(n10592) );
  AOI22D1BWP30P140LVT U15244 ( .A1(n6220), .A2(i_data_bus[540]), .B1(n10624), 
        .B2(i_data_bus[636]), .ZN(n10595) );
  AOI22D1BWP30P140LVT U15245 ( .A1(n10625), .A2(i_data_bus[604]), .B1(n10626), 
        .B2(i_data_bus[572]), .ZN(n10594) );
  AOI22D1BWP30P140LVT U15246 ( .A1(n6220), .A2(i_data_bus[515]), .B1(n10624), 
        .B2(i_data_bus[611]), .ZN(n10597) );
  AOI22D1BWP30P140LVT U15247 ( .A1(n10625), .A2(i_data_bus[579]), .B1(n10626), 
        .B2(i_data_bus[547]), .ZN(n10596) );
  AOI22D1BWP30P140LVT U15248 ( .A1(n10625), .A2(i_data_bus[582]), .B1(n10624), 
        .B2(i_data_bus[614]), .ZN(n10599) );
  AOI22D1BWP30P140LVT U15249 ( .A1(n6220), .A2(i_data_bus[518]), .B1(n10626), 
        .B2(i_data_bus[550]), .ZN(n10598) );
  AOI22D1BWP30P140LVT U15250 ( .A1(n6220), .A2(i_data_bus[527]), .B1(n10625), 
        .B2(i_data_bus[591]), .ZN(n10601) );
  AOI22D1BWP30P140LVT U15251 ( .A1(n10624), .A2(i_data_bus[623]), .B1(n10626), 
        .B2(i_data_bus[559]), .ZN(n10600) );
  AOI22D1BWP30P140LVT U15252 ( .A1(n6220), .A2(i_data_bus[513]), .B1(n10625), 
        .B2(i_data_bus[577]), .ZN(n10603) );
  AOI22D1BWP30P140LVT U15253 ( .A1(n10624), .A2(i_data_bus[609]), .B1(n10626), 
        .B2(i_data_bus[545]), .ZN(n10602) );
  AOI22D1BWP30P140LVT U15254 ( .A1(n6220), .A2(i_data_bus[519]), .B1(n10624), 
        .B2(i_data_bus[615]), .ZN(n10605) );
  AOI22D1BWP30P140LVT U15255 ( .A1(n10625), .A2(i_data_bus[583]), .B1(n10626), 
        .B2(i_data_bus[551]), .ZN(n10604) );
  AOI22D1BWP30P140LVT U15256 ( .A1(n6220), .A2(i_data_bus[528]), .B1(n10625), 
        .B2(i_data_bus[592]), .ZN(n10607) );
  AOI22D1BWP30P140LVT U15257 ( .A1(n10624), .A2(i_data_bus[624]), .B1(n10626), 
        .B2(i_data_bus[560]), .ZN(n10606) );
  AOI22D1BWP30P140LVT U15258 ( .A1(n6220), .A2(i_data_bus[535]), .B1(n10625), 
        .B2(i_data_bus[599]), .ZN(n10609) );
  AOI22D1BWP30P140LVT U15259 ( .A1(n10624), .A2(i_data_bus[631]), .B1(n10626), 
        .B2(i_data_bus[567]), .ZN(n10608) );
  AOI22D1BWP30P140LVT U15260 ( .A1(n6220), .A2(i_data_bus[537]), .B1(n10625), 
        .B2(i_data_bus[601]), .ZN(n10611) );
  AOI22D1BWP30P140LVT U15261 ( .A1(n10624), .A2(i_data_bus[633]), .B1(n10626), 
        .B2(i_data_bus[569]), .ZN(n10610) );
  AOI22D1BWP30P140LVT U15262 ( .A1(n6220), .A2(i_data_bus[526]), .B1(n10624), 
        .B2(i_data_bus[622]), .ZN(n10613) );
  AOI22D1BWP30P140LVT U15263 ( .A1(n10625), .A2(i_data_bus[590]), .B1(n10626), 
        .B2(i_data_bus[558]), .ZN(n10612) );
  AOI22D1BWP30P140LVT U15264 ( .A1(n6220), .A2(i_data_bus[539]), .B1(n10624), 
        .B2(i_data_bus[635]), .ZN(n10615) );
  AOI22D1BWP30P140LVT U15265 ( .A1(n10625), .A2(i_data_bus[603]), .B1(n10626), 
        .B2(i_data_bus[571]), .ZN(n10614) );
  AOI22D1BWP30P140LVT U15266 ( .A1(n10625), .A2(i_data_bus[593]), .B1(n10624), 
        .B2(i_data_bus[625]), .ZN(n10617) );
  AOI22D1BWP30P140LVT U15267 ( .A1(n6220), .A2(i_data_bus[529]), .B1(n10626), 
        .B2(i_data_bus[561]), .ZN(n10616) );
  AOI22D1BWP30P140LVT U15268 ( .A1(n6220), .A2(i_data_bus[541]), .B1(n10625), 
        .B2(i_data_bus[605]), .ZN(n10619) );
  AOI22D1BWP30P140LVT U15269 ( .A1(n10624), .A2(i_data_bus[637]), .B1(n10626), 
        .B2(i_data_bus[573]), .ZN(n10618) );
  AOI22D1BWP30P140LVT U15270 ( .A1(n10625), .A2(i_data_bus[580]), .B1(n10624), 
        .B2(i_data_bus[612]), .ZN(n10621) );
  AOI22D1BWP30P140LVT U15271 ( .A1(n6220), .A2(i_data_bus[516]), .B1(n10626), 
        .B2(i_data_bus[548]), .ZN(n10620) );
  AOI22D1BWP30P140LVT U15272 ( .A1(n6220), .A2(i_data_bus[524]), .B1(n10625), 
        .B2(i_data_bus[588]), .ZN(n10623) );
  AOI22D1BWP30P140LVT U15273 ( .A1(n10624), .A2(i_data_bus[620]), .B1(n10626), 
        .B2(i_data_bus[556]), .ZN(n10622) );
  AOI22D1BWP30P140LVT U15274 ( .A1(n10625), .A2(i_data_bus[594]), .B1(n10624), 
        .B2(i_data_bus[626]), .ZN(n10628) );
  AOI22D1BWP30P140LVT U15275 ( .A1(n6220), .A2(i_data_bus[530]), .B1(n10626), 
        .B2(i_data_bus[562]), .ZN(n10627) );
  NR3D0P7BWP30P140LVT U15276 ( .A1(i_cmd[23]), .A2(i_cmd[15]), .A3(i_cmd[31]), 
        .ZN(n10934) );
  NR4D1BWP30P140LVT U15277 ( .A1(i_cmd[15]), .A2(n10630), .A3(n10631), .A4(
        n10633), .ZN(n10811) );
  AOI22D1BWP30P140LVT U15278 ( .A1(i_data_bus[24]), .A2(n10812), .B1(
        i_data_bus[120]), .B2(n10811), .ZN(n10637) );
  INR4D1BWP30P140LVT U15279 ( .A1(i_cmd[23]), .B1(i_cmd[7]), .B2(n10632), .B3(
        n10938), .ZN(n10810) );
  NR4D1BWP30P140LVT U15280 ( .A1(i_cmd[31]), .A2(n10635), .A3(n10634), .A4(
        n10633), .ZN(n10813) );
  AOI22D1BWP30P140LVT U15281 ( .A1(i_data_bus[88]), .A2(n10810), .B1(
        i_data_bus[56]), .B2(n10813), .ZN(n10636) );
  ND2D1BWP30P140LVT U15282 ( .A1(n10637), .A2(n10636), .ZN(N10513) );
  AOI22D1BWP30P140LVT U15283 ( .A1(i_data_bus[26]), .A2(n10812), .B1(
        i_data_bus[90]), .B2(n10810), .ZN(n10639) );
  AOI22D1BWP30P140LVT U15284 ( .A1(i_data_bus[122]), .A2(n10811), .B1(
        i_data_bus[58]), .B2(n10813), .ZN(n10638) );
  ND2D1BWP30P140LVT U15285 ( .A1(n10639), .A2(n10638), .ZN(N10515) );
  AOI22D1BWP30P140LVT U15286 ( .A1(i_data_bus[25]), .A2(n10812), .B1(
        i_data_bus[121]), .B2(n10811), .ZN(n10641) );
  AOI22D1BWP30P140LVT U15287 ( .A1(i_data_bus[89]), .A2(n10810), .B1(
        i_data_bus[57]), .B2(n10813), .ZN(n10640) );
  ND2D1BWP30P140LVT U15288 ( .A1(n10641), .A2(n10640), .ZN(N10514) );
  AOI22D1BWP30P140LVT U15289 ( .A1(i_data_bus[5]), .A2(n10812), .B1(
        i_data_bus[101]), .B2(n10811), .ZN(n10643) );
  AOI22D1BWP30P140LVT U15290 ( .A1(i_data_bus[69]), .A2(n10810), .B1(
        i_data_bus[37]), .B2(n10813), .ZN(n10642) );
  ND2D1BWP30P140LVT U15291 ( .A1(n10643), .A2(n10642), .ZN(N10494) );
  AOI22D1BWP30P140LVT U15292 ( .A1(i_data_bus[9]), .A2(n10812), .B1(
        i_data_bus[105]), .B2(n10811), .ZN(n10645) );
  AOI22D1BWP30P140LVT U15293 ( .A1(i_data_bus[73]), .A2(n10810), .B1(
        i_data_bus[41]), .B2(n10813), .ZN(n10644) );
  ND2D1BWP30P140LVT U15294 ( .A1(n10645), .A2(n10644), .ZN(N10498) );
  AOI22D1BWP30P140LVT U15295 ( .A1(i_data_bus[20]), .A2(n10812), .B1(
        i_data_bus[52]), .B2(n10813), .ZN(n10647) );
  AOI22D1BWP30P140LVT U15296 ( .A1(i_data_bus[84]), .A2(n10810), .B1(
        i_data_bus[116]), .B2(n10811), .ZN(n10646) );
  ND2D1BWP30P140LVT U15297 ( .A1(n10647), .A2(n10646), .ZN(N10509) );
  AOI22D1BWP30P140LVT U15298 ( .A1(i_data_bus[17]), .A2(n10812), .B1(
        i_data_bus[49]), .B2(n10813), .ZN(n10649) );
  AOI22D1BWP30P140LVT U15299 ( .A1(i_data_bus[81]), .A2(n10810), .B1(
        i_data_bus[113]), .B2(n10811), .ZN(n10648) );
  ND2D1BWP30P140LVT U15300 ( .A1(n10649), .A2(n10648), .ZN(N10506) );
  AOI22D1BWP30P140LVT U15301 ( .A1(i_data_bus[19]), .A2(n10812), .B1(
        i_data_bus[83]), .B2(n10810), .ZN(n10651) );
  AOI22D1BWP30P140LVT U15302 ( .A1(i_data_bus[51]), .A2(n10813), .B1(
        i_data_bus[115]), .B2(n10811), .ZN(n10650) );
  ND2D1BWP30P140LVT U15303 ( .A1(n10651), .A2(n10650), .ZN(N10508) );
  AOI22D1BWP30P140LVT U15304 ( .A1(i_data_bus[30]), .A2(n10812), .B1(
        i_data_bus[94]), .B2(n10810), .ZN(n10653) );
  AOI22D1BWP30P140LVT U15305 ( .A1(i_data_bus[62]), .A2(n10813), .B1(
        i_data_bus[126]), .B2(n10811), .ZN(n10652) );
  ND2D1BWP30P140LVT U15306 ( .A1(n10653), .A2(n10652), .ZN(N10519) );
  AOI22D1BWP30P140LVT U15307 ( .A1(i_data_bus[7]), .A2(n10812), .B1(
        i_data_bus[39]), .B2(n10813), .ZN(n10655) );
  AOI22D1BWP30P140LVT U15308 ( .A1(i_data_bus[71]), .A2(n10810), .B1(
        i_data_bus[103]), .B2(n10811), .ZN(n10654) );
  ND2D1BWP30P140LVT U15309 ( .A1(n10655), .A2(n10654), .ZN(N10496) );
  AOI22D1BWP30P140LVT U15310 ( .A1(i_data_bus[28]), .A2(n10812), .B1(
        i_data_bus[124]), .B2(n10811), .ZN(n10657) );
  AOI22D1BWP30P140LVT U15311 ( .A1(i_data_bus[60]), .A2(n10813), .B1(
        i_data_bus[92]), .B2(n10810), .ZN(n10656) );
  ND2D1BWP30P140LVT U15312 ( .A1(n10657), .A2(n10656), .ZN(N10517) );
  AOI22D1BWP30P140LVT U15313 ( .A1(i_data_bus[1]), .A2(n10812), .B1(
        i_data_bus[33]), .B2(n10813), .ZN(n10659) );
  AOI22D1BWP30P140LVT U15314 ( .A1(i_data_bus[97]), .A2(n10811), .B1(
        i_data_bus[65]), .B2(n10810), .ZN(n10658) );
  ND2D1BWP30P140LVT U15315 ( .A1(n10659), .A2(n10658), .ZN(N10490) );
  AOI22D1BWP30P140LVT U15316 ( .A1(i_data_bus[11]), .A2(n10812), .B1(
        i_data_bus[107]), .B2(n10811), .ZN(n10661) );
  AOI22D1BWP30P140LVT U15317 ( .A1(i_data_bus[43]), .A2(n10813), .B1(
        i_data_bus[75]), .B2(n10810), .ZN(n10660) );
  ND2D1BWP30P140LVT U15318 ( .A1(n10661), .A2(n10660), .ZN(N10500) );
  NR4D1BWP30P140LVT U15319 ( .A1(i_cmd[63]), .A2(n10665), .A3(n10664), .A4(
        n10668), .ZN(n10829) );
  AOI22D1BWP30P140LVT U15320 ( .A1(i_data_bus[149]), .A2(n10830), .B1(
        i_data_bus[181]), .B2(n10829), .ZN(n10672) );
  INR4D1BWP30P140LVT U15321 ( .A1(i_cmd[55]), .B1(i_cmd[39]), .B2(n10667), 
        .B3(n10666), .ZN(n10828) );
  NR4D1BWP30P140LVT U15322 ( .A1(i_cmd[47]), .A2(n10670), .A3(n10669), .A4(
        n10668), .ZN(n10831) );
  AOI22D1BWP30P140LVT U15323 ( .A1(i_data_bus[213]), .A2(n10828), .B1(
        i_data_bus[245]), .B2(n10831), .ZN(n10671) );
  ND2D1BWP30P140LVT U15324 ( .A1(n10672), .A2(n10671), .ZN(N10598) );
  AOI22D1BWP30P140LVT U15325 ( .A1(i_data_bus[142]), .A2(n10830), .B1(
        i_data_bus[206]), .B2(n10828), .ZN(n10674) );
  AOI22D1BWP30P140LVT U15326 ( .A1(i_data_bus[174]), .A2(n10829), .B1(
        i_data_bus[238]), .B2(n10831), .ZN(n10673) );
  ND2D1BWP30P140LVT U15327 ( .A1(n10674), .A2(n10673), .ZN(N10591) );
  AOI22D1BWP30P140LVT U15328 ( .A1(i_data_bus[154]), .A2(n10830), .B1(
        i_data_bus[218]), .B2(n10828), .ZN(n10676) );
  AOI22D1BWP30P140LVT U15329 ( .A1(i_data_bus[186]), .A2(n10829), .B1(
        i_data_bus[250]), .B2(n10831), .ZN(n10675) );
  ND2D1BWP30P140LVT U15330 ( .A1(n10676), .A2(n10675), .ZN(N10603) );
  AOI22D1BWP30P140LVT U15331 ( .A1(i_data_bus[152]), .A2(n10830), .B1(
        i_data_bus[216]), .B2(n10828), .ZN(n10678) );
  AOI22D1BWP30P140LVT U15332 ( .A1(i_data_bus[184]), .A2(n10829), .B1(
        i_data_bus[248]), .B2(n10831), .ZN(n10677) );
  ND2D1BWP30P140LVT U15333 ( .A1(n10678), .A2(n10677), .ZN(N10601) );
  AOI22D1BWP30P140LVT U15334 ( .A1(i_data_bus[145]), .A2(n10830), .B1(
        i_data_bus[241]), .B2(n10831), .ZN(n10680) );
  AOI22D1BWP30P140LVT U15335 ( .A1(i_data_bus[209]), .A2(n10828), .B1(
        i_data_bus[177]), .B2(n10829), .ZN(n10679) );
  ND2D1BWP30P140LVT U15336 ( .A1(n10680), .A2(n10679), .ZN(N10594) );
  AOI22D1BWP30P140LVT U15337 ( .A1(i_data_bus[150]), .A2(n10830), .B1(
        i_data_bus[246]), .B2(n10831), .ZN(n10682) );
  AOI22D1BWP30P140LVT U15338 ( .A1(i_data_bus[214]), .A2(n10828), .B1(
        i_data_bus[182]), .B2(n10829), .ZN(n10681) );
  ND2D1BWP30P140LVT U15339 ( .A1(n10682), .A2(n10681), .ZN(N10599) );
  AOI22D1BWP30P140LVT U15340 ( .A1(i_data_bus[146]), .A2(n10830), .B1(
        i_data_bus[242]), .B2(n10831), .ZN(n10684) );
  AOI22D1BWP30P140LVT U15341 ( .A1(i_data_bus[210]), .A2(n10828), .B1(
        i_data_bus[178]), .B2(n10829), .ZN(n10683) );
  ND2D1BWP30P140LVT U15342 ( .A1(n10684), .A2(n10683), .ZN(N10595) );
  AOI22D1BWP30P140LVT U15343 ( .A1(i_data_bus[131]), .A2(n10830), .B1(
        i_data_bus[195]), .B2(n10828), .ZN(n10686) );
  AOI22D1BWP30P140LVT U15344 ( .A1(i_data_bus[227]), .A2(n10831), .B1(
        i_data_bus[163]), .B2(n10829), .ZN(n10685) );
  ND2D1BWP30P140LVT U15345 ( .A1(n10686), .A2(n10685), .ZN(N10580) );
  AOI22D1BWP30P140LVT U15346 ( .A1(i_data_bus[134]), .A2(n10830), .B1(
        i_data_bus[198]), .B2(n10828), .ZN(n10688) );
  AOI22D1BWP30P140LVT U15347 ( .A1(i_data_bus[230]), .A2(n10831), .B1(
        i_data_bus[166]), .B2(n10829), .ZN(n10687) );
  ND2D1BWP30P140LVT U15348 ( .A1(n10688), .A2(n10687), .ZN(N10583) );
  AOI22D1BWP30P140LVT U15349 ( .A1(i_data_bus[137]), .A2(n10830), .B1(
        i_data_bus[169]), .B2(n10829), .ZN(n10690) );
  AOI22D1BWP30P140LVT U15350 ( .A1(i_data_bus[233]), .A2(n10831), .B1(
        i_data_bus[201]), .B2(n10828), .ZN(n10689) );
  ND2D1BWP30P140LVT U15351 ( .A1(n10690), .A2(n10689), .ZN(N10586) );
  NR3D0P7BWP30P140LVT U15352 ( .A1(i_cmd[143]), .A2(i_cmd[159]), .A3(
        i_cmd[151]), .ZN(n10922) );
  INR4D1BWP30P140LVT U15353 ( .A1(i_cmd[151]), .B1(i_cmd[135]), .B2(n10692), 
        .B3(n10926), .ZN(n10850) );
  AOI22D1BWP30P140LVT U15354 ( .A1(i_data_bus[512]), .A2(n10852), .B1(
        i_data_bus[576]), .B2(n10850), .ZN(n10699) );
  NR4D1BWP30P140LVT U15355 ( .A1(i_cmd[143]), .A2(n10694), .A3(n10693), .A4(
        n10695), .ZN(n10853) );
  NR4D1BWP30P140LVT U15356 ( .A1(i_cmd[159]), .A2(n10697), .A3(n10696), .A4(
        n10695), .ZN(n10851) );
  AOI22D1BWP30P140LVT U15357 ( .A1(i_data_bus[608]), .A2(n10853), .B1(
        i_data_bus[544]), .B2(n10851), .ZN(n10698) );
  ND2D1BWP30P140LVT U15358 ( .A1(n10699), .A2(n10698), .ZN(N10841) );
  AOI22D1BWP30P140LVT U15359 ( .A1(i_data_bus[525]), .A2(n10852), .B1(
        i_data_bus[589]), .B2(n10850), .ZN(n10701) );
  AOI22D1BWP30P140LVT U15360 ( .A1(i_data_bus[621]), .A2(n10853), .B1(
        i_data_bus[557]), .B2(n10851), .ZN(n10700) );
  ND2D1BWP30P140LVT U15361 ( .A1(n10701), .A2(n10700), .ZN(N10854) );
  AOI22D1BWP30P140LVT U15362 ( .A1(i_data_bus[521]), .A2(n10852), .B1(
        i_data_bus[617]), .B2(n10853), .ZN(n10703) );
  AOI22D1BWP30P140LVT U15363 ( .A1(i_data_bus[585]), .A2(n10850), .B1(
        i_data_bus[553]), .B2(n10851), .ZN(n10702) );
  ND2D1BWP30P140LVT U15364 ( .A1(n10703), .A2(n10702), .ZN(N10850) );
  AOI22D1BWP30P140LVT U15365 ( .A1(i_data_bus[530]), .A2(n10852), .B1(
        i_data_bus[562]), .B2(n10851), .ZN(n10705) );
  AOI22D1BWP30P140LVT U15366 ( .A1(i_data_bus[594]), .A2(n10850), .B1(
        i_data_bus[626]), .B2(n10853), .ZN(n10704) );
  ND2D1BWP30P140LVT U15367 ( .A1(n10705), .A2(n10704), .ZN(N10859) );
  AOI22D1BWP30P140LVT U15368 ( .A1(i_data_bus[514]), .A2(n10852), .B1(
        i_data_bus[546]), .B2(n10851), .ZN(n10707) );
  AOI22D1BWP30P140LVT U15369 ( .A1(i_data_bus[578]), .A2(n10850), .B1(
        i_data_bus[610]), .B2(n10853), .ZN(n10706) );
  ND2D1BWP30P140LVT U15370 ( .A1(n10707), .A2(n10706), .ZN(N10843) );
  AOI22D1BWP30P140LVT U15371 ( .A1(i_data_bus[518]), .A2(n10852), .B1(
        i_data_bus[614]), .B2(n10853), .ZN(n10709) );
  AOI22D1BWP30P140LVT U15372 ( .A1(i_data_bus[550]), .A2(n10851), .B1(
        i_data_bus[582]), .B2(n10850), .ZN(n10708) );
  ND2D1BWP30P140LVT U15373 ( .A1(n10709), .A2(n10708), .ZN(N10847) );
  AOI22D1BWP30P140LVT U15374 ( .A1(i_data_bus[123]), .A2(n10811), .B1(
        i_data_bus[91]), .B2(n10810), .ZN(n10711) );
  AOI22D1BWP30P140LVT U15375 ( .A1(i_data_bus[27]), .A2(n10812), .B1(
        i_data_bus[59]), .B2(n10813), .ZN(n10710) );
  ND2D1BWP30P140LVT U15376 ( .A1(n10711), .A2(n10710), .ZN(N10516) );
  AOI22D1BWP30P140LVT U15377 ( .A1(i_data_bus[79]), .A2(n10810), .B1(
        i_data_bus[47]), .B2(n10813), .ZN(n10713) );
  AOI22D1BWP30P140LVT U15378 ( .A1(i_data_bus[15]), .A2(n10812), .B1(
        i_data_bus[111]), .B2(n10811), .ZN(n10712) );
  ND2D1BWP30P140LVT U15379 ( .A1(n10713), .A2(n10712), .ZN(N10504) );
  AOI22D1BWP30P140LVT U15380 ( .A1(i_data_bus[78]), .A2(n10810), .B1(
        i_data_bus[110]), .B2(n10811), .ZN(n10715) );
  AOI22D1BWP30P140LVT U15381 ( .A1(i_data_bus[14]), .A2(n10812), .B1(
        i_data_bus[46]), .B2(n10813), .ZN(n10714) );
  ND2D1BWP30P140LVT U15382 ( .A1(n10715), .A2(n10714), .ZN(N10503) );
  AOI22D1BWP30P140LVT U15383 ( .A1(i_data_bus[117]), .A2(n10811), .B1(
        i_data_bus[53]), .B2(n10813), .ZN(n10717) );
  AOI22D1BWP30P140LVT U15384 ( .A1(i_data_bus[21]), .A2(n10812), .B1(
        i_data_bus[85]), .B2(n10810), .ZN(n10716) );
  ND2D1BWP30P140LVT U15385 ( .A1(n10717), .A2(n10716), .ZN(N10510) );
  AOI22D1BWP30P140LVT U15386 ( .A1(i_data_bus[104]), .A2(n10811), .B1(
        i_data_bus[72]), .B2(n10810), .ZN(n10719) );
  AOI22D1BWP30P140LVT U15387 ( .A1(i_data_bus[8]), .A2(n10812), .B1(
        i_data_bus[40]), .B2(n10813), .ZN(n10718) );
  ND2D1BWP30P140LVT U15388 ( .A1(n10719), .A2(n10718), .ZN(N10497) );
  AOI22D1BWP30P140LVT U15389 ( .A1(i_data_bus[77]), .A2(n10810), .B1(
        i_data_bus[109]), .B2(n10811), .ZN(n10721) );
  AOI22D1BWP30P140LVT U15390 ( .A1(i_data_bus[13]), .A2(n10812), .B1(
        i_data_bus[45]), .B2(n10813), .ZN(n10720) );
  ND2D1BWP30P140LVT U15391 ( .A1(n10721), .A2(n10720), .ZN(N10502) );
  AOI22D1BWP30P140LVT U15392 ( .A1(i_data_bus[112]), .A2(n10811), .B1(
        i_data_bus[80]), .B2(n10810), .ZN(n10723) );
  AOI22D1BWP30P140LVT U15393 ( .A1(i_data_bus[16]), .A2(n10812), .B1(
        i_data_bus[48]), .B2(n10813), .ZN(n10722) );
  ND2D1BWP30P140LVT U15394 ( .A1(n10723), .A2(n10722), .ZN(N10505) );
  AOI22D1BWP30P140LVT U15395 ( .A1(i_data_bus[36]), .A2(n10813), .B1(
        i_data_bus[100]), .B2(n10811), .ZN(n10725) );
  AOI22D1BWP30P140LVT U15396 ( .A1(i_data_bus[4]), .A2(n10812), .B1(
        i_data_bus[68]), .B2(n10810), .ZN(n10724) );
  ND2D1BWP30P140LVT U15397 ( .A1(n10725), .A2(n10724), .ZN(N10493) );
  AOI22D1BWP30P140LVT U15398 ( .A1(i_data_bus[102]), .A2(n10811), .B1(
        i_data_bus[70]), .B2(n10810), .ZN(n10727) );
  AOI22D1BWP30P140LVT U15399 ( .A1(i_data_bus[6]), .A2(n10812), .B1(
        i_data_bus[38]), .B2(n10813), .ZN(n10726) );
  ND2D1BWP30P140LVT U15400 ( .A1(n10727), .A2(n10726), .ZN(N10495) );
  AOI22D1BWP30P140LVT U15401 ( .A1(i_data_bus[34]), .A2(n10813), .B1(
        i_data_bus[98]), .B2(n10811), .ZN(n10729) );
  AOI22D1BWP30P140LVT U15402 ( .A1(i_data_bus[2]), .A2(n10812), .B1(
        i_data_bus[66]), .B2(n10810), .ZN(n10728) );
  ND2D1BWP30P140LVT U15403 ( .A1(n10729), .A2(n10728), .ZN(N10491) );
  AOI22D1BWP30P140LVT U15404 ( .A1(i_data_bus[74]), .A2(n10810), .B1(
        i_data_bus[106]), .B2(n10811), .ZN(n10731) );
  AOI22D1BWP30P140LVT U15405 ( .A1(i_data_bus[10]), .A2(n10812), .B1(
        i_data_bus[42]), .B2(n10813), .ZN(n10730) );
  ND2D1BWP30P140LVT U15406 ( .A1(n10731), .A2(n10730), .ZN(N10499) );
  AOI22D1BWP30P140LVT U15407 ( .A1(i_data_bus[32]), .A2(n10813), .B1(
        i_data_bus[96]), .B2(n10811), .ZN(n10733) );
  AOI22D1BWP30P140LVT U15408 ( .A1(i_data_bus[0]), .A2(n10812), .B1(
        i_data_bus[64]), .B2(n10810), .ZN(n10732) );
  ND2D1BWP30P140LVT U15409 ( .A1(n10733), .A2(n10732), .ZN(N10489) );
  AOI22D1BWP30P140LVT U15410 ( .A1(i_data_bus[50]), .A2(n10813), .B1(
        i_data_bus[82]), .B2(n10810), .ZN(n10735) );
  AOI22D1BWP30P140LVT U15411 ( .A1(i_data_bus[18]), .A2(n10812), .B1(
        i_data_bus[114]), .B2(n10811), .ZN(n10734) );
  ND2D1BWP30P140LVT U15412 ( .A1(n10735), .A2(n10734), .ZN(N10507) );
  AOI22D1BWP30P140LVT U15413 ( .A1(i_data_bus[187]), .A2(n10829), .B1(
        i_data_bus[219]), .B2(n10828), .ZN(n10737) );
  AOI22D1BWP30P140LVT U15414 ( .A1(i_data_bus[155]), .A2(n10830), .B1(
        i_data_bus[251]), .B2(n10831), .ZN(n10736) );
  ND2D1BWP30P140LVT U15415 ( .A1(n10737), .A2(n10736), .ZN(N10604) );
  AOI22D1BWP30P140LVT U15416 ( .A1(i_data_bus[247]), .A2(n10831), .B1(
        i_data_bus[183]), .B2(n10829), .ZN(n10739) );
  AOI22D1BWP30P140LVT U15417 ( .A1(i_data_bus[151]), .A2(n10830), .B1(
        i_data_bus[215]), .B2(n10828), .ZN(n10738) );
  ND2D1BWP30P140LVT U15418 ( .A1(n10739), .A2(n10738), .ZN(N10600) );
  AOI22D1BWP30P140LVT U15419 ( .A1(i_data_bus[234]), .A2(n10831), .B1(
        i_data_bus[202]), .B2(n10828), .ZN(n10741) );
  AOI22D1BWP30P140LVT U15420 ( .A1(i_data_bus[138]), .A2(n10830), .B1(
        i_data_bus[170]), .B2(n10829), .ZN(n10740) );
  ND2D1BWP30P140LVT U15421 ( .A1(n10741), .A2(n10740), .ZN(N10587) );
  AOI22D1BWP30P140LVT U15422 ( .A1(i_data_bus[172]), .A2(n10829), .B1(
        i_data_bus[204]), .B2(n10828), .ZN(n10743) );
  AOI22D1BWP30P140LVT U15423 ( .A1(i_data_bus[140]), .A2(n10830), .B1(
        i_data_bus[236]), .B2(n10831), .ZN(n10742) );
  ND2D1BWP30P140LVT U15424 ( .A1(n10743), .A2(n10742), .ZN(N10589) );
  AOI22D1BWP30P140LVT U15425 ( .A1(i_data_bus[239]), .A2(n10831), .B1(
        i_data_bus[207]), .B2(n10828), .ZN(n10745) );
  AOI22D1BWP30P140LVT U15426 ( .A1(i_data_bus[143]), .A2(n10830), .B1(
        i_data_bus[175]), .B2(n10829), .ZN(n10744) );
  ND2D1BWP30P140LVT U15427 ( .A1(n10745), .A2(n10744), .ZN(N10592) );
  AOI22D1BWP30P140LVT U15428 ( .A1(i_data_bus[232]), .A2(n10831), .B1(
        i_data_bus[200]), .B2(n10828), .ZN(n10747) );
  AOI22D1BWP30P140LVT U15429 ( .A1(i_data_bus[136]), .A2(n10830), .B1(
        i_data_bus[168]), .B2(n10829), .ZN(n10746) );
  ND2D1BWP30P140LVT U15430 ( .A1(n10747), .A2(n10746), .ZN(N10585) );
  AOI22D1BWP30P140LVT U15431 ( .A1(i_data_bus[171]), .A2(n10829), .B1(
        i_data_bus[203]), .B2(n10828), .ZN(n10749) );
  AOI22D1BWP30P140LVT U15432 ( .A1(i_data_bus[139]), .A2(n10830), .B1(
        i_data_bus[235]), .B2(n10831), .ZN(n10748) );
  ND2D1BWP30P140LVT U15433 ( .A1(n10749), .A2(n10748), .ZN(N10588) );
  AOI22D1BWP30P140LVT U15434 ( .A1(i_data_bus[240]), .A2(n10831), .B1(
        i_data_bus[208]), .B2(n10828), .ZN(n10751) );
  AOI22D1BWP30P140LVT U15435 ( .A1(i_data_bus[144]), .A2(n10830), .B1(
        i_data_bus[176]), .B2(n10829), .ZN(n10750) );
  ND2D1BWP30P140LVT U15436 ( .A1(n10751), .A2(n10750), .ZN(N10593) );
  AOI22D1BWP30P140LVT U15437 ( .A1(i_data_bus[253]), .A2(n10831), .B1(
        i_data_bus[189]), .B2(n10829), .ZN(n10753) );
  AOI22D1BWP30P140LVT U15438 ( .A1(i_data_bus[157]), .A2(n10830), .B1(
        i_data_bus[221]), .B2(n10828), .ZN(n10752) );
  ND2D1BWP30P140LVT U15439 ( .A1(n10753), .A2(n10752), .ZN(N10606) );
  AOI22D1BWP30P140LVT U15440 ( .A1(i_data_bus[570]), .A2(n10851), .B1(
        i_data_bus[602]), .B2(n10850), .ZN(n10755) );
  AOI22D1BWP30P140LVT U15441 ( .A1(i_data_bus[538]), .A2(n10852), .B1(
        i_data_bus[634]), .B2(n10853), .ZN(n10754) );
  ND2D1BWP30P140LVT U15442 ( .A1(n10755), .A2(n10754), .ZN(N10867) );
  AOI22D1BWP30P140LVT U15443 ( .A1(i_data_bus[581]), .A2(n10850), .B1(
        i_data_bus[613]), .B2(n10853), .ZN(n10757) );
  AOI22D1BWP30P140LVT U15444 ( .A1(i_data_bus[517]), .A2(n10852), .B1(
        i_data_bus[549]), .B2(n10851), .ZN(n10756) );
  ND2D1BWP30P140LVT U15445 ( .A1(n10757), .A2(n10756), .ZN(N10846) );
  AOI22D1BWP30P140LVT U15446 ( .A1(i_data_bus[566]), .A2(n10851), .B1(
        i_data_bus[598]), .B2(n10850), .ZN(n10759) );
  AOI22D1BWP30P140LVT U15447 ( .A1(i_data_bus[534]), .A2(n10852), .B1(
        i_data_bus[630]), .B2(n10853), .ZN(n10758) );
  ND2D1BWP30P140LVT U15448 ( .A1(n10759), .A2(n10758), .ZN(N10863) );
  AOI22D1BWP30P140LVT U15449 ( .A1(i_data_bus[629]), .A2(n10853), .B1(
        i_data_bus[597]), .B2(n10850), .ZN(n10761) );
  AOI22D1BWP30P140LVT U15450 ( .A1(i_data_bus[533]), .A2(n10852), .B1(
        i_data_bus[565]), .B2(n10851), .ZN(n10760) );
  ND2D1BWP30P140LVT U15451 ( .A1(n10761), .A2(n10760), .ZN(N10862) );
  AOI22D1BWP30P140LVT U15452 ( .A1(i_data_bus[561]), .A2(n10851), .B1(
        i_data_bus[625]), .B2(n10853), .ZN(n10763) );
  AOI22D1BWP30P140LVT U15453 ( .A1(i_data_bus[529]), .A2(n10852), .B1(
        i_data_bus[593]), .B2(n10850), .ZN(n10762) );
  ND2D1BWP30P140LVT U15454 ( .A1(n10763), .A2(n10762), .ZN(N10858) );
  AOI22D1BWP30P140LVT U15455 ( .A1(i_data_bus[627]), .A2(n10853), .B1(
        i_data_bus[563]), .B2(n10851), .ZN(n10765) );
  AOI22D1BWP30P140LVT U15456 ( .A1(i_data_bus[531]), .A2(n10852), .B1(
        i_data_bus[595]), .B2(n10850), .ZN(n10764) );
  ND2D1BWP30P140LVT U15457 ( .A1(n10765), .A2(n10764), .ZN(N10860) );
  AOI22D1BWP30P140LVT U15458 ( .A1(i_data_bus[548]), .A2(n10851), .B1(
        i_data_bus[580]), .B2(n10850), .ZN(n10767) );
  AOI22D1BWP30P140LVT U15459 ( .A1(i_data_bus[516]), .A2(n10852), .B1(
        i_data_bus[612]), .B2(n10853), .ZN(n10766) );
  ND2D1BWP30P140LVT U15460 ( .A1(n10767), .A2(n10766), .ZN(N10845) );
  AOI22D1BWP30P140LVT U15461 ( .A1(i_data_bus[628]), .A2(n10853), .B1(
        i_data_bus[596]), .B2(n10850), .ZN(n10769) );
  AOI22D1BWP30P140LVT U15462 ( .A1(i_data_bus[532]), .A2(n10852), .B1(
        i_data_bus[564]), .B2(n10851), .ZN(n10768) );
  ND2D1BWP30P140LVT U15463 ( .A1(n10769), .A2(n10768), .ZN(N10861) );
  AOI22D1BWP30P140LVT U15464 ( .A1(i_data_bus[571]), .A2(n10851), .B1(
        i_data_bus[603]), .B2(n10850), .ZN(n10771) );
  AOI22D1BWP30P140LVT U15465 ( .A1(i_data_bus[539]), .A2(n10852), .B1(
        i_data_bus[635]), .B2(n10853), .ZN(n10770) );
  ND2D1BWP30P140LVT U15466 ( .A1(n10771), .A2(n10770), .ZN(N10868) );
  AOI22D1BWP30P140LVT U15467 ( .A1(i_data_bus[93]), .A2(n10810), .B1(
        i_data_bus[29]), .B2(n10812), .ZN(n10773) );
  AOI22D1BWP30P140LVT U15468 ( .A1(i_data_bus[61]), .A2(n10813), .B1(
        i_data_bus[125]), .B2(n10811), .ZN(n10772) );
  ND2D1BWP30P140LVT U15469 ( .A1(n10773), .A2(n10772), .ZN(N10518) );
  AOI22D1BWP30P140LVT U15470 ( .A1(i_data_bus[164]), .A2(n10829), .B1(
        i_data_bus[132]), .B2(n10830), .ZN(n10775) );
  AOI22D1BWP30P140LVT U15471 ( .A1(i_data_bus[196]), .A2(n10828), .B1(
        i_data_bus[228]), .B2(n10831), .ZN(n10774) );
  ND2D1BWP30P140LVT U15472 ( .A1(n10775), .A2(n10774), .ZN(N10581) );
  AOI22D1BWP30P140LVT U15473 ( .A1(i_data_bus[229]), .A2(n10831), .B1(
        i_data_bus[133]), .B2(n10830), .ZN(n10777) );
  AOI22D1BWP30P140LVT U15474 ( .A1(i_data_bus[197]), .A2(n10828), .B1(
        i_data_bus[165]), .B2(n10829), .ZN(n10776) );
  ND2D1BWP30P140LVT U15475 ( .A1(n10777), .A2(n10776), .ZN(N10582) );
  AOI22D1BWP30P140LVT U15476 ( .A1(i_data_bus[254]), .A2(n10831), .B1(
        i_data_bus[158]), .B2(n10830), .ZN(n10779) );
  AOI22D1BWP30P140LVT U15477 ( .A1(i_data_bus[222]), .A2(n10828), .B1(
        i_data_bus[190]), .B2(n10829), .ZN(n10778) );
  ND2D1BWP30P140LVT U15478 ( .A1(n10779), .A2(n10778), .ZN(N10607) );
  AOI22D1BWP30P140LVT U15479 ( .A1(i_data_bus[225]), .A2(n10831), .B1(
        i_data_bus[129]), .B2(n10830), .ZN(n10781) );
  AOI22D1BWP30P140LVT U15480 ( .A1(i_data_bus[161]), .A2(n10829), .B1(
        i_data_bus[193]), .B2(n10828), .ZN(n10780) );
  ND2D1BWP30P140LVT U15481 ( .A1(n10781), .A2(n10780), .ZN(N10578) );
  AOI22D1BWP30P140LVT U15482 ( .A1(i_data_bus[179]), .A2(n10829), .B1(
        i_data_bus[147]), .B2(n10830), .ZN(n10783) );
  AOI22D1BWP30P140LVT U15483 ( .A1(i_data_bus[243]), .A2(n10831), .B1(
        i_data_bus[211]), .B2(n10828), .ZN(n10782) );
  ND2D1BWP30P140LVT U15484 ( .A1(n10783), .A2(n10782), .ZN(N10596) );
  AOI22D1BWP30P140LVT U15485 ( .A1(i_data_bus[188]), .A2(n10829), .B1(
        i_data_bus[156]), .B2(n10830), .ZN(n10785) );
  AOI22D1BWP30P140LVT U15486 ( .A1(i_data_bus[252]), .A2(n10831), .B1(
        i_data_bus[220]), .B2(n10828), .ZN(n10784) );
  ND2D1BWP30P140LVT U15487 ( .A1(n10785), .A2(n10784), .ZN(N10605) );
  AOI22D1BWP30P140LVT U15488 ( .A1(i_data_bus[587]), .A2(n10850), .B1(
        i_data_bus[523]), .B2(n10852), .ZN(n10787) );
  AOI22D1BWP30P140LVT U15489 ( .A1(i_data_bus[619]), .A2(n10853), .B1(
        i_data_bus[555]), .B2(n10851), .ZN(n10786) );
  ND2D1BWP30P140LVT U15490 ( .A1(n10787), .A2(n10786), .ZN(N10852) );
  AOI22D1BWP30P140LVT U15491 ( .A1(i_data_bus[638]), .A2(n10853), .B1(
        i_data_bus[542]), .B2(n10852), .ZN(n10789) );
  AOI22D1BWP30P140LVT U15492 ( .A1(i_data_bus[606]), .A2(n10850), .B1(
        i_data_bus[574]), .B2(n10851), .ZN(n10788) );
  ND2D1BWP30P140LVT U15493 ( .A1(n10789), .A2(n10788), .ZN(N10871) );
  AOI22D1BWP30P140LVT U15494 ( .A1(i_data_bus[568]), .A2(n10851), .B1(
        i_data_bus[536]), .B2(n10852), .ZN(n10791) );
  AOI22D1BWP30P140LVT U15495 ( .A1(i_data_bus[600]), .A2(n10850), .B1(
        i_data_bus[632]), .B2(n10853), .ZN(n10790) );
  ND2D1BWP30P140LVT U15496 ( .A1(n10791), .A2(n10790), .ZN(N10865) );
  AOI22D1BWP30P140LVT U15497 ( .A1(i_data_bus[583]), .A2(n10850), .B1(
        i_data_bus[519]), .B2(n10852), .ZN(n10793) );
  AOI22D1BWP30P140LVT U15498 ( .A1(i_data_bus[551]), .A2(n10851), .B1(
        i_data_bus[615]), .B2(n10853), .ZN(n10792) );
  ND2D1BWP30P140LVT U15499 ( .A1(n10793), .A2(n10792), .ZN(N10848) );
  AOI22D1BWP30P140LVT U15500 ( .A1(i_data_bus[579]), .A2(n10850), .B1(
        i_data_bus[515]), .B2(n10852), .ZN(n10795) );
  AOI22D1BWP30P140LVT U15501 ( .A1(i_data_bus[547]), .A2(n10851), .B1(
        i_data_bus[611]), .B2(n10853), .ZN(n10794) );
  ND2D1BWP30P140LVT U15502 ( .A1(n10795), .A2(n10794), .ZN(N10844) );
  AOI22D1BWP30P140LVT U15503 ( .A1(i_data_bus[590]), .A2(n10850), .B1(
        i_data_bus[526]), .B2(n10852), .ZN(n10797) );
  AOI22D1BWP30P140LVT U15504 ( .A1(i_data_bus[558]), .A2(n10851), .B1(
        i_data_bus[622]), .B2(n10853), .ZN(n10796) );
  ND2D1BWP30P140LVT U15505 ( .A1(n10797), .A2(n10796), .ZN(N10855) );
  AOI22D1BWP30P140LVT U15506 ( .A1(i_data_bus[631]), .A2(n10853), .B1(
        i_data_bus[535]), .B2(n10852), .ZN(n10799) );
  AOI22D1BWP30P140LVT U15507 ( .A1(i_data_bus[567]), .A2(n10851), .B1(
        i_data_bus[599]), .B2(n10850), .ZN(n10798) );
  ND2D1BWP30P140LVT U15508 ( .A1(n10799), .A2(n10798), .ZN(N10864) );
  AOI22D1BWP30P140LVT U15509 ( .A1(i_data_bus[609]), .A2(n10853), .B1(
        i_data_bus[513]), .B2(n10852), .ZN(n10801) );
  AOI22D1BWP30P140LVT U15510 ( .A1(i_data_bus[545]), .A2(n10851), .B1(
        i_data_bus[577]), .B2(n10850), .ZN(n10800) );
  ND2D1BWP30P140LVT U15511 ( .A1(n10801), .A2(n10800), .ZN(N10842) );
  AOI22D1BWP30P140LVT U15512 ( .A1(i_data_bus[108]), .A2(n10811), .B1(
        i_data_bus[44]), .B2(n10813), .ZN(n10803) );
  AOI22D1BWP30P140LVT U15513 ( .A1(i_data_bus[76]), .A2(n10810), .B1(
        i_data_bus[12]), .B2(n10812), .ZN(n10802) );
  ND2D1BWP30P140LVT U15514 ( .A1(n10803), .A2(n10802), .ZN(N10501) );
  AOI22D1BWP30P140LVT U15515 ( .A1(i_data_bus[95]), .A2(n10810), .B1(
        i_data_bus[63]), .B2(n10813), .ZN(n10805) );
  AOI22D1BWP30P140LVT U15516 ( .A1(i_data_bus[127]), .A2(n10811), .B1(
        i_data_bus[31]), .B2(n10812), .ZN(n10804) );
  ND2D1BWP30P140LVT U15517 ( .A1(n10805), .A2(n10804), .ZN(N10520) );
  AOI22D1BWP30P140LVT U15518 ( .A1(i_data_bus[118]), .A2(n10811), .B1(
        i_data_bus[54]), .B2(n10813), .ZN(n10807) );
  AOI22D1BWP30P140LVT U15519 ( .A1(i_data_bus[86]), .A2(n10810), .B1(
        i_data_bus[22]), .B2(n10812), .ZN(n10806) );
  ND2D1BWP30P140LVT U15520 ( .A1(n10807), .A2(n10806), .ZN(N10511) );
  AOI22D1BWP30P140LVT U15521 ( .A1(i_data_bus[55]), .A2(n10813), .B1(
        i_data_bus[119]), .B2(n10811), .ZN(n10809) );
  AOI22D1BWP30P140LVT U15522 ( .A1(i_data_bus[87]), .A2(n10810), .B1(
        i_data_bus[23]), .B2(n10812), .ZN(n10808) );
  ND2D1BWP30P140LVT U15523 ( .A1(n10809), .A2(n10808), .ZN(N10512) );
  AOI22D1BWP30P140LVT U15524 ( .A1(i_data_bus[99]), .A2(n10811), .B1(
        i_data_bus[67]), .B2(n10810), .ZN(n10815) );
  AOI22D1BWP30P140LVT U15525 ( .A1(i_data_bus[35]), .A2(n10813), .B1(
        i_data_bus[3]), .B2(n10812), .ZN(n10814) );
  ND2D1BWP30P140LVT U15526 ( .A1(n10815), .A2(n10814), .ZN(N10492) );
  AOI22D1BWP30P140LVT U15527 ( .A1(i_data_bus[255]), .A2(n10831), .B1(
        i_data_bus[191]), .B2(n10829), .ZN(n10817) );
  AOI22D1BWP30P140LVT U15528 ( .A1(i_data_bus[223]), .A2(n10828), .B1(
        i_data_bus[159]), .B2(n10830), .ZN(n10816) );
  ND2D1BWP30P140LVT U15529 ( .A1(n10817), .A2(n10816), .ZN(N10608) );
  AOI22D1BWP30P140LVT U15530 ( .A1(i_data_bus[231]), .A2(n10831), .B1(
        i_data_bus[167]), .B2(n10829), .ZN(n10819) );
  AOI22D1BWP30P140LVT U15531 ( .A1(i_data_bus[199]), .A2(n10828), .B1(
        i_data_bus[135]), .B2(n10830), .ZN(n10818) );
  ND2D1BWP30P140LVT U15532 ( .A1(n10819), .A2(n10818), .ZN(N10584) );
  AOI22D1BWP30P140LVT U15533 ( .A1(i_data_bus[173]), .A2(n10829), .B1(
        i_data_bus[237]), .B2(n10831), .ZN(n10821) );
  AOI22D1BWP30P140LVT U15534 ( .A1(i_data_bus[205]), .A2(n10828), .B1(
        i_data_bus[141]), .B2(n10830), .ZN(n10820) );
  ND2D1BWP30P140LVT U15535 ( .A1(n10821), .A2(n10820), .ZN(N10590) );
  AOI22D1BWP30P140LVT U15536 ( .A1(i_data_bus[217]), .A2(n10828), .B1(
        i_data_bus[185]), .B2(n10829), .ZN(n10823) );
  AOI22D1BWP30P140LVT U15537 ( .A1(i_data_bus[249]), .A2(n10831), .B1(
        i_data_bus[153]), .B2(n10830), .ZN(n10822) );
  ND2D1BWP30P140LVT U15538 ( .A1(n10823), .A2(n10822), .ZN(N10602) );
  AOI22D1BWP30P140LVT U15539 ( .A1(i_data_bus[162]), .A2(n10829), .B1(
        i_data_bus[226]), .B2(n10831), .ZN(n10825) );
  AOI22D1BWP30P140LVT U15540 ( .A1(i_data_bus[194]), .A2(n10828), .B1(
        i_data_bus[130]), .B2(n10830), .ZN(n10824) );
  ND2D1BWP30P140LVT U15541 ( .A1(n10825), .A2(n10824), .ZN(N10579) );
  AOI22D1BWP30P140LVT U15542 ( .A1(i_data_bus[244]), .A2(n10831), .B1(
        i_data_bus[180]), .B2(n10829), .ZN(n10827) );
  AOI22D1BWP30P140LVT U15543 ( .A1(i_data_bus[212]), .A2(n10828), .B1(
        i_data_bus[148]), .B2(n10830), .ZN(n10826) );
  ND2D1BWP30P140LVT U15544 ( .A1(n10827), .A2(n10826), .ZN(N10597) );
  AOI22D1BWP30P140LVT U15545 ( .A1(i_data_bus[160]), .A2(n10829), .B1(
        i_data_bus[192]), .B2(n10828), .ZN(n10833) );
  AOI22D1BWP30P140LVT U15546 ( .A1(i_data_bus[224]), .A2(n10831), .B1(
        i_data_bus[128]), .B2(n10830), .ZN(n10832) );
  ND2D1BWP30P140LVT U15547 ( .A1(n10833), .A2(n10832), .ZN(N10577) );
  AOI22D1BWP30P140LVT U15548 ( .A1(i_data_bus[618]), .A2(n10853), .B1(
        i_data_bus[554]), .B2(n10851), .ZN(n10835) );
  AOI22D1BWP30P140LVT U15549 ( .A1(i_data_bus[586]), .A2(n10850), .B1(
        i_data_bus[522]), .B2(n10852), .ZN(n10834) );
  ND2D1BWP30P140LVT U15550 ( .A1(n10835), .A2(n10834), .ZN(N10851) );
  AOI22D1BWP30P140LVT U15551 ( .A1(i_data_bus[560]), .A2(n10851), .B1(
        i_data_bus[592]), .B2(n10850), .ZN(n10837) );
  AOI22D1BWP30P140LVT U15552 ( .A1(i_data_bus[624]), .A2(n10853), .B1(
        i_data_bus[528]), .B2(n10852), .ZN(n10836) );
  ND2D1BWP30P140LVT U15553 ( .A1(n10837), .A2(n10836), .ZN(N10857) );
  AOI22D1BWP30P140LVT U15554 ( .A1(i_data_bus[556]), .A2(n10851), .B1(
        i_data_bus[588]), .B2(n10850), .ZN(n10839) );
  AOI22D1BWP30P140LVT U15555 ( .A1(i_data_bus[620]), .A2(n10853), .B1(
        i_data_bus[524]), .B2(n10852), .ZN(n10838) );
  ND2D1BWP30P140LVT U15556 ( .A1(n10839), .A2(n10838), .ZN(N10853) );
  AOI22D1BWP30P140LVT U15557 ( .A1(i_data_bus[623]), .A2(n10853), .B1(
        i_data_bus[591]), .B2(n10850), .ZN(n10841) );
  AOI22D1BWP30P140LVT U15558 ( .A1(i_data_bus[559]), .A2(n10851), .B1(
        i_data_bus[527]), .B2(n10852), .ZN(n10840) );
  ND2D1BWP30P140LVT U15559 ( .A1(n10841), .A2(n10840), .ZN(N10856) );
  AOI22D1BWP30P140LVT U15560 ( .A1(i_data_bus[584]), .A2(n10850), .B1(
        i_data_bus[552]), .B2(n10851), .ZN(n10843) );
  AOI22D1BWP30P140LVT U15561 ( .A1(i_data_bus[616]), .A2(n10853), .B1(
        i_data_bus[520]), .B2(n10852), .ZN(n10842) );
  ND2D1BWP30P140LVT U15562 ( .A1(n10843), .A2(n10842), .ZN(N10849) );
  AOI22D1BWP30P140LVT U15563 ( .A1(i_data_bus[604]), .A2(n10850), .B1(
        i_data_bus[636]), .B2(n10853), .ZN(n10845) );
  AOI22D1BWP30P140LVT U15564 ( .A1(i_data_bus[572]), .A2(n10851), .B1(
        i_data_bus[540]), .B2(n10852), .ZN(n10844) );
  ND2D1BWP30P140LVT U15565 ( .A1(n10845), .A2(n10844), .ZN(N10869) );
  AOI22D1BWP30P140LVT U15566 ( .A1(i_data_bus[637]), .A2(n10853), .B1(
        i_data_bus[605]), .B2(n10850), .ZN(n10847) );
  AOI22D1BWP30P140LVT U15567 ( .A1(i_data_bus[573]), .A2(n10851), .B1(
        i_data_bus[541]), .B2(n10852), .ZN(n10846) );
  ND2D1BWP30P140LVT U15568 ( .A1(n10847), .A2(n10846), .ZN(N10870) );
  AOI22D1BWP30P140LVT U15569 ( .A1(i_data_bus[607]), .A2(n10850), .B1(
        i_data_bus[575]), .B2(n10851), .ZN(n10849) );
  AOI22D1BWP30P140LVT U15570 ( .A1(i_data_bus[639]), .A2(n10853), .B1(
        i_data_bus[543]), .B2(n10852), .ZN(n10848) );
  ND2D1BWP30P140LVT U15571 ( .A1(n10849), .A2(n10848), .ZN(N10872) );
  AOI22D1BWP30P140LVT U15572 ( .A1(i_data_bus[569]), .A2(n10851), .B1(
        i_data_bus[601]), .B2(n10850), .ZN(n10855) );
  AOI22D1BWP30P140LVT U15573 ( .A1(i_data_bus[633]), .A2(n10853), .B1(
        i_data_bus[537]), .B2(n10852), .ZN(n10854) );
  ND2D1BWP30P140LVT U15574 ( .A1(n10855), .A2(n10854), .ZN(N10866) );
  NR4D0BWP30P140LVT U15575 ( .A1(inner_first_stage_valid_reg[10]), .A2(
        inner_first_stage_valid_reg[11]), .A3(inner_first_stage_valid_reg[13]), 
        .A4(inner_first_stage_valid_reg[9]), .ZN(n10862) );
  INR3D2BWP30P140LVT U15576 ( .A1(inner_first_stage_valid_reg[15]), .B1(
        inner_first_stage_valid_reg[14]), .B2(n10857), .ZN(n11481) );
  INR3D2BWP30P140LVT U15577 ( .A1(inner_first_stage_valid_reg[14]), .B1(
        inner_first_stage_valid_reg[15]), .B2(n10857), .ZN(n11480) );
  NR2D1BWP30P140LVT U15578 ( .A1(inner_first_stage_valid_reg[13]), .A2(
        inner_first_stage_valid_reg[9]), .ZN(n10858) );
  NR3D0P7BWP30P140LVT U15579 ( .A1(inner_first_stage_valid_reg[8]), .A2(
        inner_first_stage_valid_reg[14]), .A3(inner_first_stage_valid_reg[15]), 
        .ZN(n10863) );
  INR3D0BWP30P140LVT U15580 ( .A1(n10863), .B1(inner_first_stage_valid_reg[12]), .B2(n11173), .ZN(n10859) );
  INR3D2BWP30P140LVT U15581 ( .A1(inner_first_stage_valid_reg[11]), .B1(
        inner_first_stage_valid_reg[10]), .B2(n10865), .ZN(n11483) );
  NR2D1BWP30P140LVT U15582 ( .A1(inner_first_stage_valid_reg[10]), .A2(
        inner_first_stage_valid_reg[11]), .ZN(n10860) );
  INR3D2BWP30P140LVT U15583 ( .A1(inner_first_stage_valid_reg[13]), .B1(
        inner_first_stage_valid_reg[9]), .B2(n10864), .ZN(n11482) );
  NR4D0BWP30P140LVT U15584 ( .A1(n11481), .A2(n11480), .A3(n11483), .A4(n11482), .ZN(n10867) );
  INR4D1BWP30P140LVT U15585 ( .A1(inner_first_stage_valid_reg[8]), .B1(
        inner_first_stage_valid_reg[15]), .B2(inner_first_stage_valid_reg[14]), 
        .B3(n10861), .ZN(n11477) );
  INR3D2BWP30P140LVT U15586 ( .A1(inner_first_stage_valid_reg[9]), .B1(
        inner_first_stage_valid_reg[13]), .B2(n10864), .ZN(n11479) );
  INR3D2BWP30P140LVT U15587 ( .A1(inner_first_stage_valid_reg[10]), .B1(
        inner_first_stage_valid_reg[11]), .B2(n10865), .ZN(n11478) );
  NR4D0BWP30P140LVT U15588 ( .A1(n11477), .A2(n11476), .A3(n11479), .A4(n11478), .ZN(n10866) );
  INVD1BWP30P140LVT U15589 ( .I(inner_first_stage_valid_reg[38]), .ZN(n10870)
         );
  NR4D0BWP30P140LVT U15590 ( .A1(inner_first_stage_valid_reg[34]), .A2(
        inner_first_stage_valid_reg[35]), .A3(inner_first_stage_valid_reg[32]), 
        .A4(n10878), .ZN(n10875) );
  INVD1BWP30P140LVT U15591 ( .I(inner_first_stage_valid_reg[36]), .ZN(n10874)
         );
  ND3D1BWP30P140LVT U15592 ( .A1(n12302), .A2(n10875), .A3(n10874), .ZN(n10868) );
  ND3D1BWP30P140LVT U15593 ( .A1(n10870), .A2(n12303), .A3(n10869), .ZN(n10873) );
  NR4D0BWP30P140LVT U15594 ( .A1(inner_first_stage_valid_reg[34]), .A2(
        inner_first_stage_valid_reg[36]), .A3(inner_first_stage_valid_reg[35]), 
        .A4(n10873), .ZN(n10879) );
  INR3D2BWP30P140LVT U15595 ( .A1(inner_first_stage_valid_reg[37]), .B1(
        inner_first_stage_valid_reg[33]), .B2(n10871), .ZN(n11891) );
  INR3D2BWP30P140LVT U15596 ( .A1(inner_first_stage_valid_reg[33]), .B1(
        inner_first_stage_valid_reg[37]), .B2(n10871), .ZN(n11890) );
  NR4D0BWP30P140LVT U15597 ( .A1(n11889), .A2(n11888), .A3(n11891), .A4(n11890), .ZN(n10881) );
  NR4D0BWP30P140LVT U15598 ( .A1(inner_first_stage_valid_reg[38]), .A2(
        inner_first_stage_valid_reg[36]), .A3(inner_first_stage_valid_reg[39]), 
        .A4(n10878), .ZN(n10872) );
  INR4D1BWP30P140LVT U15599 ( .A1(inner_first_stage_valid_reg[34]), .B1(
        inner_first_stage_valid_reg[32]), .B2(inner_first_stage_valid_reg[35]), 
        .B3(n10876), .ZN(n11885) );
  INR4D1BWP30P140LVT U15600 ( .A1(inner_first_stage_valid_reg[35]), .B1(
        inner_first_stage_valid_reg[34]), .B2(inner_first_stage_valid_reg[32]), 
        .B3(n10876), .ZN(n11884) );
  INR3D2BWP30P140LVT U15601 ( .A1(n10879), .B1(n10878), .B2(n10877), .ZN(
        n11886) );
  NR4D0BWP30P140LVT U15602 ( .A1(n11885), .A2(n11887), .A3(n11884), .A4(n11886), .ZN(n10880) );
  NR3D0P7BWP30P140LVT U15603 ( .A1(inner_first_stage_valid_reg[17]), .A2(
        inner_first_stage_valid_reg[18]), .A3(inner_first_stage_valid_reg[19]), 
        .ZN(n10887) );
  NR2D1BWP30P140LVT U15604 ( .A1(inner_first_stage_valid_reg[21]), .A2(
        inner_first_stage_valid_reg[16]), .ZN(n10882) );
  INR3D2BWP30P140LVT U15605 ( .A1(inner_first_stage_valid_reg[22]), .B1(
        inner_first_stage_valid_reg[23]), .B2(n10883), .ZN(n11617) );
  INR3D2BWP30P140LVT U15606 ( .A1(inner_first_stage_valid_reg[23]), .B1(
        inner_first_stage_valid_reg[22]), .B2(n10883), .ZN(n11619) );
  NR3D0P7BWP30P140LVT U15607 ( .A1(inner_first_stage_valid_reg[16]), .A2(
        inner_first_stage_valid_reg[20]), .A3(n10892), .ZN(n10886) );
  NR2D1BWP30P140LVT U15608 ( .A1(inner_first_stage_valid_reg[17]), .A2(
        inner_first_stage_valid_reg[21]), .ZN(n10884) );
  INR3D2BWP30P140LVT U15609 ( .A1(inner_first_stage_valid_reg[18]), .B1(
        inner_first_stage_valid_reg[19]), .B2(n10885), .ZN(n11616) );
  INR3D2BWP30P140LVT U15610 ( .A1(inner_first_stage_valid_reg[19]), .B1(
        inner_first_stage_valid_reg[18]), .B2(n10885), .ZN(n11618) );
  NR4D0BWP30P140LVT U15611 ( .A1(n11617), .A2(n11619), .A3(n11616), .A4(n11618), .ZN(n10895) );
  NR2D1BWP30P140LVT U15612 ( .A1(inner_first_stage_valid_reg[18]), .A2(
        inner_first_stage_valid_reg[19]), .ZN(n10890) );
  ND3D1BWP30P140LVT U15613 ( .A1(n10890), .A2(n10889), .A3(n10888), .ZN(n10893) );
  INR4D1BWP30P140LVT U15614 ( .A1(inner_first_stage_valid_reg[16]), .B1(
        inner_first_stage_valid_reg[17]), .B2(inner_first_stage_valid_reg[21]), 
        .B3(n10893), .ZN(n11613) );
  INR3D2BWP30P140LVT U15615 ( .A1(inner_first_stage_valid_reg[20]), .B1(n10892), .B2(n10891), .ZN(n11614) );
  INR4D1BWP30P140LVT U15616 ( .A1(inner_first_stage_valid_reg[17]), .B1(
        inner_first_stage_valid_reg[16]), .B2(inner_first_stage_valid_reg[21]), 
        .B3(n10893), .ZN(n11612) );
  NR4D0BWP30P140LVT U15617 ( .A1(n11615), .A2(n11613), .A3(n11614), .A4(n11612), .ZN(n10894) );
  NR3D0P7BWP30P140LVT U15618 ( .A1(inner_first_stage_valid_reg[46]), .A2(
        inner_first_stage_valid_reg[47]), .A3(n11173), .ZN(n10900) );
  NR2D1BWP30P140LVT U15619 ( .A1(inner_first_stage_valid_reg[41]), .A2(
        inner_first_stage_valid_reg[45]), .ZN(n10896) );
  IND4D1BWP30P140LVT U15620 ( .A1(inner_first_stage_valid_reg[44]), .B1(n10900), .B2(n10896), .B3(n10907), .ZN(n10897) );
  INR3D2BWP30P140LVT U15621 ( .A1(inner_first_stage_valid_reg[43]), .B1(
        inner_first_stage_valid_reg[42]), .B2(n10897), .ZN(n12025) );
  INR3D2BWP30P140LVT U15622 ( .A1(inner_first_stage_valid_reg[42]), .B1(
        inner_first_stage_valid_reg[43]), .B2(n10897), .ZN(n12024) );
  INVD1BWP30P140LVT U15623 ( .I(inner_first_stage_valid_reg[41]), .ZN(n10905)
         );
  NR4D0BWP30P140LVT U15624 ( .A1(inner_first_stage_valid_reg[42]), .A2(
        inner_first_stage_valid_reg[43]), .A3(inner_first_stage_valid_reg[45]), 
        .A4(n10898), .ZN(n10901) );
  INR3D2BWP30P140LVT U15625 ( .A1(inner_first_stage_valid_reg[47]), .B1(
        inner_first_stage_valid_reg[46]), .B2(n10899), .ZN(n12027) );
  INR3D2BWP30P140LVT U15626 ( .A1(inner_first_stage_valid_reg[46]), .B1(
        inner_first_stage_valid_reg[47]), .B2(n10899), .ZN(n12026) );
  NR4D0BWP30P140LVT U15627 ( .A1(n12025), .A2(n12024), .A3(n12027), .A4(n12026), .ZN(n10909) );
  ND3D1BWP30P140LVT U15628 ( .A1(n10904), .A2(n10903), .A3(n10902), .ZN(n10906) );
  NR4D1BWP30P140LVT U15629 ( .A1(inner_first_stage_valid_reg[45]), .A2(
        inner_first_stage_valid_reg[40]), .A3(n10905), .A4(n10906), .ZN(n12023) );
  INR4D1BWP30P140LVT U15630 ( .A1(inner_first_stage_valid_reg[45]), .B1(
        inner_first_stage_valid_reg[41]), .B2(inner_first_stage_valid_reg[40]), 
        .B3(n10906), .ZN(n12020) );
  NR4D1BWP30P140LVT U15631 ( .A1(inner_first_stage_valid_reg[41]), .A2(
        inner_first_stage_valid_reg[45]), .A3(n10907), .A4(n10906), .ZN(n12022) );
  NR4D0BWP30P140LVT U15632 ( .A1(n12021), .A2(n12023), .A3(n12020), .A4(n12022), .ZN(n10908) );
  AOI211D1BWP30P140LVT U15633 ( .A1(i_cmd[255]), .A2(i_cmd[239]), .B(
        i_cmd[231]), .C(n10910), .ZN(n10911) );
  INR2D1BWP30P140LVT U15634 ( .A1(n10912), .B1(n10911), .ZN(n10913) );
  AOI211D1BWP30P140LVT U15635 ( .A1(i_cmd[247]), .A2(n10914), .B(n10913), .C(
        n11181), .ZN(N11104) );
  AOI211D1BWP30P140LVT U15636 ( .A1(i_cmd[215]), .A2(n10916), .B(i_cmd[199]), 
        .C(n10915), .ZN(n10917) );
  OAI21D1BWP30P140LVT U15637 ( .A1(n10919), .A2(n10918), .B(n10917), .ZN(
        n10920) );
  AOI21D1BWP30P140LVT U15638 ( .A1(n10921), .A2(n10920), .B(n11173), .ZN(
        N11016) );
  AOI211D1BWP30P140LVT U15639 ( .A1(i_cmd[159]), .A2(i_cmd[143]), .B(
        i_cmd[135]), .C(n10922), .ZN(n10923) );
  INR2D1BWP30P140LVT U15640 ( .A1(n10924), .B1(n10923), .ZN(n10925) );
  AOI211D1BWP30P140LVT U15641 ( .A1(i_cmd[151]), .A2(n10926), .B(n10925), .C(
        n11181), .ZN(N10840) );
  AOI211D1BWP30P140LVT U15642 ( .A1(i_cmd[87]), .A2(n10928), .B(i_cmd[71]), 
        .C(n10927), .ZN(n10929) );
  OAI21D1BWP30P140LVT U15643 ( .A1(n10931), .A2(n10930), .B(n10929), .ZN(
        n10932) );
  AOI21D1BWP30P140LVT U15644 ( .A1(n10933), .A2(n10932), .B(n11173), .ZN(
        N10664) );
  AOI211D1BWP30P140LVT U15645 ( .A1(i_cmd[31]), .A2(i_cmd[15]), .B(n10934), 
        .C(i_cmd[7]), .ZN(n10935) );
  INR2D1BWP30P140LVT U15646 ( .A1(n10936), .B1(n10935), .ZN(n10937) );
  AOI211D1BWP30P140LVT U15647 ( .A1(i_cmd[23]), .A2(n10938), .B(n10937), .C(
        n11181), .ZN(N10488) );
  AOI211D1BWP30P140LVT U15648 ( .A1(i_cmd[254]), .A2(i_cmd[238]), .B(n10939), 
        .C(i_cmd[230]), .ZN(n10940) );
  INR2D1BWP30P140LVT U15649 ( .A1(n10941), .B1(n10940), .ZN(n10942) );
  AOI211D1BWP30P140LVT U15650 ( .A1(i_cmd[246]), .A2(n10943), .B(n10942), .C(
        n11181), .ZN(N10254) );
  AOI211D1BWP30P140LVT U15651 ( .A1(i_cmd[190]), .A2(i_cmd[174]), .B(
        i_cmd[166]), .C(n10944), .ZN(n10945) );
  INR2D1BWP30P140LVT U15652 ( .A1(n10946), .B1(n10945), .ZN(n10947) );
  AOI211D1BWP30P140LVT U15653 ( .A1(i_cmd[182]), .A2(n10948), .B(n10947), .C(
        n11181), .ZN(N9822) );
  AOI211D1BWP30P140LVT U15654 ( .A1(i_cmd[150]), .A2(n10950), .B(i_cmd[134]), 
        .C(n10949), .ZN(n10951) );
  OAI21D1BWP30P140LVT U15655 ( .A1(n10953), .A2(n10952), .B(n10951), .ZN(
        n10954) );
  AOI21D1BWP30P140LVT U15656 ( .A1(n10955), .A2(n10954), .B(n11181), .ZN(N9606) );
  AOI211D1BWP30P140LVT U15657 ( .A1(i_cmd[86]), .A2(n10957), .B(i_cmd[70]), 
        .C(n10956), .ZN(n10958) );
  OAI21D1BWP30P140LVT U15658 ( .A1(n10960), .A2(n10959), .B(n10958), .ZN(
        n10961) );
  AOI21D1BWP30P140LVT U15659 ( .A1(n10962), .A2(n10961), .B(n11181), .ZN(N9174) );
  AOI211D1BWP30P140LVT U15660 ( .A1(i_cmd[30]), .A2(i_cmd[14]), .B(i_cmd[6]), 
        .C(n10963), .ZN(n10964) );
  INR2D1BWP30P140LVT U15661 ( .A1(n10965), .B1(n10964), .ZN(n10966) );
  AOI211D1BWP30P140LVT U15662 ( .A1(i_cmd[22]), .A2(n10967), .B(n10966), .C(
        n11181), .ZN(N8742) );
  AOI211D1BWP30P140LVT U15663 ( .A1(i_cmd[237]), .A2(i_cmd[253]), .B(
        i_cmd[229]), .C(n10968), .ZN(n10969) );
  INR2D1BWP30P140LVT U15664 ( .A1(n10970), .B1(n10969), .ZN(n10971) );
  AOI211D1BWP30P140LVT U15665 ( .A1(i_cmd[245]), .A2(n10972), .B(n10971), .C(
        n11181), .ZN(N8380) );
  AOI211D1BWP30P140LVT U15666 ( .A1(i_cmd[221]), .A2(i_cmd[205]), .B(
        i_cmd[197]), .C(n10973), .ZN(n10974) );
  INR2D1BWP30P140LVT U15667 ( .A1(n10975), .B1(n10974), .ZN(n10976) );
  AOI211D1BWP30P140LVT U15668 ( .A1(i_cmd[213]), .A2(n10977), .B(n10976), .C(
        n11181), .ZN(N8292) );
  AOI211D1BWP30P140LVT U15669 ( .A1(i_cmd[181]), .A2(n10979), .B(i_cmd[165]), 
        .C(n10978), .ZN(n10980) );
  OAI21D1BWP30P140LVT U15670 ( .A1(n10982), .A2(n10981), .B(n10980), .ZN(
        n10983) );
  AOI21D1BWP30P140LVT U15671 ( .A1(n10984), .A2(n10983), .B(n11181), .ZN(N8204) );
  AOI211D1BWP30P140LVT U15672 ( .A1(i_cmd[157]), .A2(i_cmd[141]), .B(
        i_cmd[133]), .C(n10985), .ZN(n10986) );
  INR2D1BWP30P140LVT U15673 ( .A1(n10987), .B1(n10986), .ZN(n10988) );
  AOI211D1BWP30P140LVT U15674 ( .A1(i_cmd[149]), .A2(n10989), .B(n10988), .C(
        n11181), .ZN(N8116) );
  AOI211D1BWP30P140LVT U15675 ( .A1(i_cmd[117]), .A2(n10991), .B(i_cmd[101]), 
        .C(n10990), .ZN(n10992) );
  OAI21D1BWP30P140LVT U15676 ( .A1(n10994), .A2(n10993), .B(n10992), .ZN(
        n10995) );
  AOI21D1BWP30P140LVT U15677 ( .A1(n10996), .A2(n10995), .B(n11057), .ZN(N8028) );
  AOI211D1BWP30P140LVT U15678 ( .A1(i_cmd[85]), .A2(n10998), .B(i_cmd[69]), 
        .C(n10997), .ZN(n10999) );
  OAI21D1BWP30P140LVT U15679 ( .A1(n11001), .A2(n11000), .B(n10999), .ZN(
        n11002) );
  AOI21D1BWP30P140LVT U15680 ( .A1(n11003), .A2(n11002), .B(n11181), .ZN(N7940) );
  AOI211D1BWP30P140LVT U15681 ( .A1(i_cmd[61]), .A2(i_cmd[45]), .B(i_cmd[37]), 
        .C(n11004), .ZN(n11005) );
  INR2D1BWP30P140LVT U15682 ( .A1(n11006), .B1(n11005), .ZN(n11007) );
  AOI211D1BWP30P140LVT U15683 ( .A1(i_cmd[53]), .A2(n11008), .B(n11007), .C(
        n11181), .ZN(N7852) );
  AOI211D1BWP30P140LVT U15684 ( .A1(i_cmd[29]), .A2(i_cmd[13]), .B(i_cmd[5]), 
        .C(n11009), .ZN(n11010) );
  INR2D1BWP30P140LVT U15685 ( .A1(n11011), .B1(n11010), .ZN(n11012) );
  AOI211D1BWP30P140LVT U15686 ( .A1(i_cmd[21]), .A2(n11013), .B(n11012), .C(
        n11181), .ZN(N7764) );
  AOI211D1BWP30P140LVT U15687 ( .A1(i_cmd[220]), .A2(i_cmd[204]), .B(n11014), 
        .C(i_cmd[196]), .ZN(n11015) );
  INR2D1BWP30P140LVT U15688 ( .A1(n11016), .B1(n11015), .ZN(n11017) );
  AOI211D1BWP30P140LVT U15689 ( .A1(i_cmd[212]), .A2(n11018), .B(n11017), .C(
        n11181), .ZN(N7314) );
  AOI211D1BWP30P140LVT U15690 ( .A1(i_cmd[180]), .A2(n11020), .B(i_cmd[164]), 
        .C(n11019), .ZN(n11021) );
  OAI21D1BWP30P140LVT U15691 ( .A1(n11023), .A2(n11022), .B(n11021), .ZN(
        n11024) );
  AOI21D1BWP30P140LVT U15692 ( .A1(n11025), .A2(n11024), .B(n11057), .ZN(N7098) );
  AOI211D1BWP30P140LVT U15693 ( .A1(i_cmd[148]), .A2(n11027), .B(i_cmd[132]), 
        .C(n11026), .ZN(n11028) );
  OAI21D1BWP30P140LVT U15694 ( .A1(n11030), .A2(n11029), .B(n11028), .ZN(
        n11031) );
  AOI21D1BWP30P140LVT U15695 ( .A1(n11032), .A2(n11031), .B(n11173), .ZN(N6882) );
  AOI211D1BWP30P140LVT U15696 ( .A1(i_cmd[84]), .A2(n11034), .B(i_cmd[68]), 
        .C(n11033), .ZN(n11035) );
  OAI21D1BWP30P140LVT U15697 ( .A1(n11037), .A2(n11036), .B(n11035), .ZN(
        n11038) );
  AOI21D1BWP30P140LVT U15698 ( .A1(n11039), .A2(n11038), .B(n11181), .ZN(N6450) );
  AOI211D1BWP30P140LVT U15699 ( .A1(i_cmd[60]), .A2(i_cmd[44]), .B(n11040), 
        .C(i_cmd[36]), .ZN(n11041) );
  INR2D1BWP30P140LVT U15700 ( .A1(n11042), .B1(n11041), .ZN(n11043) );
  AOI211D1BWP30P140LVT U15701 ( .A1(i_cmd[52]), .A2(n11044), .B(n11043), .C(
        n11181), .ZN(N6234) );
  AOI211D1BWP30P140LVT U15702 ( .A1(i_cmd[20]), .A2(n11046), .B(i_cmd[4]), .C(
        n11045), .ZN(n11047) );
  OAI21D1BWP30P140LVT U15703 ( .A1(n11049), .A2(n11048), .B(n11047), .ZN(
        n11050) );
  AOI21D1BWP30P140LVT U15704 ( .A1(n11051), .A2(n11050), .B(n11181), .ZN(N6018) );
  AOI211D1BWP30P140LVT U15705 ( .A1(i_cmd[243]), .A2(n11053), .B(i_cmd[227]), 
        .C(n11052), .ZN(n11054) );
  OAI21D1BWP30P140LVT U15706 ( .A1(n11056), .A2(n11055), .B(n11054), .ZN(
        n11058) );
  AOI21D1BWP30P140LVT U15707 ( .A1(n11059), .A2(n11058), .B(n11057), .ZN(N5656) );
  AOI211D1BWP30P140LVT U15708 ( .A1(i_cmd[219]), .A2(i_cmd[203]), .B(
        i_cmd[195]), .C(n11060), .ZN(n11061) );
  INR2D1BWP30P140LVT U15709 ( .A1(n11062), .B1(n11061), .ZN(n11063) );
  AOI211D1BWP30P140LVT U15710 ( .A1(i_cmd[211]), .A2(n11064), .B(n11063), .C(
        n11181), .ZN(N5568) );
  AOI211D1BWP30P140LVT U15711 ( .A1(i_cmd[171]), .A2(i_cmd[187]), .B(
        i_cmd[163]), .C(n11065), .ZN(n11066) );
  INR2D1BWP30P140LVT U15712 ( .A1(n11067), .B1(n11066), .ZN(n11068) );
  AOI211D1BWP30P140LVT U15713 ( .A1(i_cmd[179]), .A2(n11069), .B(n11068), .C(
        n11181), .ZN(N5480) );
  AOI211D1BWP30P140LVT U15714 ( .A1(i_cmd[155]), .A2(i_cmd[139]), .B(
        i_cmd[131]), .C(n11070), .ZN(n11071) );
  INR2D1BWP30P140LVT U15715 ( .A1(n11072), .B1(n11071), .ZN(n11073) );
  AOI211D1BWP30P140LVT U15716 ( .A1(i_cmd[147]), .A2(n11074), .B(n11073), .C(
        n11181), .ZN(N5392) );
  AOI211D1BWP30P140LVT U15717 ( .A1(i_cmd[115]), .A2(n11076), .B(i_cmd[99]), 
        .C(n11075), .ZN(n11077) );
  OAI21D1BWP30P140LVT U15718 ( .A1(n11079), .A2(n11078), .B(n11077), .ZN(
        n11080) );
  AOI21D1BWP30P140LVT U15719 ( .A1(n11081), .A2(n11080), .B(n11181), .ZN(N5304) );
  AOI211D1BWP30P140LVT U15720 ( .A1(i_cmd[83]), .A2(n11083), .B(i_cmd[67]), 
        .C(n11082), .ZN(n11084) );
  OAI21D1BWP30P140LVT U15721 ( .A1(n11086), .A2(n11085), .B(n11084), .ZN(
        n11087) );
  AOI21D1BWP30P140LVT U15722 ( .A1(n11088), .A2(n11087), .B(n11181), .ZN(N5216) );
  AOI211D1BWP30P140LVT U15723 ( .A1(i_cmd[51]), .A2(n11090), .B(i_cmd[35]), 
        .C(n11089), .ZN(n11091) );
  OAI21D1BWP30P140LVT U15724 ( .A1(n11093), .A2(n11092), .B(n11091), .ZN(
        n11094) );
  AOI21D1BWP30P140LVT U15725 ( .A1(n11095), .A2(n11094), .B(n11181), .ZN(N5128) );
  AOI211D1BWP30P140LVT U15726 ( .A1(i_cmd[218]), .A2(i_cmd[202]), .B(n11096), 
        .C(i_cmd[194]), .ZN(n11097) );
  INR2D1BWP30P140LVT U15727 ( .A1(n11098), .B1(n11097), .ZN(n11099) );
  AOI211D1BWP30P140LVT U15728 ( .A1(i_cmd[210]), .A2(n11100), .B(n11099), .C(
        n11181), .ZN(N4590) );
  AOI211D1BWP30P140LVT U15729 ( .A1(i_cmd[122]), .A2(i_cmd[106]), .B(i_cmd[98]), .C(n11101), .ZN(n11102) );
  INR2D1BWP30P140LVT U15730 ( .A1(n11103), .B1(n11102), .ZN(n11104) );
  AOI211D1BWP30P140LVT U15731 ( .A1(i_cmd[114]), .A2(n11105), .B(n11104), .C(
        n11181), .ZN(N3942) );
  AOI211D1BWP30P140LVT U15732 ( .A1(i_cmd[50]), .A2(n11107), .B(i_cmd[34]), 
        .C(n11106), .ZN(n11108) );
  OAI21D1BWP30P140LVT U15733 ( .A1(n11110), .A2(n11109), .B(n11108), .ZN(
        n11111) );
  AOI21D1BWP30P140LVT U15734 ( .A1(n11112), .A2(n11111), .B(n11173), .ZN(N3510) );
  AOI211D1BWP30P140LVT U15735 ( .A1(i_cmd[241]), .A2(n11114), .B(i_cmd[225]), 
        .C(n11113), .ZN(n11115) );
  OAI21D1BWP30P140LVT U15736 ( .A1(n11117), .A2(n11116), .B(n11115), .ZN(
        n11118) );
  AOI21D1BWP30P140LVT U15737 ( .A1(n11119), .A2(n11118), .B(n11173), .ZN(N2932) );
  AOI211D1BWP30P140LVT U15738 ( .A1(i_cmd[201]), .A2(i_cmd[217]), .B(
        i_cmd[193]), .C(n11120), .ZN(n11121) );
  INR2D1BWP30P140LVT U15739 ( .A1(n11122), .B1(n11121), .ZN(n11123) );
  AOI211D1BWP30P140LVT U15740 ( .A1(i_cmd[209]), .A2(n11124), .B(n11123), .C(
        n11181), .ZN(N2844) );
  AOI211D1BWP30P140LVT U15741 ( .A1(i_cmd[145]), .A2(n11126), .B(i_cmd[129]), 
        .C(n11125), .ZN(n11127) );
  OAI21D1BWP30P140LVT U15742 ( .A1(n11129), .A2(n11128), .B(n11127), .ZN(
        n11130) );
  AOI21D1BWP30P140LVT U15743 ( .A1(n11131), .A2(n11130), .B(n11173), .ZN(N2668) );
  AOI211D1BWP30P140LVT U15744 ( .A1(i_cmd[89]), .A2(i_cmd[73]), .B(n11132), 
        .C(i_cmd[65]), .ZN(n11133) );
  INR2D1BWP30P140LVT U15745 ( .A1(n11134), .B1(n11133), .ZN(n11135) );
  AOI211D1BWP30P140LVT U15746 ( .A1(i_cmd[81]), .A2(n11136), .B(n11135), .C(
        n11181), .ZN(N2492) );
  AOI211D1BWP30P140LVT U15747 ( .A1(i_cmd[49]), .A2(n11138), .B(i_cmd[33]), 
        .C(n11137), .ZN(n11139) );
  OAI21D1BWP30P140LVT U15748 ( .A1(n11141), .A2(n11140), .B(n11139), .ZN(
        n11142) );
  AOI21D1BWP30P140LVT U15749 ( .A1(n11143), .A2(n11142), .B(n11173), .ZN(N2404) );
  AOI211D1BWP30P140LVT U15750 ( .A1(i_cmd[17]), .A2(n11145), .B(i_cmd[1]), .C(
        n11144), .ZN(n11146) );
  OAI21D1BWP30P140LVT U15751 ( .A1(n11148), .A2(n11147), .B(n11146), .ZN(
        n11149) );
  AOI21D1BWP30P140LVT U15752 ( .A1(n11150), .A2(n11149), .B(n11173), .ZN(N2316) );
  AOI211D1BWP30P140LVT U15753 ( .A1(i_cmd[216]), .A2(i_cmd[200]), .B(
        i_cmd[192]), .C(n11151), .ZN(n11152) );
  INR2D1BWP30P140LVT U15754 ( .A1(n11153), .B1(n11152), .ZN(n11154) );
  AOI211D1BWP30P140LVT U15755 ( .A1(i_cmd[208]), .A2(n11155), .B(n11154), .C(
        n11181), .ZN(N1862) );
  AOI211D1BWP30P140LVT U15756 ( .A1(i_cmd[168]), .A2(i_cmd[184]), .B(
        i_cmd[160]), .C(n11156), .ZN(n11157) );
  INR2D1BWP30P140LVT U15757 ( .A1(n11158), .B1(n11157), .ZN(n11159) );
  AOI211D1BWP30P140LVT U15758 ( .A1(i_cmd[176]), .A2(n11160), .B(n11159), .C(
        n11181), .ZN(N1642) );
  AOI211D1BWP30P140LVT U15759 ( .A1(i_cmd[144]), .A2(n11162), .B(i_cmd[128]), 
        .C(n11161), .ZN(n11163) );
  OAI21D1BWP30P140LVT U15760 ( .A1(n11165), .A2(n11164), .B(n11163), .ZN(
        n11166) );
  AOI21D1BWP30P140LVT U15761 ( .A1(n11167), .A2(n11166), .B(n11173), .ZN(N1422) );
  AOI211D1BWP30P140LVT U15762 ( .A1(i_cmd[80]), .A2(n11169), .B(i_cmd[64]), 
        .C(n11168), .ZN(n11170) );
  OAI21D1BWP30P140LVT U15763 ( .A1(n11172), .A2(n11171), .B(n11170), .ZN(
        n11174) );
  AOI21D1BWP30P140LVT U15764 ( .A1(n11175), .A2(n11174), .B(n11173), .ZN(N982)
         );
  AOI211D1BWP30P140LVT U15765 ( .A1(i_cmd[48]), .A2(n11177), .B(i_cmd[32]), 
        .C(n11176), .ZN(n11178) );
  OAI21D1BWP30P140LVT U15766 ( .A1(n11180), .A2(n11179), .B(n11178), .ZN(
        n11182) );
  AOI21D1BWP30P140LVT U15767 ( .A1(n11183), .A2(n11182), .B(n11181), .ZN(N762)
         );
  AOI22D1BWP30P140LVT U15768 ( .A1(n11339), .A2(inner_first_stage_data_reg[64]), .B1(n11342), .B2(inner_first_stage_data_reg[96]), .ZN(n11187) );
  AOI22D1BWP30P140LVT U15769 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[128]), .B1(n11345), .B2(
        inner_first_stage_data_reg[0]), .ZN(n11186) );
  AOI22D1BWP30P140LVT U15770 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[192]), .B1(n11343), .B2(
        inner_first_stage_data_reg[224]), .ZN(n11185) );
  ND4D1BWP30P140LVT U15771 ( .A1(n11187), .A2(n11186), .A3(n11185), .A4(n11184), .ZN(n11188) );
  AO21D1BWP30P140LVT U15772 ( .A1(n11351), .A2(inner_first_stage_data_reg[160]), .B(n11188), .Z(N2229) );
  AOI22D1BWP30P140LVT U15773 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[129]), .B1(n11342), .B2(
        inner_first_stage_data_reg[97]), .ZN(n11192) );
  AOI22D1BWP30P140LVT U15774 ( .A1(n11339), .A2(inner_first_stage_data_reg[65]), .B1(n11341), .B2(inner_first_stage_data_reg[193]), .ZN(n11191) );
  AOI22D1BWP30P140LVT U15775 ( .A1(n11345), .A2(inner_first_stage_data_reg[1]), 
        .B1(n11343), .B2(inner_first_stage_data_reg[225]), .ZN(n11190) );
  ND4D1BWP30P140LVT U15776 ( .A1(n11192), .A2(n11191), .A3(n11190), .A4(n11189), .ZN(n11193) );
  AO21D1BWP30P140LVT U15777 ( .A1(n11344), .A2(inner_first_stage_data_reg[33]), 
        .B(n11193), .Z(N2230) );
  AOI22D1BWP30P140LVT U15778 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[130]), .B1(n11339), .B2(
        inner_first_stage_data_reg[66]), .ZN(n11197) );
  AOI22D1BWP30P140LVT U15779 ( .A1(n11345), .A2(inner_first_stage_data_reg[2]), 
        .B1(n11342), .B2(inner_first_stage_data_reg[98]), .ZN(n11196) );
  AOI22D1BWP30P140LVT U15780 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[194]), .B1(n11343), .B2(
        inner_first_stage_data_reg[226]), .ZN(n11195) );
  ND4D1BWP30P140LVT U15781 ( .A1(n11197), .A2(n11196), .A3(n11195), .A4(n11194), .ZN(n11198) );
  AO21D1BWP30P140LVT U15782 ( .A1(n11344), .A2(inner_first_stage_data_reg[34]), 
        .B(n11198), .Z(N2231) );
  AOI22D1BWP30P140LVT U15783 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[131]), .B1(n11339), .B2(
        inner_first_stage_data_reg[67]), .ZN(n11202) );
  AOI22D1BWP30P140LVT U15784 ( .A1(n11342), .A2(inner_first_stage_data_reg[99]), .B1(n11343), .B2(inner_first_stage_data_reg[227]), .ZN(n11201) );
  AOI22D1BWP30P140LVT U15785 ( .A1(n11345), .A2(inner_first_stage_data_reg[3]), 
        .B1(n11344), .B2(inner_first_stage_data_reg[35]), .ZN(n11200) );
  ND2D1BWP30P140LVT U15786 ( .A1(n11341), .A2(inner_first_stage_data_reg[195]), 
        .ZN(n11199) );
  ND4D1BWP30P140LVT U15787 ( .A1(n11202), .A2(n11201), .A3(n11200), .A4(n11199), .ZN(n11203) );
  AO21D1BWP30P140LVT U15788 ( .A1(n11351), .A2(inner_first_stage_data_reg[163]), .B(n11203), .Z(N2232) );
  AOI22D1BWP30P140LVT U15789 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[132]), .B1(n11342), .B2(
        inner_first_stage_data_reg[100]), .ZN(n11207) );
  AOI22D1BWP30P140LVT U15790 ( .A1(n11345), .A2(inner_first_stage_data_reg[4]), 
        .B1(n11339), .B2(inner_first_stage_data_reg[68]), .ZN(n11206) );
  AOI22D1BWP30P140LVT U15791 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[196]), .B1(n11343), .B2(
        inner_first_stage_data_reg[228]), .ZN(n11205) );
  ND4D1BWP30P140LVT U15792 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(n11208) );
  AO21D1BWP30P140LVT U15793 ( .A1(n11351), .A2(inner_first_stage_data_reg[164]), .B(n11208), .Z(N2233) );
  AOI22D1BWP30P140LVT U15794 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[133]), .B1(n11339), .B2(
        inner_first_stage_data_reg[69]), .ZN(n11212) );
  AOI22D1BWP30P140LVT U15795 ( .A1(n11342), .A2(
        inner_first_stage_data_reg[101]), .B1(n11341), .B2(
        inner_first_stage_data_reg[197]), .ZN(n11211) );
  AOI22D1BWP30P140LVT U15796 ( .A1(n11351), .A2(
        inner_first_stage_data_reg[165]), .B1(n11343), .B2(
        inner_first_stage_data_reg[229]), .ZN(n11210) );
  ND4D1BWP30P140LVT U15797 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(n11213) );
  AO21D1BWP30P140LVT U15798 ( .A1(n11344), .A2(inner_first_stage_data_reg[37]), 
        .B(n11213), .Z(N2234) );
  AOI22D1BWP30P140LVT U15799 ( .A1(n11339), .A2(inner_first_stage_data_reg[70]), .B1(n11342), .B2(inner_first_stage_data_reg[102]), .ZN(n11217) );
  AOI22D1BWP30P140LVT U15800 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[134]), .B1(n11345), .B2(
        inner_first_stage_data_reg[6]), .ZN(n11216) );
  AOI22D1BWP30P140LVT U15801 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[198]), .B1(n11343), .B2(
        inner_first_stage_data_reg[230]), .ZN(n11215) );
  ND4D1BWP30P140LVT U15802 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(n11218) );
  AO21D1BWP30P140LVT U15803 ( .A1(n11344), .A2(inner_first_stage_data_reg[38]), 
        .B(n11218), .Z(N2235) );
  AOI22D1BWP30P140LVT U15804 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[135]), .B1(n11342), .B2(
        inner_first_stage_data_reg[103]), .ZN(n11222) );
  AOI22D1BWP30P140LVT U15805 ( .A1(n11339), .A2(inner_first_stage_data_reg[71]), .B1(n11341), .B2(inner_first_stage_data_reg[199]), .ZN(n11221) );
  AOI22D1BWP30P140LVT U15806 ( .A1(n11351), .A2(
        inner_first_stage_data_reg[167]), .B1(n11345), .B2(
        inner_first_stage_data_reg[7]), .ZN(n11220) );
  ND2D1BWP30P140LVT U15807 ( .A1(n11343), .A2(inner_first_stage_data_reg[231]), 
        .ZN(n11219) );
  ND4D1BWP30P140LVT U15808 ( .A1(n11222), .A2(n11221), .A3(n11220), .A4(n11219), .ZN(n11223) );
  AO21D1BWP30P140LVT U15809 ( .A1(n11344), .A2(inner_first_stage_data_reg[39]), 
        .B(n11223), .Z(N2236) );
  AOI22D1BWP30P140LVT U15810 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[136]), .B1(n11339), .B2(
        inner_first_stage_data_reg[72]), .ZN(n11227) );
  AOI22D1BWP30P140LVT U15811 ( .A1(n11345), .A2(inner_first_stage_data_reg[8]), 
        .B1(n11342), .B2(inner_first_stage_data_reg[104]), .ZN(n11226) );
  AOI22D1BWP30P140LVT U15812 ( .A1(n11351), .A2(
        inner_first_stage_data_reg[168]), .B1(n11341), .B2(
        inner_first_stage_data_reg[200]), .ZN(n11225) );
  ND2D1BWP30P140LVT U15813 ( .A1(n11343), .A2(inner_first_stage_data_reg[232]), 
        .ZN(n11224) );
  ND4D1BWP30P140LVT U15814 ( .A1(n11227), .A2(n11226), .A3(n11225), .A4(n11224), .ZN(n11228) );
  AO21D1BWP30P140LVT U15815 ( .A1(n11344), .A2(inner_first_stage_data_reg[40]), 
        .B(n11228), .Z(N2237) );
  AOI22D1BWP30P140LVT U15816 ( .A1(n11339), .A2(inner_first_stage_data_reg[73]), .B1(n11342), .B2(inner_first_stage_data_reg[105]), .ZN(n11232) );
  AOI22D1BWP30P140LVT U15817 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[137]), .B1(n11341), .B2(
        inner_first_stage_data_reg[201]), .ZN(n11231) );
  AOI22D1BWP30P140LVT U15818 ( .A1(n11345), .A2(inner_first_stage_data_reg[9]), 
        .B1(n11343), .B2(inner_first_stage_data_reg[233]), .ZN(n11230) );
  ND4D1BWP30P140LVT U15819 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(n11233) );
  AO21D1BWP30P140LVT U15820 ( .A1(n11344), .A2(inner_first_stage_data_reg[41]), 
        .B(n11233), .Z(N2238) );
  AOI22D1BWP30P140LVT U15821 ( .A1(n11339), .A2(inner_first_stage_data_reg[74]), .B1(n11342), .B2(inner_first_stage_data_reg[106]), .ZN(n11237) );
  AOI22D1BWP30P140LVT U15822 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[138]), .B1(n11345), .B2(
        inner_first_stage_data_reg[10]), .ZN(n11236) );
  AOI22D1BWP30P140LVT U15823 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[202]), .B1(n11343), .B2(
        inner_first_stage_data_reg[234]), .ZN(n11235) );
  ND4D1BWP30P140LVT U15824 ( .A1(n11237), .A2(n11236), .A3(n11235), .A4(n11234), .ZN(n11238) );
  AO21D1BWP30P140LVT U15825 ( .A1(n11344), .A2(inner_first_stage_data_reg[42]), 
        .B(n11238), .Z(N2239) );
  AOI22D1BWP30P140LVT U15826 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[139]), .B1(n11342), .B2(
        inner_first_stage_data_reg[107]), .ZN(n11242) );
  AOI22D1BWP30P140LVT U15827 ( .A1(n11345), .A2(inner_first_stage_data_reg[11]), .B1(n11339), .B2(inner_first_stage_data_reg[75]), .ZN(n11241) );
  AOI22D1BWP30P140LVT U15828 ( .A1(n11344), .A2(inner_first_stage_data_reg[43]), .B1(n11341), .B2(inner_first_stage_data_reg[203]), .ZN(n11240) );
  ND2D1BWP30P140LVT U15829 ( .A1(n11343), .A2(inner_first_stage_data_reg[235]), 
        .ZN(n11239) );
  ND4D1BWP30P140LVT U15830 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(n11243) );
  AO21D1BWP30P140LVT U15831 ( .A1(n11351), .A2(inner_first_stage_data_reg[171]), .B(n11243), .Z(N2240) );
  AOI22D1BWP30P140LVT U15832 ( .A1(n11339), .A2(inner_first_stage_data_reg[76]), .B1(n11342), .B2(inner_first_stage_data_reg[108]), .ZN(n11247) );
  AOI22D1BWP30P140LVT U15833 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[140]), .B1(n11343), .B2(
        inner_first_stage_data_reg[236]), .ZN(n11246) );
  AOI22D1BWP30P140LVT U15834 ( .A1(n11344), .A2(inner_first_stage_data_reg[44]), .B1(n11341), .B2(inner_first_stage_data_reg[204]), .ZN(n11245) );
  ND4D1BWP30P140LVT U15835 ( .A1(n11247), .A2(n11246), .A3(n11245), .A4(n11244), .ZN(n11248) );
  AO21D1BWP30P140LVT U15836 ( .A1(n11351), .A2(inner_first_stage_data_reg[172]), .B(n11248), .Z(N2241) );
  AOI22D1BWP30P140LVT U15837 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[141]), .B1(n11339), .B2(
        inner_first_stage_data_reg[77]), .ZN(n11252) );
  AOI22D1BWP30P140LVT U15838 ( .A1(n11345), .A2(inner_first_stage_data_reg[13]), .B1(n11342), .B2(inner_first_stage_data_reg[109]), .ZN(n11251) );
  AOI22D1BWP30P140LVT U15839 ( .A1(n11344), .A2(inner_first_stage_data_reg[45]), .B1(n11343), .B2(inner_first_stage_data_reg[237]), .ZN(n11250) );
  ND2D1BWP30P140LVT U15840 ( .A1(n11341), .A2(inner_first_stage_data_reg[205]), 
        .ZN(n11249) );
  ND4D1BWP30P140LVT U15841 ( .A1(n11252), .A2(n11251), .A3(n11250), .A4(n11249), .ZN(n11253) );
  AO21D1BWP30P140LVT U15842 ( .A1(n11351), .A2(inner_first_stage_data_reg[173]), .B(n11253), .Z(N2242) );
  AOI22D1BWP30P140LVT U15843 ( .A1(n11339), .A2(inner_first_stage_data_reg[78]), .B1(n11342), .B2(inner_first_stage_data_reg[110]), .ZN(n11257) );
  AOI22D1BWP30P140LVT U15844 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[142]), .B1(n11345), .B2(
        inner_first_stage_data_reg[14]), .ZN(n11256) );
  AOI22D1BWP30P140LVT U15845 ( .A1(n11351), .A2(
        inner_first_stage_data_reg[174]), .B1(n11343), .B2(
        inner_first_stage_data_reg[238]), .ZN(n11255) );
  ND2D1BWP30P140LVT U15846 ( .A1(n11341), .A2(inner_first_stage_data_reg[206]), 
        .ZN(n11254) );
  ND4D1BWP30P140LVT U15847 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(n11258) );
  AO21D1BWP30P140LVT U15848 ( .A1(n11344), .A2(inner_first_stage_data_reg[46]), 
        .B(n11258), .Z(N2243) );
  AOI22D1BWP30P140LVT U15849 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[143]), .B1(n11339), .B2(
        inner_first_stage_data_reg[79]), .ZN(n11262) );
  AOI22D1BWP30P140LVT U15850 ( .A1(n11345), .A2(inner_first_stage_data_reg[15]), .B1(n11342), .B2(inner_first_stage_data_reg[111]), .ZN(n11261) );
  AOI22D1BWP30P140LVT U15851 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[207]), .B1(n11343), .B2(
        inner_first_stage_data_reg[239]), .ZN(n11260) );
  ND4D1BWP30P140LVT U15852 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n11259), .ZN(n11263) );
  AO21D1BWP30P140LVT U15853 ( .A1(n11344), .A2(inner_first_stage_data_reg[47]), 
        .B(n11263), .Z(N2244) );
  AOI22D1BWP30P140LVT U15854 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[144]), .B1(n11339), .B2(
        inner_first_stage_data_reg[80]), .ZN(n11267) );
  AOI22D1BWP30P140LVT U15855 ( .A1(n11345), .A2(inner_first_stage_data_reg[16]), .B1(n11342), .B2(inner_first_stage_data_reg[112]), .ZN(n11266) );
  AOI22D1BWP30P140LVT U15856 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[208]), .B1(n11343), .B2(
        inner_first_stage_data_reg[240]), .ZN(n11265) );
  ND4D1BWP30P140LVT U15857 ( .A1(n11267), .A2(n11266), .A3(n11265), .A4(n11264), .ZN(n11268) );
  AO21D1BWP30P140LVT U15858 ( .A1(n11344), .A2(inner_first_stage_data_reg[48]), 
        .B(n11268), .Z(N2245) );
  AOI22D1BWP30P140LVT U15859 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[145]), .B1(n11342), .B2(
        inner_first_stage_data_reg[113]), .ZN(n11272) );
  AOI22D1BWP30P140LVT U15860 ( .A1(n11339), .A2(inner_first_stage_data_reg[81]), .B1(n11341), .B2(inner_first_stage_data_reg[209]), .ZN(n11271) );
  AOI22D1BWP30P140LVT U15861 ( .A1(n11345), .A2(inner_first_stage_data_reg[17]), .B1(n11343), .B2(inner_first_stage_data_reg[241]), .ZN(n11270) );
  ND4D1BWP30P140LVT U15862 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(n11273) );
  AO21D1BWP30P140LVT U15863 ( .A1(n11344), .A2(inner_first_stage_data_reg[49]), 
        .B(n11273), .Z(N2246) );
  AOI22D1BWP30P140LVT U15864 ( .A1(n11339), .A2(inner_first_stage_data_reg[82]), .B1(n11342), .B2(inner_first_stage_data_reg[114]), .ZN(n11277) );
  AOI22D1BWP30P140LVT U15865 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[146]), .B1(n11345), .B2(
        inner_first_stage_data_reg[18]), .ZN(n11276) );
  AOI22D1BWP30P140LVT U15866 ( .A1(n11351), .A2(
        inner_first_stage_data_reg[178]), .B1(n11341), .B2(
        inner_first_stage_data_reg[210]), .ZN(n11275) );
  ND2D1BWP30P140LVT U15867 ( .A1(n11343), .A2(inner_first_stage_data_reg[242]), 
        .ZN(n11274) );
  ND4D1BWP30P140LVT U15868 ( .A1(n11277), .A2(n11276), .A3(n11275), .A4(n11274), .ZN(n11278) );
  AO21D1BWP30P140LVT U15869 ( .A1(n11344), .A2(inner_first_stage_data_reg[50]), 
        .B(n11278), .Z(N2247) );
  AOI22D1BWP30P140LVT U15870 ( .A1(n11339), .A2(inner_first_stage_data_reg[83]), .B1(n11342), .B2(inner_first_stage_data_reg[115]), .ZN(n11282) );
  AOI22D1BWP30P140LVT U15871 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[147]), .B1(n11343), .B2(
        inner_first_stage_data_reg[243]), .ZN(n11281) );
  AOI22D1BWP30P140LVT U15872 ( .A1(n11351), .A2(
        inner_first_stage_data_reg[179]), .B1(n11345), .B2(
        inner_first_stage_data_reg[19]), .ZN(n11280) );
  ND2D1BWP30P140LVT U15873 ( .A1(n11341), .A2(inner_first_stage_data_reg[211]), 
        .ZN(n11279) );
  ND4D1BWP30P140LVT U15874 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(n11283) );
  AO21D1BWP30P140LVT U15875 ( .A1(n11344), .A2(inner_first_stage_data_reg[51]), 
        .B(n11283), .Z(N2248) );
  AOI22D1BWP30P140LVT U15876 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[148]), .B1(n11342), .B2(
        inner_first_stage_data_reg[116]), .ZN(n11287) );
  AOI22D1BWP30P140LVT U15877 ( .A1(n11339), .A2(inner_first_stage_data_reg[84]), .B1(n11341), .B2(inner_first_stage_data_reg[212]), .ZN(n11286) );
  AOI22D1BWP30P140LVT U15878 ( .A1(n11345), .A2(inner_first_stage_data_reg[20]), .B1(n11343), .B2(inner_first_stage_data_reg[244]), .ZN(n11285) );
  ND4D1BWP30P140LVT U15879 ( .A1(n11287), .A2(n11286), .A3(n11285), .A4(n11284), .ZN(n11288) );
  AO21D1BWP30P140LVT U15880 ( .A1(n11344), .A2(inner_first_stage_data_reg[52]), 
        .B(n11288), .Z(N2249) );
  AOI22D1BWP30P140LVT U15881 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[149]), .B1(n11342), .B2(
        inner_first_stage_data_reg[117]), .ZN(n11292) );
  AOI22D1BWP30P140LVT U15882 ( .A1(n11339), .A2(inner_first_stage_data_reg[85]), .B1(n11341), .B2(inner_first_stage_data_reg[213]), .ZN(n11291) );
  AOI22D1BWP30P140LVT U15883 ( .A1(n11345), .A2(inner_first_stage_data_reg[21]), .B1(n11343), .B2(inner_first_stage_data_reg[245]), .ZN(n11290) );
  ND4D1BWP30P140LVT U15884 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(n11293) );
  AO21D1BWP30P140LVT U15885 ( .A1(n11351), .A2(inner_first_stage_data_reg[181]), .B(n11293), .Z(N2250) );
  AOI22D1BWP30P140LVT U15886 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[150]), .B1(n11342), .B2(
        inner_first_stage_data_reg[118]), .ZN(n11297) );
  AOI22D1BWP30P140LVT U15887 ( .A1(n11339), .A2(inner_first_stage_data_reg[86]), .B1(n11343), .B2(inner_first_stage_data_reg[246]), .ZN(n11296) );
  AOI22D1BWP30P140LVT U15888 ( .A1(n11345), .A2(inner_first_stage_data_reg[22]), .B1(n11341), .B2(inner_first_stage_data_reg[214]), .ZN(n11295) );
  ND4D1BWP30P140LVT U15889 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(n11298) );
  AO21D1BWP30P140LVT U15890 ( .A1(n11351), .A2(inner_first_stage_data_reg[182]), .B(n11298), .Z(N2251) );
  AOI22D1BWP30P140LVT U15891 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[151]), .B1(n11339), .B2(
        inner_first_stage_data_reg[87]), .ZN(n11302) );
  AOI22D1BWP30P140LVT U15892 ( .A1(n11342), .A2(
        inner_first_stage_data_reg[119]), .B1(n11341), .B2(
        inner_first_stage_data_reg[215]), .ZN(n11301) );
  AOI22D1BWP30P140LVT U15893 ( .A1(n11345), .A2(inner_first_stage_data_reg[23]), .B1(n11343), .B2(inner_first_stage_data_reg[247]), .ZN(n11300) );
  ND4D1BWP30P140LVT U15894 ( .A1(n11302), .A2(n11301), .A3(n11300), .A4(n11299), .ZN(n11303) );
  AO21D1BWP30P140LVT U15895 ( .A1(n11351), .A2(inner_first_stage_data_reg[183]), .B(n11303), .Z(N2252) );
  AOI22D1BWP30P140LVT U15896 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[152]), .B1(n11339), .B2(
        inner_first_stage_data_reg[88]), .ZN(n11307) );
  AOI22D1BWP30P140LVT U15897 ( .A1(n11345), .A2(inner_first_stage_data_reg[24]), .B1(n11342), .B2(inner_first_stage_data_reg[120]), .ZN(n11306) );
  AOI22D1BWP30P140LVT U15898 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[216]), .B1(n11343), .B2(
        inner_first_stage_data_reg[248]), .ZN(n11305) );
  ND4D1BWP30P140LVT U15899 ( .A1(n11307), .A2(n11306), .A3(n11305), .A4(n11304), .ZN(n11308) );
  AO21D1BWP30P140LVT U15900 ( .A1(n11344), .A2(inner_first_stage_data_reg[56]), 
        .B(n11308), .Z(N2253) );
  AOI22D1BWP30P140LVT U15901 ( .A1(n11339), .A2(inner_first_stage_data_reg[89]), .B1(n11342), .B2(inner_first_stage_data_reg[121]), .ZN(n11312) );
  AOI22D1BWP30P140LVT U15902 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[153]), .B1(n11343), .B2(
        inner_first_stage_data_reg[249]), .ZN(n11311) );
  AOI22D1BWP30P140LVT U15903 ( .A1(n11345), .A2(inner_first_stage_data_reg[25]), .B1(n11341), .B2(inner_first_stage_data_reg[217]), .ZN(n11310) );
  ND4D1BWP30P140LVT U15904 ( .A1(n11312), .A2(n11311), .A3(n11310), .A4(n11309), .ZN(n11313) );
  AO21D1BWP30P140LVT U15905 ( .A1(n11351), .A2(inner_first_stage_data_reg[185]), .B(n11313), .Z(N2254) );
  AOI22D1BWP30P140LVT U15906 ( .A1(n11339), .A2(inner_first_stage_data_reg[90]), .B1(n11342), .B2(inner_first_stage_data_reg[122]), .ZN(n11317) );
  AOI22D1BWP30P140LVT U15907 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[154]), .B1(n11341), .B2(
        inner_first_stage_data_reg[218]), .ZN(n11316) );
  AOI22D1BWP30P140LVT U15908 ( .A1(n11345), .A2(inner_first_stage_data_reg[26]), .B1(n11343), .B2(inner_first_stage_data_reg[250]), .ZN(n11315) );
  ND4D1BWP30P140LVT U15909 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(n11318) );
  AO21D1BWP30P140LVT U15910 ( .A1(n11344), .A2(inner_first_stage_data_reg[58]), 
        .B(n11318), .Z(N2255) );
  AOI22D1BWP30P140LVT U15911 ( .A1(n11339), .A2(inner_first_stage_data_reg[91]), .B1(n11342), .B2(inner_first_stage_data_reg[123]), .ZN(n11322) );
  AOI22D1BWP30P140LVT U15912 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[155]), .B1(n11345), .B2(
        inner_first_stage_data_reg[27]), .ZN(n11321) );
  AOI22D1BWP30P140LVT U15913 ( .A1(n11351), .A2(
        inner_first_stage_data_reg[187]), .B1(n11341), .B2(
        inner_first_stage_data_reg[219]), .ZN(n11320) );
  ND2D1BWP30P140LVT U15914 ( .A1(n11343), .A2(inner_first_stage_data_reg[251]), 
        .ZN(n11319) );
  ND4D1BWP30P140LVT U15915 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(n11323) );
  AO21D1BWP30P140LVT U15916 ( .A1(n11344), .A2(inner_first_stage_data_reg[59]), 
        .B(n11323), .Z(N2256) );
  AOI22D1BWP30P140LVT U15917 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[156]), .B1(n11339), .B2(
        inner_first_stage_data_reg[92]), .ZN(n11327) );
  AOI22D1BWP30P140LVT U15918 ( .A1(n11342), .A2(
        inner_first_stage_data_reg[124]), .B1(n11341), .B2(
        inner_first_stage_data_reg[220]), .ZN(n11326) );
  AOI22D1BWP30P140LVT U15919 ( .A1(n11345), .A2(inner_first_stage_data_reg[28]), .B1(n11343), .B2(inner_first_stage_data_reg[252]), .ZN(n11325) );
  ND4D1BWP30P140LVT U15920 ( .A1(n11327), .A2(n11326), .A3(n11325), .A4(n11324), .ZN(n11328) );
  AO21D1BWP30P140LVT U15921 ( .A1(n11351), .A2(inner_first_stage_data_reg[188]), .B(n11328), .Z(N2257) );
  AOI22D1BWP30P140LVT U15922 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[157]), .B1(n11342), .B2(
        inner_first_stage_data_reg[125]), .ZN(n11332) );
  AOI22D1BWP30P140LVT U15923 ( .A1(n11345), .A2(inner_first_stage_data_reg[29]), .B1(n11339), .B2(inner_first_stage_data_reg[93]), .ZN(n11331) );
  AOI22D1BWP30P140LVT U15924 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[221]), .B1(n11343), .B2(
        inner_first_stage_data_reg[253]), .ZN(n11330) );
  ND4D1BWP30P140LVT U15925 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(n11333) );
  AO21D1BWP30P140LVT U15926 ( .A1(n11344), .A2(inner_first_stage_data_reg[61]), 
        .B(n11333), .Z(N2258) );
  AOI22D1BWP30P140LVT U15927 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[158]), .B1(n11339), .B2(
        inner_first_stage_data_reg[94]), .ZN(n11337) );
  AOI22D1BWP30P140LVT U15928 ( .A1(n11345), .A2(inner_first_stage_data_reg[30]), .B1(n11342), .B2(inner_first_stage_data_reg[126]), .ZN(n11336) );
  AOI22D1BWP30P140LVT U15929 ( .A1(n11341), .A2(
        inner_first_stage_data_reg[222]), .B1(n11343), .B2(
        inner_first_stage_data_reg[254]), .ZN(n11335) );
  ND4D1BWP30P140LVT U15930 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(n11338) );
  AO21D1BWP30P140LVT U15931 ( .A1(n11344), .A2(inner_first_stage_data_reg[62]), 
        .B(n11338), .Z(N2259) );
  AOI22D1BWP30P140LVT U15932 ( .A1(n11340), .A2(
        inner_first_stage_data_reg[159]), .B1(n11339), .B2(
        inner_first_stage_data_reg[95]), .ZN(n11349) );
  AOI22D1BWP30P140LVT U15933 ( .A1(n11342), .A2(
        inner_first_stage_data_reg[127]), .B1(n11341), .B2(
        inner_first_stage_data_reg[223]), .ZN(n11348) );
  AOI22D1BWP30P140LVT U15934 ( .A1(n11344), .A2(inner_first_stage_data_reg[63]), .B1(n11343), .B2(inner_first_stage_data_reg[255]), .ZN(n11347) );
  ND4D1BWP30P140LVT U15935 ( .A1(n11349), .A2(n11348), .A3(n11347), .A4(n11346), .ZN(n11350) );
  AO21D1BWP30P140LVT U15936 ( .A1(n11351), .A2(inner_first_stage_data_reg[191]), .B(n11350), .Z(N2260) );
  AOI22D1BWP30P140LVT U15937 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[256]), .B1(n11476), .B2(
        inner_first_stage_data_reg[384]), .ZN(n11355) );
  AOI22D1BWP30P140LVT U15938 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[288]), .B1(n11481), .B2(
        inner_first_stage_data_reg[480]), .ZN(n11354) );
  AOI22D1BWP30P140LVT U15939 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[448]), .B1(n11478), .B2(
        inner_first_stage_data_reg[320]), .ZN(n11353) );
  AOI22D1BWP30P140LVT U15940 ( .A1(n11483), .A2(
        inner_first_stage_data_reg[352]), .B1(n11482), .B2(
        inner_first_stage_data_reg[416]), .ZN(n11352) );
  ND4D1BWP30P140LVT U15941 ( .A1(n11355), .A2(n11354), .A3(n11353), .A4(n11352), .ZN(N3079) );
  AOI22D1BWP30P140LVT U15942 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[257]), .B1(n11476), .B2(
        inner_first_stage_data_reg[385]), .ZN(n11359) );
  AOI22D1BWP30P140LVT U15943 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[449]), .B1(n11482), .B2(
        inner_first_stage_data_reg[417]), .ZN(n11358) );
  AOI22D1BWP30P140LVT U15944 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[289]), .B1(n11478), .B2(
        inner_first_stage_data_reg[321]), .ZN(n11357) );
  AOI22D1BWP30P140LVT U15945 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[481]), .B1(n11483), .B2(
        inner_first_stage_data_reg[353]), .ZN(n11356) );
  ND4D1BWP30P140LVT U15946 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(N3080) );
  AOI22D1BWP30P140LVT U15947 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[258]), .B1(n11476), .B2(
        inner_first_stage_data_reg[386]), .ZN(n11363) );
  AOI22D1BWP30P140LVT U15948 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[290]), .B1(n11480), .B2(
        inner_first_stage_data_reg[450]), .ZN(n11362) );
  AOI22D1BWP30P140LVT U15949 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[322]), .B1(n11482), .B2(
        inner_first_stage_data_reg[418]), .ZN(n11361) );
  AOI22D1BWP30P140LVT U15950 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[482]), .B1(n11483), .B2(
        inner_first_stage_data_reg[354]), .ZN(n11360) );
  ND4D1BWP30P140LVT U15951 ( .A1(n11363), .A2(n11362), .A3(n11361), .A4(n11360), .ZN(N3081) );
  AOI22D1BWP30P140LVT U15952 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[259]), .B1(n11476), .B2(
        inner_first_stage_data_reg[387]), .ZN(n11367) );
  AOI22D1BWP30P140LVT U15953 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[291]), .B1(n11482), .B2(
        inner_first_stage_data_reg[419]), .ZN(n11366) );
  AOI22D1BWP30P140LVT U15954 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[451]), .B1(n11478), .B2(
        inner_first_stage_data_reg[323]), .ZN(n11365) );
  AOI22D1BWP30P140LVT U15955 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[483]), .B1(n11483), .B2(
        inner_first_stage_data_reg[355]), .ZN(n11364) );
  ND4D1BWP30P140LVT U15956 ( .A1(n11367), .A2(n11366), .A3(n11365), .A4(n11364), .ZN(N3082) );
  AOI22D1BWP30P140LVT U15957 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[260]), .B1(n11476), .B2(
        inner_first_stage_data_reg[388]), .ZN(n11371) );
  AOI22D1BWP30P140LVT U15958 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[292]), .B1(n11482), .B2(
        inner_first_stage_data_reg[420]), .ZN(n11370) );
  AOI22D1BWP30P140LVT U15959 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[484]), .B1(n11483), .B2(
        inner_first_stage_data_reg[356]), .ZN(n11369) );
  AOI22D1BWP30P140LVT U15960 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[452]), .B1(n11478), .B2(
        inner_first_stage_data_reg[324]), .ZN(n11368) );
  ND4D1BWP30P140LVT U15961 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(N3083) );
  AOI22D1BWP30P140LVT U15962 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[261]), .B1(n11476), .B2(
        inner_first_stage_data_reg[389]), .ZN(n11375) );
  AOI22D1BWP30P140LVT U15963 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[453]), .B1(n11482), .B2(
        inner_first_stage_data_reg[421]), .ZN(n11374) );
  AOI22D1BWP30P140LVT U15964 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[293]), .B1(n11483), .B2(
        inner_first_stage_data_reg[357]), .ZN(n11373) );
  AOI22D1BWP30P140LVT U15965 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[485]), .B1(n11478), .B2(
        inner_first_stage_data_reg[325]), .ZN(n11372) );
  ND4D1BWP30P140LVT U15966 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(N3084) );
  AOI22D1BWP30P140LVT U15967 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[262]), .B1(n11476), .B2(
        inner_first_stage_data_reg[390]), .ZN(n11379) );
  AOI22D1BWP30P140LVT U15968 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[326]), .B1(n11483), .B2(
        inner_first_stage_data_reg[358]), .ZN(n11378) );
  AOI22D1BWP30P140LVT U15969 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[294]), .B1(n11481), .B2(
        inner_first_stage_data_reg[486]), .ZN(n11377) );
  AOI22D1BWP30P140LVT U15970 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[454]), .B1(n11482), .B2(
        inner_first_stage_data_reg[422]), .ZN(n11376) );
  ND4D1BWP30P140LVT U15971 ( .A1(n11379), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(N3085) );
  AOI22D1BWP30P140LVT U15972 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[263]), .B1(n11476), .B2(
        inner_first_stage_data_reg[391]), .ZN(n11383) );
  AOI22D1BWP30P140LVT U15973 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[487]), .B1(n11478), .B2(
        inner_first_stage_data_reg[327]), .ZN(n11382) );
  AOI22D1BWP30P140LVT U15974 ( .A1(n11483), .A2(
        inner_first_stage_data_reg[359]), .B1(n11482), .B2(
        inner_first_stage_data_reg[423]), .ZN(n11381) );
  AOI22D1BWP30P140LVT U15975 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[295]), .B1(n11480), .B2(
        inner_first_stage_data_reg[455]), .ZN(n11380) );
  ND4D1BWP30P140LVT U15976 ( .A1(n11383), .A2(n11382), .A3(n11381), .A4(n11380), .ZN(N3086) );
  AOI22D1BWP30P140LVT U15977 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[264]), .B1(n11476), .B2(
        inner_first_stage_data_reg[392]), .ZN(n11387) );
  AOI22D1BWP30P140LVT U15978 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[488]), .B1(n11483), .B2(
        inner_first_stage_data_reg[360]), .ZN(n11386) );
  AOI22D1BWP30P140LVT U15979 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[296]), .B1(n11482), .B2(
        inner_first_stage_data_reg[424]), .ZN(n11385) );
  AOI22D1BWP30P140LVT U15980 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[456]), .B1(n11478), .B2(
        inner_first_stage_data_reg[328]), .ZN(n11384) );
  ND4D1BWP30P140LVT U15981 ( .A1(n11387), .A2(n11386), .A3(n11385), .A4(n11384), .ZN(N3087) );
  AOI22D1BWP30P140LVT U15982 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[265]), .B1(n11476), .B2(
        inner_first_stage_data_reg[393]), .ZN(n11391) );
  AOI22D1BWP30P140LVT U15983 ( .A1(n11483), .A2(
        inner_first_stage_data_reg[361]), .B1(n11482), .B2(
        inner_first_stage_data_reg[425]), .ZN(n11390) );
  AOI22D1BWP30P140LVT U15984 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[297]), .B1(n11480), .B2(
        inner_first_stage_data_reg[457]), .ZN(n11389) );
  AOI22D1BWP30P140LVT U15985 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[489]), .B1(n11478), .B2(
        inner_first_stage_data_reg[329]), .ZN(n11388) );
  ND4D1BWP30P140LVT U15986 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(N3088) );
  AOI22D1BWP30P140LVT U15987 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[266]), .B1(n11476), .B2(
        inner_first_stage_data_reg[394]), .ZN(n11395) );
  AOI22D1BWP30P140LVT U15988 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[298]), .B1(n11481), .B2(
        inner_first_stage_data_reg[490]), .ZN(n11394) );
  AOI22D1BWP30P140LVT U15989 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[330]), .B1(n11482), .B2(
        inner_first_stage_data_reg[426]), .ZN(n11393) );
  AOI22D1BWP30P140LVT U15990 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[458]), .B1(n11483), .B2(
        inner_first_stage_data_reg[362]), .ZN(n11392) );
  ND4D1BWP30P140LVT U15991 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(N3089) );
  AOI22D1BWP30P140LVT U15992 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[267]), .B1(n11476), .B2(
        inner_first_stage_data_reg[395]), .ZN(n11399) );
  AOI22D1BWP30P140LVT U15993 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[491]), .B1(n11480), .B2(
        inner_first_stage_data_reg[459]), .ZN(n11398) );
  AOI22D1BWP30P140LVT U15994 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[331]), .B1(n11482), .B2(
        inner_first_stage_data_reg[427]), .ZN(n11397) );
  AOI22D1BWP30P140LVT U15995 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[299]), .B1(n11483), .B2(
        inner_first_stage_data_reg[363]), .ZN(n11396) );
  ND4D1BWP30P140LVT U15996 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(N3090) );
  AOI22D1BWP30P140LVT U15997 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[268]), .B1(n11476), .B2(
        inner_first_stage_data_reg[396]), .ZN(n11403) );
  AOI22D1BWP30P140LVT U15998 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[300]), .B1(n11482), .B2(
        inner_first_stage_data_reg[428]), .ZN(n11402) );
  AOI22D1BWP30P140LVT U15999 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[492]), .B1(n11478), .B2(
        inner_first_stage_data_reg[332]), .ZN(n11401) );
  AOI22D1BWP30P140LVT U16000 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[460]), .B1(n11483), .B2(
        inner_first_stage_data_reg[364]), .ZN(n11400) );
  ND4D1BWP30P140LVT U16001 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(N3091) );
  AOI22D1BWP30P140LVT U16002 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[269]), .B1(n11476), .B2(
        inner_first_stage_data_reg[397]), .ZN(n11407) );
  AOI22D1BWP30P140LVT U16003 ( .A1(n11483), .A2(
        inner_first_stage_data_reg[365]), .B1(n11482), .B2(
        inner_first_stage_data_reg[429]), .ZN(n11406) );
  AOI22D1BWP30P140LVT U16004 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[301]), .B1(n11481), .B2(
        inner_first_stage_data_reg[493]), .ZN(n11405) );
  AOI22D1BWP30P140LVT U16005 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[461]), .B1(n11478), .B2(
        inner_first_stage_data_reg[333]), .ZN(n11404) );
  ND4D1BWP30P140LVT U16006 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(N3092) );
  AOI22D1BWP30P140LVT U16007 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[270]), .B1(n11476), .B2(
        inner_first_stage_data_reg[398]), .ZN(n11411) );
  AOI22D1BWP30P140LVT U16008 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[494]), .B1(n11478), .B2(
        inner_first_stage_data_reg[334]), .ZN(n11410) );
  AOI22D1BWP30P140LVT U16009 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[462]), .B1(n11482), .B2(
        inner_first_stage_data_reg[430]), .ZN(n11409) );
  AOI22D1BWP30P140LVT U16010 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[302]), .B1(n11483), .B2(
        inner_first_stage_data_reg[366]), .ZN(n11408) );
  ND4D1BWP30P140LVT U16011 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(N3093) );
  AOI22D1BWP30P140LVT U16012 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[271]), .B1(n11476), .B2(
        inner_first_stage_data_reg[399]), .ZN(n11415) );
  AOI22D1BWP30P140LVT U16013 ( .A1(n11483), .A2(
        inner_first_stage_data_reg[367]), .B1(n11482), .B2(
        inner_first_stage_data_reg[431]), .ZN(n11414) );
  AOI22D1BWP30P140LVT U16014 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[463]), .B1(n11478), .B2(
        inner_first_stage_data_reg[335]), .ZN(n11413) );
  AOI22D1BWP30P140LVT U16015 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[303]), .B1(n11481), .B2(
        inner_first_stage_data_reg[495]), .ZN(n11412) );
  ND4D1BWP30P140LVT U16016 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(N3094) );
  AOI22D1BWP30P140LVT U16017 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[272]), .B1(n11476), .B2(
        inner_first_stage_data_reg[400]), .ZN(n11419) );
  AOI22D1BWP30P140LVT U16018 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[464]), .B1(n11478), .B2(
        inner_first_stage_data_reg[336]), .ZN(n11418) );
  AOI22D1BWP30P140LVT U16019 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[304]), .B1(n11481), .B2(
        inner_first_stage_data_reg[496]), .ZN(n11417) );
  AOI22D1BWP30P140LVT U16020 ( .A1(n11483), .A2(
        inner_first_stage_data_reg[368]), .B1(n11482), .B2(
        inner_first_stage_data_reg[432]), .ZN(n11416) );
  ND4D1BWP30P140LVT U16021 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(N3095) );
  AOI22D1BWP30P140LVT U16022 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[273]), .B1(n11476), .B2(
        inner_first_stage_data_reg[401]), .ZN(n11423) );
  AOI22D1BWP30P140LVT U16023 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[465]), .B1(n11482), .B2(
        inner_first_stage_data_reg[433]), .ZN(n11422) );
  AOI22D1BWP30P140LVT U16024 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[305]), .B1(n11478), .B2(
        inner_first_stage_data_reg[337]), .ZN(n11421) );
  AOI22D1BWP30P140LVT U16025 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[497]), .B1(n11483), .B2(
        inner_first_stage_data_reg[369]), .ZN(n11420) );
  ND4D1BWP30P140LVT U16026 ( .A1(n11423), .A2(n11422), .A3(n11421), .A4(n11420), .ZN(N3096) );
  AOI22D1BWP30P140LVT U16027 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[274]), .B1(n11476), .B2(
        inner_first_stage_data_reg[402]), .ZN(n11427) );
  AOI22D1BWP30P140LVT U16028 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[498]), .B1(n11483), .B2(
        inner_first_stage_data_reg[370]), .ZN(n11426) );
  AOI22D1BWP30P140LVT U16029 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[466]), .B1(n11482), .B2(
        inner_first_stage_data_reg[434]), .ZN(n11425) );
  AOI22D1BWP30P140LVT U16030 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[306]), .B1(n11478), .B2(
        inner_first_stage_data_reg[338]), .ZN(n11424) );
  ND4D1BWP30P140LVT U16031 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(N3097) );
  AOI22D1BWP30P140LVT U16032 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[275]), .B1(n11476), .B2(
        inner_first_stage_data_reg[403]), .ZN(n11431) );
  AOI22D1BWP30P140LVT U16033 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[467]), .B1(n11478), .B2(
        inner_first_stage_data_reg[339]), .ZN(n11430) );
  AOI22D1BWP30P140LVT U16034 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[499]), .B1(n11482), .B2(
        inner_first_stage_data_reg[435]), .ZN(n11429) );
  AOI22D1BWP30P140LVT U16035 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[307]), .B1(n11483), .B2(
        inner_first_stage_data_reg[371]), .ZN(n11428) );
  ND4D1BWP30P140LVT U16036 ( .A1(n11431), .A2(n11430), .A3(n11429), .A4(n11428), .ZN(N3098) );
  AOI22D1BWP30P140LVT U16037 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[276]), .B1(n11476), .B2(
        inner_first_stage_data_reg[404]), .ZN(n11435) );
  AOI22D1BWP30P140LVT U16038 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[340]), .B1(n11483), .B2(
        inner_first_stage_data_reg[372]), .ZN(n11434) );
  AOI22D1BWP30P140LVT U16039 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[308]), .B1(n11482), .B2(
        inner_first_stage_data_reg[436]), .ZN(n11433) );
  AOI22D1BWP30P140LVT U16040 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[500]), .B1(n11480), .B2(
        inner_first_stage_data_reg[468]), .ZN(n11432) );
  ND4D1BWP30P140LVT U16041 ( .A1(n11435), .A2(n11434), .A3(n11433), .A4(n11432), .ZN(N3099) );
  AOI22D1BWP30P140LVT U16042 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[277]), .B1(n11476), .B2(
        inner_first_stage_data_reg[405]), .ZN(n11439) );
  AOI22D1BWP30P140LVT U16043 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[501]), .B1(n11483), .B2(
        inner_first_stage_data_reg[373]), .ZN(n11438) );
  AOI22D1BWP30P140LVT U16044 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[341]), .B1(n11482), .B2(
        inner_first_stage_data_reg[437]), .ZN(n11437) );
  AOI22D1BWP30P140LVT U16045 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[309]), .B1(n11480), .B2(
        inner_first_stage_data_reg[469]), .ZN(n11436) );
  ND4D1BWP30P140LVT U16046 ( .A1(n11439), .A2(n11438), .A3(n11437), .A4(n11436), .ZN(N3100) );
  AOI22D1BWP30P140LVT U16047 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[278]), .B1(n11476), .B2(
        inner_first_stage_data_reg[406]), .ZN(n11443) );
  AOI22D1BWP30P140LVT U16048 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[502]), .B1(n11483), .B2(
        inner_first_stage_data_reg[374]), .ZN(n11442) );
  AOI22D1BWP30P140LVT U16049 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[310]), .B1(n11478), .B2(
        inner_first_stage_data_reg[342]), .ZN(n11441) );
  AOI22D1BWP30P140LVT U16050 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[470]), .B1(n11482), .B2(
        inner_first_stage_data_reg[438]), .ZN(n11440) );
  ND4D1BWP30P140LVT U16051 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(N3101) );
  AOI22D1BWP30P140LVT U16052 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[279]), .B1(n11476), .B2(
        inner_first_stage_data_reg[407]), .ZN(n11447) );
  AOI22D1BWP30P140LVT U16053 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[311]), .B1(n11481), .B2(
        inner_first_stage_data_reg[503]), .ZN(n11446) );
  AOI22D1BWP30P140LVT U16054 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[343]), .B1(n11482), .B2(
        inner_first_stage_data_reg[439]), .ZN(n11445) );
  AOI22D1BWP30P140LVT U16055 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[471]), .B1(n11483), .B2(
        inner_first_stage_data_reg[375]), .ZN(n11444) );
  ND4D1BWP30P140LVT U16056 ( .A1(n11447), .A2(n11446), .A3(n11445), .A4(n11444), .ZN(N3102) );
  AOI22D1BWP30P140LVT U16057 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[280]), .B1(n11476), .B2(
        inner_first_stage_data_reg[408]), .ZN(n11451) );
  AOI22D1BWP30P140LVT U16058 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[344]), .B1(n11483), .B2(
        inner_first_stage_data_reg[376]), .ZN(n11450) );
  AOI22D1BWP30P140LVT U16059 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[472]), .B1(n11482), .B2(
        inner_first_stage_data_reg[440]), .ZN(n11449) );
  AOI22D1BWP30P140LVT U16060 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[312]), .B1(n11481), .B2(
        inner_first_stage_data_reg[504]), .ZN(n11448) );
  ND4D1BWP30P140LVT U16061 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(N3103) );
  AOI22D1BWP30P140LVT U16062 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[281]), .B1(n11476), .B2(
        inner_first_stage_data_reg[409]), .ZN(n11455) );
  AOI22D1BWP30P140LVT U16063 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[313]), .B1(n11480), .B2(
        inner_first_stage_data_reg[473]), .ZN(n11454) );
  AOI22D1BWP30P140LVT U16064 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[505]), .B1(n11482), .B2(
        inner_first_stage_data_reg[441]), .ZN(n11453) );
  AOI22D1BWP30P140LVT U16065 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[345]), .B1(n11483), .B2(
        inner_first_stage_data_reg[377]), .ZN(n11452) );
  ND4D1BWP30P140LVT U16066 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(N3104) );
  AOI22D1BWP30P140LVT U16067 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[282]), .B1(n11476), .B2(
        inner_first_stage_data_reg[410]), .ZN(n11459) );
  AOI22D1BWP30P140LVT U16068 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[506]), .B1(n11480), .B2(
        inner_first_stage_data_reg[474]), .ZN(n11458) );
  AOI22D1BWP30P140LVT U16069 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[346]), .B1(n11483), .B2(
        inner_first_stage_data_reg[378]), .ZN(n11457) );
  AOI22D1BWP30P140LVT U16070 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[314]), .B1(n11482), .B2(
        inner_first_stage_data_reg[442]), .ZN(n11456) );
  ND4D1BWP30P140LVT U16071 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(N3105) );
  AOI22D1BWP30P140LVT U16072 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[283]), .B1(n11476), .B2(
        inner_first_stage_data_reg[411]), .ZN(n11463) );
  AOI22D1BWP30P140LVT U16073 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[315]), .B1(n11478), .B2(
        inner_first_stage_data_reg[347]), .ZN(n11462) );
  AOI22D1BWP30P140LVT U16074 ( .A1(n11483), .A2(
        inner_first_stage_data_reg[379]), .B1(n11482), .B2(
        inner_first_stage_data_reg[443]), .ZN(n11461) );
  AOI22D1BWP30P140LVT U16075 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[507]), .B1(n11480), .B2(
        inner_first_stage_data_reg[475]), .ZN(n11460) );
  ND4D1BWP30P140LVT U16076 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(N3106) );
  AOI22D1BWP30P140LVT U16077 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[284]), .B1(n11476), .B2(
        inner_first_stage_data_reg[412]), .ZN(n11467) );
  AOI22D1BWP30P140LVT U16078 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[476]), .B1(n11482), .B2(
        inner_first_stage_data_reg[444]), .ZN(n11466) );
  AOI22D1BWP30P140LVT U16079 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[508]), .B1(n11483), .B2(
        inner_first_stage_data_reg[380]), .ZN(n11465) );
  AOI22D1BWP30P140LVT U16080 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[316]), .B1(n11478), .B2(
        inner_first_stage_data_reg[348]), .ZN(n11464) );
  ND4D1BWP30P140LVT U16081 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(N3107) );
  AOI22D1BWP30P140LVT U16082 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[285]), .B1(n11476), .B2(
        inner_first_stage_data_reg[413]), .ZN(n11471) );
  AOI22D1BWP30P140LVT U16083 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[349]), .B1(n11482), .B2(
        inner_first_stage_data_reg[445]), .ZN(n11470) );
  AOI22D1BWP30P140LVT U16084 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[317]), .B1(n11481), .B2(
        inner_first_stage_data_reg[509]), .ZN(n11469) );
  AOI22D1BWP30P140LVT U16085 ( .A1(n11480), .A2(
        inner_first_stage_data_reg[477]), .B1(n11483), .B2(
        inner_first_stage_data_reg[381]), .ZN(n11468) );
  ND4D1BWP30P140LVT U16086 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(N3108) );
  AOI22D1BWP30P140LVT U16087 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[286]), .B1(n11476), .B2(
        inner_first_stage_data_reg[414]), .ZN(n11475) );
  AOI22D1BWP30P140LVT U16088 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[318]), .B1(n11483), .B2(
        inner_first_stage_data_reg[382]), .ZN(n11474) );
  AOI22D1BWP30P140LVT U16089 ( .A1(n11478), .A2(
        inner_first_stage_data_reg[350]), .B1(n11482), .B2(
        inner_first_stage_data_reg[446]), .ZN(n11473) );
  AOI22D1BWP30P140LVT U16090 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[510]), .B1(n11480), .B2(
        inner_first_stage_data_reg[478]), .ZN(n11472) );
  ND4D1BWP30P140LVT U16091 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(N3109) );
  AOI22D1BWP30P140LVT U16092 ( .A1(n11477), .A2(
        inner_first_stage_data_reg[287]), .B1(n11476), .B2(
        inner_first_stage_data_reg[415]), .ZN(n11487) );
  AOI22D1BWP30P140LVT U16093 ( .A1(n11479), .A2(
        inner_first_stage_data_reg[319]), .B1(n11478), .B2(
        inner_first_stage_data_reg[351]), .ZN(n11486) );
  AOI22D1BWP30P140LVT U16094 ( .A1(n11481), .A2(
        inner_first_stage_data_reg[511]), .B1(n11480), .B2(
        inner_first_stage_data_reg[479]), .ZN(n11485) );
  AOI22D1BWP30P140LVT U16095 ( .A1(n11483), .A2(
        inner_first_stage_data_reg[383]), .B1(n11482), .B2(
        inner_first_stage_data_reg[447]), .ZN(n11484) );
  ND4D1BWP30P140LVT U16096 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(N3110) );
  AOI22D1BWP30P140LVT U16097 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[672]), .B1(n11613), .B2(
        inner_first_stage_data_reg[512]), .ZN(n11491) );
  AOI22D1BWP30P140LVT U16098 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[640]), .B1(n11612), .B2(
        inner_first_stage_data_reg[544]), .ZN(n11490) );
  AOI22D1BWP30P140LVT U16099 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[704]), .B1(n11619), .B2(
        inner_first_stage_data_reg[736]), .ZN(n11489) );
  AOI22D1BWP30P140LVT U16100 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[576]), .B1(n11618), .B2(
        inner_first_stage_data_reg[608]), .ZN(n11488) );
  ND4D1BWP30P140LVT U16101 ( .A1(n11491), .A2(n11490), .A3(n11489), .A4(n11488), .ZN(N4953) );
  AOI22D1BWP30P140LVT U16102 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[513]), .B1(n11612), .B2(
        inner_first_stage_data_reg[545]), .ZN(n11495) );
  AOI22D1BWP30P140LVT U16103 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[673]), .B1(n11614), .B2(
        inner_first_stage_data_reg[641]), .ZN(n11494) );
  AOI22D1BWP30P140LVT U16104 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[737]), .B1(n11618), .B2(
        inner_first_stage_data_reg[609]), .ZN(n11493) );
  AOI22D1BWP30P140LVT U16105 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[705]), .B1(n11616), .B2(
        inner_first_stage_data_reg[577]), .ZN(n11492) );
  ND4D1BWP30P140LVT U16106 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(N4954) );
  AOI22D1BWP30P140LVT U16107 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[674]), .B1(n11614), .B2(
        inner_first_stage_data_reg[642]), .ZN(n11499) );
  AOI22D1BWP30P140LVT U16108 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[514]), .B1(n11612), .B2(
        inner_first_stage_data_reg[546]), .ZN(n11498) );
  AOI22D1BWP30P140LVT U16109 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[738]), .B1(n11616), .B2(
        inner_first_stage_data_reg[578]), .ZN(n11497) );
  AOI22D1BWP30P140LVT U16110 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[706]), .B1(n11618), .B2(
        inner_first_stage_data_reg[610]), .ZN(n11496) );
  ND4D1BWP30P140LVT U16111 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(N4955) );
  AOI22D1BWP30P140LVT U16112 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[675]), .B1(n11613), .B2(
        inner_first_stage_data_reg[515]), .ZN(n11503) );
  AOI22D1BWP30P140LVT U16113 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[643]), .B1(n11612), .B2(
        inner_first_stage_data_reg[547]), .ZN(n11502) );
  AOI22D1BWP30P140LVT U16114 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[707]), .B1(n11616), .B2(
        inner_first_stage_data_reg[579]), .ZN(n11501) );
  AOI22D1BWP30P140LVT U16115 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[739]), .B1(n11618), .B2(
        inner_first_stage_data_reg[611]), .ZN(n11500) );
  ND4D1BWP30P140LVT U16116 ( .A1(n11503), .A2(n11502), .A3(n11501), .A4(n11500), .ZN(N4956) );
  AOI22D1BWP30P140LVT U16117 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[644]), .B1(n11612), .B2(
        inner_first_stage_data_reg[548]), .ZN(n11507) );
  AOI22D1BWP30P140LVT U16118 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[676]), .B1(n11613), .B2(
        inner_first_stage_data_reg[516]), .ZN(n11506) );
  AOI22D1BWP30P140LVT U16119 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[740]), .B1(n11616), .B2(
        inner_first_stage_data_reg[580]), .ZN(n11505) );
  AOI22D1BWP30P140LVT U16120 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[708]), .B1(n11618), .B2(
        inner_first_stage_data_reg[612]), .ZN(n11504) );
  ND4D1BWP30P140LVT U16121 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(N4957) );
  AOI22D1BWP30P140LVT U16122 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[677]), .B1(n11612), .B2(
        inner_first_stage_data_reg[549]), .ZN(n11511) );
  AOI22D1BWP30P140LVT U16123 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[517]), .B1(n11614), .B2(
        inner_first_stage_data_reg[645]), .ZN(n11510) );
  AOI22D1BWP30P140LVT U16124 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[709]), .B1(n11619), .B2(
        inner_first_stage_data_reg[741]), .ZN(n11509) );
  AOI22D1BWP30P140LVT U16125 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[581]), .B1(n11618), .B2(
        inner_first_stage_data_reg[613]), .ZN(n11508) );
  ND4D1BWP30P140LVT U16126 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(N4958) );
  AOI22D1BWP30P140LVT U16127 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[646]), .B1(n11612), .B2(
        inner_first_stage_data_reg[550]), .ZN(n11515) );
  AOI22D1BWP30P140LVT U16128 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[678]), .B1(n11613), .B2(
        inner_first_stage_data_reg[518]), .ZN(n11514) );
  AOI22D1BWP30P140LVT U16129 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[582]), .B1(n11618), .B2(
        inner_first_stage_data_reg[614]), .ZN(n11513) );
  AOI22D1BWP30P140LVT U16130 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[710]), .B1(n11619), .B2(
        inner_first_stage_data_reg[742]), .ZN(n11512) );
  ND4D1BWP30P140LVT U16131 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(N4959) );
  AOI22D1BWP30P140LVT U16132 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[679]), .B1(n11613), .B2(
        inner_first_stage_data_reg[519]), .ZN(n11519) );
  AOI22D1BWP30P140LVT U16133 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[647]), .B1(n11612), .B2(
        inner_first_stage_data_reg[551]), .ZN(n11518) );
  AOI22D1BWP30P140LVT U16134 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[711]), .B1(n11618), .B2(
        inner_first_stage_data_reg[615]), .ZN(n11517) );
  AOI22D1BWP30P140LVT U16135 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[743]), .B1(n11616), .B2(
        inner_first_stage_data_reg[583]), .ZN(n11516) );
  ND4D1BWP30P140LVT U16136 ( .A1(n11519), .A2(n11518), .A3(n11517), .A4(n11516), .ZN(N4960) );
  AOI22D1BWP30P140LVT U16137 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[648]), .B1(n11612), .B2(
        inner_first_stage_data_reg[552]), .ZN(n11523) );
  AOI22D1BWP30P140LVT U16138 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[680]), .B1(n11613), .B2(
        inner_first_stage_data_reg[520]), .ZN(n11522) );
  AOI22D1BWP30P140LVT U16139 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[712]), .B1(n11618), .B2(
        inner_first_stage_data_reg[616]), .ZN(n11521) );
  AOI22D1BWP30P140LVT U16140 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[744]), .B1(n11616), .B2(
        inner_first_stage_data_reg[584]), .ZN(n11520) );
  ND4D1BWP30P140LVT U16141 ( .A1(n11523), .A2(n11522), .A3(n11521), .A4(n11520), .ZN(N4961) );
  AOI22D1BWP30P140LVT U16142 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[681]), .B1(n11613), .B2(
        inner_first_stage_data_reg[521]), .ZN(n11527) );
  AOI22D1BWP30P140LVT U16143 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[649]), .B1(n11612), .B2(
        inner_first_stage_data_reg[553]), .ZN(n11526) );
  AOI22D1BWP30P140LVT U16144 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[713]), .B1(n11616), .B2(
        inner_first_stage_data_reg[585]), .ZN(n11525) );
  AOI22D1BWP30P140LVT U16145 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[745]), .B1(n11618), .B2(
        inner_first_stage_data_reg[617]), .ZN(n11524) );
  ND4D1BWP30P140LVT U16146 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(N4962) );
  AOI22D1BWP30P140LVT U16147 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[682]), .B1(n11614), .B2(
        inner_first_stage_data_reg[650]), .ZN(n11531) );
  AOI22D1BWP30P140LVT U16148 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[522]), .B1(n11612), .B2(
        inner_first_stage_data_reg[554]), .ZN(n11530) );
  AOI22D1BWP30P140LVT U16149 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[714]), .B1(n11619), .B2(
        inner_first_stage_data_reg[746]), .ZN(n11529) );
  AOI22D1BWP30P140LVT U16150 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[586]), .B1(n11618), .B2(
        inner_first_stage_data_reg[618]), .ZN(n11528) );
  ND4D1BWP30P140LVT U16151 ( .A1(n11531), .A2(n11530), .A3(n11529), .A4(n11528), .ZN(N4963) );
  AOI22D1BWP30P140LVT U16152 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[523]), .B1(n11612), .B2(
        inner_first_stage_data_reg[555]), .ZN(n11535) );
  AOI22D1BWP30P140LVT U16153 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[683]), .B1(n11614), .B2(
        inner_first_stage_data_reg[651]), .ZN(n11534) );
  AOI22D1BWP30P140LVT U16154 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[587]), .B1(n11618), .B2(
        inner_first_stage_data_reg[619]), .ZN(n11533) );
  AOI22D1BWP30P140LVT U16155 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[715]), .B1(n11619), .B2(
        inner_first_stage_data_reg[747]), .ZN(n11532) );
  ND4D1BWP30P140LVT U16156 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(N4964) );
  AOI22D1BWP30P140LVT U16157 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[684]), .B1(n11613), .B2(
        inner_first_stage_data_reg[524]), .ZN(n11539) );
  AOI22D1BWP30P140LVT U16158 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[652]), .B1(n11612), .B2(
        inner_first_stage_data_reg[556]), .ZN(n11538) );
  AOI22D1BWP30P140LVT U16159 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[748]), .B1(n11618), .B2(
        inner_first_stage_data_reg[620]), .ZN(n11537) );
  AOI22D1BWP30P140LVT U16160 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[716]), .B1(n11616), .B2(
        inner_first_stage_data_reg[588]), .ZN(n11536) );
  ND4D1BWP30P140LVT U16161 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(N4965) );
  AOI22D1BWP30P140LVT U16162 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[685]), .B1(n11614), .B2(
        inner_first_stage_data_reg[653]), .ZN(n11543) );
  AOI22D1BWP30P140LVT U16163 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[525]), .B1(n11612), .B2(
        inner_first_stage_data_reg[557]), .ZN(n11542) );
  AOI22D1BWP30P140LVT U16164 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[589]), .B1(n11618), .B2(
        inner_first_stage_data_reg[621]), .ZN(n11541) );
  AOI22D1BWP30P140LVT U16165 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[717]), .B1(n11619), .B2(
        inner_first_stage_data_reg[749]), .ZN(n11540) );
  ND4D1BWP30P140LVT U16166 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(N4966) );
  AOI22D1BWP30P140LVT U16167 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[686]), .B1(n11614), .B2(
        inner_first_stage_data_reg[654]), .ZN(n11547) );
  AOI22D1BWP30P140LVT U16168 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[526]), .B1(n11612), .B2(
        inner_first_stage_data_reg[558]), .ZN(n11546) );
  AOI22D1BWP30P140LVT U16169 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[718]), .B1(n11618), .B2(
        inner_first_stage_data_reg[622]), .ZN(n11545) );
  AOI22D1BWP30P140LVT U16170 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[750]), .B1(n11616), .B2(
        inner_first_stage_data_reg[590]), .ZN(n11544) );
  ND4D1BWP30P140LVT U16171 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(N4967) );
  AOI22D1BWP30P140LVT U16172 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[527]), .B1(n11612), .B2(
        inner_first_stage_data_reg[559]), .ZN(n11551) );
  AOI22D1BWP30P140LVT U16173 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[687]), .B1(n11614), .B2(
        inner_first_stage_data_reg[655]), .ZN(n11550) );
  AOI22D1BWP30P140LVT U16174 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[591]), .B1(n11618), .B2(
        inner_first_stage_data_reg[623]), .ZN(n11549) );
  AOI22D1BWP30P140LVT U16175 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[719]), .B1(n11619), .B2(
        inner_first_stage_data_reg[751]), .ZN(n11548) );
  ND4D1BWP30P140LVT U16176 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(N4968) );
  AOI22D1BWP30P140LVT U16177 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[656]), .B1(n11612), .B2(
        inner_first_stage_data_reg[560]), .ZN(n11555) );
  AOI22D1BWP30P140LVT U16178 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[688]), .B1(n11613), .B2(
        inner_first_stage_data_reg[528]), .ZN(n11554) );
  AOI22D1BWP30P140LVT U16179 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[592]), .B1(n11618), .B2(
        inner_first_stage_data_reg[624]), .ZN(n11553) );
  AOI22D1BWP30P140LVT U16180 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[720]), .B1(n11619), .B2(
        inner_first_stage_data_reg[752]), .ZN(n11552) );
  ND4D1BWP30P140LVT U16181 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(N4969) );
  AOI22D1BWP30P140LVT U16182 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[657]), .B1(n11612), .B2(
        inner_first_stage_data_reg[561]), .ZN(n11559) );
  AOI22D1BWP30P140LVT U16183 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[689]), .B1(n11613), .B2(
        inner_first_stage_data_reg[529]), .ZN(n11558) );
  AOI22D1BWP30P140LVT U16184 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[753]), .B1(n11616), .B2(
        inner_first_stage_data_reg[593]), .ZN(n11557) );
  AOI22D1BWP30P140LVT U16185 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[721]), .B1(n11618), .B2(
        inner_first_stage_data_reg[625]), .ZN(n11556) );
  ND4D1BWP30P140LVT U16186 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(N4970) );
  AOI22D1BWP30P140LVT U16187 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[690]), .B1(n11613), .B2(
        inner_first_stage_data_reg[530]), .ZN(n11563) );
  AOI22D1BWP30P140LVT U16188 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[658]), .B1(n11612), .B2(
        inner_first_stage_data_reg[562]), .ZN(n11562) );
  AOI22D1BWP30P140LVT U16189 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[754]), .B1(n11618), .B2(
        inner_first_stage_data_reg[626]), .ZN(n11561) );
  AOI22D1BWP30P140LVT U16190 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[722]), .B1(n11616), .B2(
        inner_first_stage_data_reg[594]), .ZN(n11560) );
  ND4D1BWP30P140LVT U16191 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(N4971) );
  AOI22D1BWP30P140LVT U16192 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[691]), .B1(n11613), .B2(
        inner_first_stage_data_reg[531]), .ZN(n11567) );
  AOI22D1BWP30P140LVT U16193 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[659]), .B1(n11612), .B2(
        inner_first_stage_data_reg[563]), .ZN(n11566) );
  AOI22D1BWP30P140LVT U16194 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[723]), .B1(n11616), .B2(
        inner_first_stage_data_reg[595]), .ZN(n11565) );
  AOI22D1BWP30P140LVT U16195 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[755]), .B1(n11618), .B2(
        inner_first_stage_data_reg[627]), .ZN(n11564) );
  ND4D1BWP30P140LVT U16196 ( .A1(n11567), .A2(n11566), .A3(n11565), .A4(n11564), .ZN(N4972) );
  AOI22D1BWP30P140LVT U16197 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[532]), .B1(n11612), .B2(
        inner_first_stage_data_reg[564]), .ZN(n11571) );
  AOI22D1BWP30P140LVT U16198 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[692]), .B1(n11614), .B2(
        inner_first_stage_data_reg[660]), .ZN(n11570) );
  AOI22D1BWP30P140LVT U16199 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[724]), .B1(n11619), .B2(
        inner_first_stage_data_reg[756]), .ZN(n11569) );
  AOI22D1BWP30P140LVT U16200 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[596]), .B1(n11618), .B2(
        inner_first_stage_data_reg[628]), .ZN(n11568) );
  ND4D1BWP30P140LVT U16201 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(N4973) );
  AOI22D1BWP30P140LVT U16202 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[533]), .B1(n11612), .B2(
        inner_first_stage_data_reg[565]), .ZN(n11575) );
  AOI22D1BWP30P140LVT U16203 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[693]), .B1(n11614), .B2(
        inner_first_stage_data_reg[661]), .ZN(n11574) );
  AOI22D1BWP30P140LVT U16204 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[725]), .B1(n11618), .B2(
        inner_first_stage_data_reg[629]), .ZN(n11573) );
  AOI22D1BWP30P140LVT U16205 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[757]), .B1(n11616), .B2(
        inner_first_stage_data_reg[597]), .ZN(n11572) );
  ND4D1BWP30P140LVT U16206 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(N4974) );
  AOI22D1BWP30P140LVT U16207 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[534]), .B1(n11614), .B2(
        inner_first_stage_data_reg[662]), .ZN(n11579) );
  AOI22D1BWP30P140LVT U16208 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[694]), .B1(n11612), .B2(
        inner_first_stage_data_reg[566]), .ZN(n11578) );
  AOI22D1BWP30P140LVT U16209 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[758]), .B1(n11616), .B2(
        inner_first_stage_data_reg[598]), .ZN(n11577) );
  AOI22D1BWP30P140LVT U16210 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[726]), .B1(n11618), .B2(
        inner_first_stage_data_reg[630]), .ZN(n11576) );
  ND4D1BWP30P140LVT U16211 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(N4975) );
  AOI22D1BWP30P140LVT U16212 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[695]), .B1(n11614), .B2(
        inner_first_stage_data_reg[663]), .ZN(n11583) );
  AOI22D1BWP30P140LVT U16213 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[535]), .B1(n11612), .B2(
        inner_first_stage_data_reg[567]), .ZN(n11582) );
  AOI22D1BWP30P140LVT U16214 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[727]), .B1(n11619), .B2(
        inner_first_stage_data_reg[759]), .ZN(n11581) );
  AOI22D1BWP30P140LVT U16215 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[599]), .B1(n11618), .B2(
        inner_first_stage_data_reg[631]), .ZN(n11580) );
  ND4D1BWP30P140LVT U16216 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(N4976) );
  AOI22D1BWP30P140LVT U16217 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[696]), .B1(n11612), .B2(
        inner_first_stage_data_reg[568]), .ZN(n11587) );
  AOI22D1BWP30P140LVT U16218 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[536]), .B1(n11614), .B2(
        inner_first_stage_data_reg[664]), .ZN(n11586) );
  AOI22D1BWP30P140LVT U16219 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[760]), .B1(n11618), .B2(
        inner_first_stage_data_reg[632]), .ZN(n11585) );
  AOI22D1BWP30P140LVT U16220 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[728]), .B1(n11616), .B2(
        inner_first_stage_data_reg[600]), .ZN(n11584) );
  ND4D1BWP30P140LVT U16221 ( .A1(n11587), .A2(n11586), .A3(n11585), .A4(n11584), .ZN(N4977) );
  AOI22D1BWP30P140LVT U16222 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[537]), .B1(n11612), .B2(
        inner_first_stage_data_reg[569]), .ZN(n11591) );
  AOI22D1BWP30P140LVT U16223 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[697]), .B1(n11614), .B2(
        inner_first_stage_data_reg[665]), .ZN(n11590) );
  AOI22D1BWP30P140LVT U16224 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[729]), .B1(n11616), .B2(
        inner_first_stage_data_reg[601]), .ZN(n11589) );
  AOI22D1BWP30P140LVT U16225 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[761]), .B1(n11618), .B2(
        inner_first_stage_data_reg[633]), .ZN(n11588) );
  ND4D1BWP30P140LVT U16226 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(N4978) );
  AOI22D1BWP30P140LVT U16227 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[538]), .B1(n11612), .B2(
        inner_first_stage_data_reg[570]), .ZN(n11595) );
  AOI22D1BWP30P140LVT U16228 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[698]), .B1(n11614), .B2(
        inner_first_stage_data_reg[666]), .ZN(n11594) );
  AOI22D1BWP30P140LVT U16229 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[730]), .B1(n11618), .B2(
        inner_first_stage_data_reg[634]), .ZN(n11593) );
  AOI22D1BWP30P140LVT U16230 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[762]), .B1(n11616), .B2(
        inner_first_stage_data_reg[602]), .ZN(n11592) );
  ND4D1BWP30P140LVT U16231 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(N4979) );
  AOI22D1BWP30P140LVT U16232 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[539]), .B1(n11614), .B2(
        inner_first_stage_data_reg[667]), .ZN(n11599) );
  AOI22D1BWP30P140LVT U16233 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[699]), .B1(n11612), .B2(
        inner_first_stage_data_reg[571]), .ZN(n11598) );
  AOI22D1BWP30P140LVT U16234 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[731]), .B1(n11619), .B2(
        inner_first_stage_data_reg[763]), .ZN(n11597) );
  AOI22D1BWP30P140LVT U16235 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[603]), .B1(n11618), .B2(
        inner_first_stage_data_reg[635]), .ZN(n11596) );
  ND4D1BWP30P140LVT U16236 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(N4980) );
  AOI22D1BWP30P140LVT U16237 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[540]), .B1(n11612), .B2(
        inner_first_stage_data_reg[572]), .ZN(n11603) );
  AOI22D1BWP30P140LVT U16238 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[700]), .B1(n11614), .B2(
        inner_first_stage_data_reg[668]), .ZN(n11602) );
  AOI22D1BWP30P140LVT U16239 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[604]), .B1(n11618), .B2(
        inner_first_stage_data_reg[636]), .ZN(n11601) );
  AOI22D1BWP30P140LVT U16240 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[732]), .B1(n11619), .B2(
        inner_first_stage_data_reg[764]), .ZN(n11600) );
  ND4D1BWP30P140LVT U16241 ( .A1(n11603), .A2(n11602), .A3(n11601), .A4(n11600), .ZN(N4981) );
  AOI22D1BWP30P140LVT U16242 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[701]), .B1(n11613), .B2(
        inner_first_stage_data_reg[541]), .ZN(n11607) );
  AOI22D1BWP30P140LVT U16243 ( .A1(n11614), .A2(
        inner_first_stage_data_reg[669]), .B1(n11612), .B2(
        inner_first_stage_data_reg[573]), .ZN(n11606) );
  AOI22D1BWP30P140LVT U16244 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[733]), .B1(n11619), .B2(
        inner_first_stage_data_reg[765]), .ZN(n11605) );
  AOI22D1BWP30P140LVT U16245 ( .A1(n11616), .A2(
        inner_first_stage_data_reg[605]), .B1(n11618), .B2(
        inner_first_stage_data_reg[637]), .ZN(n11604) );
  ND4D1BWP30P140LVT U16246 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(N4982) );
  AOI22D1BWP30P140LVT U16247 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[702]), .B1(n11612), .B2(
        inner_first_stage_data_reg[574]), .ZN(n11611) );
  AOI22D1BWP30P140LVT U16248 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[542]), .B1(n11614), .B2(
        inner_first_stage_data_reg[670]), .ZN(n11610) );
  AOI22D1BWP30P140LVT U16249 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[766]), .B1(n11618), .B2(
        inner_first_stage_data_reg[638]), .ZN(n11609) );
  AOI22D1BWP30P140LVT U16250 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[734]), .B1(n11616), .B2(
        inner_first_stage_data_reg[606]), .ZN(n11608) );
  ND4D1BWP30P140LVT U16251 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(N4983) );
  AOI22D1BWP30P140LVT U16252 ( .A1(n11613), .A2(
        inner_first_stage_data_reg[543]), .B1(n11612), .B2(
        inner_first_stage_data_reg[575]), .ZN(n11623) );
  AOI22D1BWP30P140LVT U16253 ( .A1(n11615), .A2(
        inner_first_stage_data_reg[703]), .B1(n11614), .B2(
        inner_first_stage_data_reg[671]), .ZN(n11622) );
  AOI22D1BWP30P140LVT U16254 ( .A1(n11617), .A2(
        inner_first_stage_data_reg[735]), .B1(n11616), .B2(
        inner_first_stage_data_reg[607]), .ZN(n11621) );
  AOI22D1BWP30P140LVT U16255 ( .A1(n11619), .A2(
        inner_first_stage_data_reg[767]), .B1(n11618), .B2(
        inner_first_stage_data_reg[639]), .ZN(n11620) );
  ND4D1BWP30P140LVT U16256 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(N4984) );
  AOI22D1BWP30P140LVT U16257 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[992]), .B1(n11748), .B2(
        inner_first_stage_data_reg[960]), .ZN(n11627) );
  AOI22D1BWP30P140LVT U16258 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[768]), .B1(n11750), .B2(
        inner_first_stage_data_reg[896]), .ZN(n11626) );
  AOI22D1BWP30P140LVT U16259 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[800]), .B1(n11753), .B2(
        inner_first_stage_data_reg[928]), .ZN(n11625) );
  AOI22D1BWP30P140LVT U16260 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[832]), .B1(n11752), .B2(
        inner_first_stage_data_reg[864]), .ZN(n11624) );
  ND4D1BWP30P140LVT U16261 ( .A1(n11627), .A2(n11626), .A3(n11625), .A4(n11624), .ZN(N5803) );
  AOI22D1BWP30P140LVT U16262 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[993]), .B1(n11750), .B2(
        inner_first_stage_data_reg[897]), .ZN(n11631) );
  AOI22D1BWP30P140LVT U16263 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[961]), .B1(n11751), .B2(
        inner_first_stage_data_reg[769]), .ZN(n11630) );
  AOI22D1BWP30P140LVT U16264 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[929]), .B1(n11752), .B2(
        inner_first_stage_data_reg[865]), .ZN(n11629) );
  AOI22D1BWP30P140LVT U16265 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[801]), .B1(n11754), .B2(
        inner_first_stage_data_reg[833]), .ZN(n11628) );
  ND4D1BWP30P140LVT U16266 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(N5804) );
  AOI22D1BWP30P140LVT U16267 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[994]), .B1(n11751), .B2(
        inner_first_stage_data_reg[770]), .ZN(n11635) );
  AOI22D1BWP30P140LVT U16268 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[962]), .B1(n11750), .B2(
        inner_first_stage_data_reg[898]), .ZN(n11634) );
  AOI22D1BWP30P140LVT U16269 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[834]), .B1(n11752), .B2(
        inner_first_stage_data_reg[866]), .ZN(n11633) );
  AOI22D1BWP30P140LVT U16270 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[802]), .B1(n11753), .B2(
        inner_first_stage_data_reg[930]), .ZN(n11632) );
  ND4D1BWP30P140LVT U16271 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(N5805) );
  AOI22D1BWP30P140LVT U16272 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[963]), .B1(n11751), .B2(
        inner_first_stage_data_reg[771]), .ZN(n11639) );
  AOI22D1BWP30P140LVT U16273 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[995]), .B1(n11750), .B2(
        inner_first_stage_data_reg[899]), .ZN(n11638) );
  AOI22D1BWP30P140LVT U16274 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[835]), .B1(n11752), .B2(
        inner_first_stage_data_reg[867]), .ZN(n11637) );
  AOI22D1BWP30P140LVT U16275 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[803]), .B1(n11753), .B2(
        inner_first_stage_data_reg[931]), .ZN(n11636) );
  ND4D1BWP30P140LVT U16276 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(N5806) );
  AOI22D1BWP30P140LVT U16277 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[772]), .B1(n11750), .B2(
        inner_first_stage_data_reg[900]), .ZN(n11643) );
  AOI22D1BWP30P140LVT U16278 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[996]), .B1(n11748), .B2(
        inner_first_stage_data_reg[964]), .ZN(n11642) );
  AOI22D1BWP30P140LVT U16279 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[804]), .B1(n11752), .B2(
        inner_first_stage_data_reg[868]), .ZN(n11641) );
  AOI22D1BWP30P140LVT U16280 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[932]), .B1(n11754), .B2(
        inner_first_stage_data_reg[836]), .ZN(n11640) );
  ND4D1BWP30P140LVT U16281 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(N5807) );
  AOI22D1BWP30P140LVT U16282 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[773]), .B1(n11750), .B2(
        inner_first_stage_data_reg[901]), .ZN(n11647) );
  AOI22D1BWP30P140LVT U16283 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[997]), .B1(n11748), .B2(
        inner_first_stage_data_reg[965]), .ZN(n11646) );
  AOI22D1BWP30P140LVT U16284 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[805]), .B1(n11752), .B2(
        inner_first_stage_data_reg[869]), .ZN(n11645) );
  AOI22D1BWP30P140LVT U16285 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[933]), .B1(n11754), .B2(
        inner_first_stage_data_reg[837]), .ZN(n11644) );
  ND4D1BWP30P140LVT U16286 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(N5808) );
  AOI22D1BWP30P140LVT U16287 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[966]), .B1(n11751), .B2(
        inner_first_stage_data_reg[774]), .ZN(n11651) );
  AOI22D1BWP30P140LVT U16288 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[998]), .B1(n11750), .B2(
        inner_first_stage_data_reg[902]), .ZN(n11650) );
  AOI22D1BWP30P140LVT U16289 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[806]), .B1(n11752), .B2(
        inner_first_stage_data_reg[870]), .ZN(n11649) );
  AOI22D1BWP30P140LVT U16290 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[934]), .B1(n11754), .B2(
        inner_first_stage_data_reg[838]), .ZN(n11648) );
  ND4D1BWP30P140LVT U16291 ( .A1(n11651), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(N5809) );
  AOI22D1BWP30P140LVT U16292 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[775]), .B1(n11750), .B2(
        inner_first_stage_data_reg[903]), .ZN(n11655) );
  AOI22D1BWP30P140LVT U16293 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[999]), .B1(n11748), .B2(
        inner_first_stage_data_reg[967]), .ZN(n11654) );
  AOI22D1BWP30P140LVT U16294 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[935]), .B1(n11752), .B2(
        inner_first_stage_data_reg[871]), .ZN(n11653) );
  AOI22D1BWP30P140LVT U16295 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[807]), .B1(n11754), .B2(
        inner_first_stage_data_reg[839]), .ZN(n11652) );
  ND4D1BWP30P140LVT U16296 ( .A1(n11655), .A2(n11654), .A3(n11653), .A4(n11652), .ZN(N5810) );
  AOI22D1BWP30P140LVT U16297 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1000]), .B1(n11750), .B2(
        inner_first_stage_data_reg[904]), .ZN(n11659) );
  AOI22D1BWP30P140LVT U16298 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[968]), .B1(n11751), .B2(
        inner_first_stage_data_reg[776]), .ZN(n11658) );
  AOI22D1BWP30P140LVT U16299 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[936]), .B1(n11752), .B2(
        inner_first_stage_data_reg[872]), .ZN(n11657) );
  AOI22D1BWP30P140LVT U16300 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[808]), .B1(n11754), .B2(
        inner_first_stage_data_reg[840]), .ZN(n11656) );
  ND4D1BWP30P140LVT U16301 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(N5811) );
  AOI22D1BWP30P140LVT U16302 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1001]), .B1(n11751), .B2(
        inner_first_stage_data_reg[777]), .ZN(n11663) );
  AOI22D1BWP30P140LVT U16303 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[969]), .B1(n11750), .B2(
        inner_first_stage_data_reg[905]), .ZN(n11662) );
  AOI22D1BWP30P140LVT U16304 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[841]), .B1(n11752), .B2(
        inner_first_stage_data_reg[873]), .ZN(n11661) );
  AOI22D1BWP30P140LVT U16305 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[809]), .B1(n11753), .B2(
        inner_first_stage_data_reg[937]), .ZN(n11660) );
  ND4D1BWP30P140LVT U16306 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(N5812) );
  AOI22D1BWP30P140LVT U16307 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1002]), .B1(n11751), .B2(
        inner_first_stage_data_reg[778]), .ZN(n11667) );
  AOI22D1BWP30P140LVT U16308 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[970]), .B1(n11750), .B2(
        inner_first_stage_data_reg[906]), .ZN(n11666) );
  AOI22D1BWP30P140LVT U16309 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[810]), .B1(n11752), .B2(
        inner_first_stage_data_reg[874]), .ZN(n11665) );
  AOI22D1BWP30P140LVT U16310 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[938]), .B1(n11754), .B2(
        inner_first_stage_data_reg[842]), .ZN(n11664) );
  ND4D1BWP30P140LVT U16311 ( .A1(n11667), .A2(n11666), .A3(n11665), .A4(n11664), .ZN(N5813) );
  AOI22D1BWP30P140LVT U16312 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1003]), .B1(n11751), .B2(
        inner_first_stage_data_reg[779]), .ZN(n11671) );
  AOI22D1BWP30P140LVT U16313 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[971]), .B1(n11750), .B2(
        inner_first_stage_data_reg[907]), .ZN(n11670) );
  AOI22D1BWP30P140LVT U16314 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[811]), .B1(n11754), .B2(
        inner_first_stage_data_reg[843]), .ZN(n11669) );
  AOI22D1BWP30P140LVT U16315 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[939]), .B1(n11752), .B2(
        inner_first_stage_data_reg[875]), .ZN(n11668) );
  ND4D1BWP30P140LVT U16316 ( .A1(n11671), .A2(n11670), .A3(n11669), .A4(n11668), .ZN(N5814) );
  AOI22D1BWP30P140LVT U16317 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[780]), .B1(n11750), .B2(
        inner_first_stage_data_reg[908]), .ZN(n11675) );
  AOI22D1BWP30P140LVT U16318 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1004]), .B1(n11748), .B2(
        inner_first_stage_data_reg[972]), .ZN(n11674) );
  AOI22D1BWP30P140LVT U16319 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[844]), .B1(n11752), .B2(
        inner_first_stage_data_reg[876]), .ZN(n11673) );
  AOI22D1BWP30P140LVT U16320 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[812]), .B1(n11753), .B2(
        inner_first_stage_data_reg[940]), .ZN(n11672) );
  ND4D1BWP30P140LVT U16321 ( .A1(n11675), .A2(n11674), .A3(n11673), .A4(n11672), .ZN(N5815) );
  AOI22D1BWP30P140LVT U16322 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1005]), .B1(n11751), .B2(
        inner_first_stage_data_reg[781]), .ZN(n11679) );
  AOI22D1BWP30P140LVT U16323 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[973]), .B1(n11750), .B2(
        inner_first_stage_data_reg[909]), .ZN(n11678) );
  AOI22D1BWP30P140LVT U16324 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[813]), .B1(n11754), .B2(
        inner_first_stage_data_reg[845]), .ZN(n11677) );
  AOI22D1BWP30P140LVT U16325 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[941]), .B1(n11752), .B2(
        inner_first_stage_data_reg[877]), .ZN(n11676) );
  ND4D1BWP30P140LVT U16326 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(N5816) );
  AOI22D1BWP30P140LVT U16327 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1006]), .B1(n11750), .B2(
        inner_first_stage_data_reg[910]), .ZN(n11683) );
  AOI22D1BWP30P140LVT U16328 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[974]), .B1(n11751), .B2(
        inner_first_stage_data_reg[782]), .ZN(n11682) );
  AOI22D1BWP30P140LVT U16329 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[942]), .B1(n11754), .B2(
        inner_first_stage_data_reg[846]), .ZN(n11681) );
  AOI22D1BWP30P140LVT U16330 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[814]), .B1(n11752), .B2(
        inner_first_stage_data_reg[878]), .ZN(n11680) );
  ND4D1BWP30P140LVT U16331 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(N5817) );
  AOI22D1BWP30P140LVT U16332 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1007]), .B1(n11748), .B2(
        inner_first_stage_data_reg[975]), .ZN(n11687) );
  AOI22D1BWP30P140LVT U16333 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[783]), .B1(n11750), .B2(
        inner_first_stage_data_reg[911]), .ZN(n11686) );
  AOI22D1BWP30P140LVT U16334 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[847]), .B1(n11752), .B2(
        inner_first_stage_data_reg[879]), .ZN(n11685) );
  AOI22D1BWP30P140LVT U16335 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[815]), .B1(n11753), .B2(
        inner_first_stage_data_reg[943]), .ZN(n11684) );
  ND4D1BWP30P140LVT U16336 ( .A1(n11687), .A2(n11686), .A3(n11685), .A4(n11684), .ZN(N5818) );
  AOI22D1BWP30P140LVT U16337 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[976]), .B1(n11751), .B2(
        inner_first_stage_data_reg[784]), .ZN(n11691) );
  AOI22D1BWP30P140LVT U16338 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1008]), .B1(n11750), .B2(
        inner_first_stage_data_reg[912]), .ZN(n11690) );
  AOI22D1BWP30P140LVT U16339 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[944]), .B1(n11752), .B2(
        inner_first_stage_data_reg[880]), .ZN(n11689) );
  AOI22D1BWP30P140LVT U16340 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[816]), .B1(n11754), .B2(
        inner_first_stage_data_reg[848]), .ZN(n11688) );
  ND4D1BWP30P140LVT U16341 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(N5819) );
  AOI22D1BWP30P140LVT U16342 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1009]), .B1(n11748), .B2(
        inner_first_stage_data_reg[977]), .ZN(n11695) );
  AOI22D1BWP30P140LVT U16343 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[785]), .B1(n11750), .B2(
        inner_first_stage_data_reg[913]), .ZN(n11694) );
  AOI22D1BWP30P140LVT U16344 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[817]), .B1(n11753), .B2(
        inner_first_stage_data_reg[945]), .ZN(n11693) );
  AOI22D1BWP30P140LVT U16345 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[849]), .B1(n11752), .B2(
        inner_first_stage_data_reg[881]), .ZN(n11692) );
  ND4D1BWP30P140LVT U16346 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(N5820) );
  AOI22D1BWP30P140LVT U16347 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[978]), .B1(n11751), .B2(
        inner_first_stage_data_reg[786]), .ZN(n11699) );
  AOI22D1BWP30P140LVT U16348 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1010]), .B1(n11750), .B2(
        inner_first_stage_data_reg[914]), .ZN(n11698) );
  AOI22D1BWP30P140LVT U16349 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[946]), .B1(n11752), .B2(
        inner_first_stage_data_reg[882]), .ZN(n11697) );
  AOI22D1BWP30P140LVT U16350 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[818]), .B1(n11754), .B2(
        inner_first_stage_data_reg[850]), .ZN(n11696) );
  ND4D1BWP30P140LVT U16351 ( .A1(n11699), .A2(n11698), .A3(n11697), .A4(n11696), .ZN(N5821) );
  AOI22D1BWP30P140LVT U16352 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1011]), .B1(n11751), .B2(
        inner_first_stage_data_reg[787]), .ZN(n11703) );
  AOI22D1BWP30P140LVT U16353 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[979]), .B1(n11750), .B2(
        inner_first_stage_data_reg[915]), .ZN(n11702) );
  AOI22D1BWP30P140LVT U16354 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[819]), .B1(n11754), .B2(
        inner_first_stage_data_reg[851]), .ZN(n11701) );
  AOI22D1BWP30P140LVT U16355 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[947]), .B1(n11752), .B2(
        inner_first_stage_data_reg[883]), .ZN(n11700) );
  ND4D1BWP30P140LVT U16356 ( .A1(n11703), .A2(n11702), .A3(n11701), .A4(n11700), .ZN(N5822) );
  AOI22D1BWP30P140LVT U16357 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[980]), .B1(n11751), .B2(
        inner_first_stage_data_reg[788]), .ZN(n11707) );
  AOI22D1BWP30P140LVT U16358 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1012]), .B1(n11750), .B2(
        inner_first_stage_data_reg[916]), .ZN(n11706) );
  AOI22D1BWP30P140LVT U16359 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[820]), .B1(n11754), .B2(
        inner_first_stage_data_reg[852]), .ZN(n11705) );
  AOI22D1BWP30P140LVT U16360 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[948]), .B1(n11752), .B2(
        inner_first_stage_data_reg[884]), .ZN(n11704) );
  ND4D1BWP30P140LVT U16361 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(N5823) );
  AOI22D1BWP30P140LVT U16362 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1013]), .B1(n11748), .B2(
        inner_first_stage_data_reg[981]), .ZN(n11711) );
  AOI22D1BWP30P140LVT U16363 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[789]), .B1(n11750), .B2(
        inner_first_stage_data_reg[917]), .ZN(n11710) );
  AOI22D1BWP30P140LVT U16364 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[949]), .B1(n11754), .B2(
        inner_first_stage_data_reg[853]), .ZN(n11709) );
  AOI22D1BWP30P140LVT U16365 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[821]), .B1(n11752), .B2(
        inner_first_stage_data_reg[885]), .ZN(n11708) );
  ND4D1BWP30P140LVT U16366 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(N5824) );
  AOI22D1BWP30P140LVT U16367 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1014]), .B1(n11751), .B2(
        inner_first_stage_data_reg[790]), .ZN(n11715) );
  AOI22D1BWP30P140LVT U16368 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[982]), .B1(n11750), .B2(
        inner_first_stage_data_reg[918]), .ZN(n11714) );
  AOI22D1BWP30P140LVT U16369 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[854]), .B1(n11752), .B2(
        inner_first_stage_data_reg[886]), .ZN(n11713) );
  AOI22D1BWP30P140LVT U16370 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[822]), .B1(n11753), .B2(
        inner_first_stage_data_reg[950]), .ZN(n11712) );
  ND4D1BWP30P140LVT U16371 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(N5825) );
  AOI22D1BWP30P140LVT U16372 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[983]), .B1(n11750), .B2(
        inner_first_stage_data_reg[919]), .ZN(n11719) );
  AOI22D1BWP30P140LVT U16373 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1015]), .B1(n11751), .B2(
        inner_first_stage_data_reg[791]), .ZN(n11718) );
  AOI22D1BWP30P140LVT U16374 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[951]), .B1(n11754), .B2(
        inner_first_stage_data_reg[855]), .ZN(n11717) );
  AOI22D1BWP30P140LVT U16375 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[823]), .B1(n11752), .B2(
        inner_first_stage_data_reg[887]), .ZN(n11716) );
  ND4D1BWP30P140LVT U16376 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(N5826) );
  AOI22D1BWP30P140LVT U16377 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1016]), .B1(n11748), .B2(
        inner_first_stage_data_reg[984]), .ZN(n11723) );
  AOI22D1BWP30P140LVT U16378 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[792]), .B1(n11750), .B2(
        inner_first_stage_data_reg[920]), .ZN(n11722) );
  AOI22D1BWP30P140LVT U16379 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[952]), .B1(n11752), .B2(
        inner_first_stage_data_reg[888]), .ZN(n11721) );
  AOI22D1BWP30P140LVT U16380 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[824]), .B1(n11754), .B2(
        inner_first_stage_data_reg[856]), .ZN(n11720) );
  ND4D1BWP30P140LVT U16381 ( .A1(n11723), .A2(n11722), .A3(n11721), .A4(n11720), .ZN(N5827) );
  AOI22D1BWP30P140LVT U16382 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1017]), .B1(n11750), .B2(
        inner_first_stage_data_reg[921]), .ZN(n11727) );
  AOI22D1BWP30P140LVT U16383 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[985]), .B1(n11751), .B2(
        inner_first_stage_data_reg[793]), .ZN(n11726) );
  AOI22D1BWP30P140LVT U16384 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[953]), .B1(n11752), .B2(
        inner_first_stage_data_reg[889]), .ZN(n11725) );
  AOI22D1BWP30P140LVT U16385 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[825]), .B1(n11754), .B2(
        inner_first_stage_data_reg[857]), .ZN(n11724) );
  ND4D1BWP30P140LVT U16386 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(N5828) );
  AOI22D1BWP30P140LVT U16387 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1018]), .B1(n11748), .B2(
        inner_first_stage_data_reg[986]), .ZN(n11731) );
  AOI22D1BWP30P140LVT U16388 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[794]), .B1(n11750), .B2(
        inner_first_stage_data_reg[922]), .ZN(n11730) );
  AOI22D1BWP30P140LVT U16389 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[826]), .B1(n11753), .B2(
        inner_first_stage_data_reg[954]), .ZN(n11729) );
  AOI22D1BWP30P140LVT U16390 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[858]), .B1(n11752), .B2(
        inner_first_stage_data_reg[890]), .ZN(n11728) );
  ND4D1BWP30P140LVT U16391 ( .A1(n11731), .A2(n11730), .A3(n11729), .A4(n11728), .ZN(N5829) );
  AOI22D1BWP30P140LVT U16392 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1019]), .B1(n11750), .B2(
        inner_first_stage_data_reg[923]), .ZN(n11735) );
  AOI22D1BWP30P140LVT U16393 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[987]), .B1(n11751), .B2(
        inner_first_stage_data_reg[795]), .ZN(n11734) );
  AOI22D1BWP30P140LVT U16394 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[955]), .B1(n11754), .B2(
        inner_first_stage_data_reg[859]), .ZN(n11733) );
  AOI22D1BWP30P140LVT U16395 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[827]), .B1(n11752), .B2(
        inner_first_stage_data_reg[891]), .ZN(n11732) );
  ND4D1BWP30P140LVT U16396 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(N5830) );
  AOI22D1BWP30P140LVT U16397 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[796]), .B1(n11750), .B2(
        inner_first_stage_data_reg[924]), .ZN(n11739) );
  AOI22D1BWP30P140LVT U16398 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1020]), .B1(n11748), .B2(
        inner_first_stage_data_reg[988]), .ZN(n11738) );
  AOI22D1BWP30P140LVT U16399 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[956]), .B1(n11752), .B2(
        inner_first_stage_data_reg[892]), .ZN(n11737) );
  AOI22D1BWP30P140LVT U16400 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[828]), .B1(n11754), .B2(
        inner_first_stage_data_reg[860]), .ZN(n11736) );
  ND4D1BWP30P140LVT U16401 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(N5831) );
  AOI22D1BWP30P140LVT U16402 ( .A1(n11748), .A2(
        inner_first_stage_data_reg[989]), .B1(n11751), .B2(
        inner_first_stage_data_reg[797]), .ZN(n11743) );
  AOI22D1BWP30P140LVT U16403 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1021]), .B1(n11750), .B2(
        inner_first_stage_data_reg[925]), .ZN(n11742) );
  AOI22D1BWP30P140LVT U16404 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[829]), .B1(n11754), .B2(
        inner_first_stage_data_reg[861]), .ZN(n11741) );
  AOI22D1BWP30P140LVT U16405 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[957]), .B1(n11752), .B2(
        inner_first_stage_data_reg[893]), .ZN(n11740) );
  ND4D1BWP30P140LVT U16406 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(N5832) );
  AOI22D1BWP30P140LVT U16407 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1022]), .B1(n11748), .B2(
        inner_first_stage_data_reg[990]), .ZN(n11747) );
  AOI22D1BWP30P140LVT U16408 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[798]), .B1(n11750), .B2(
        inner_first_stage_data_reg[926]), .ZN(n11746) );
  AOI22D1BWP30P140LVT U16409 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[830]), .B1(n11753), .B2(
        inner_first_stage_data_reg[958]), .ZN(n11745) );
  AOI22D1BWP30P140LVT U16410 ( .A1(n11754), .A2(
        inner_first_stage_data_reg[862]), .B1(n11752), .B2(
        inner_first_stage_data_reg[894]), .ZN(n11744) );
  ND4D1BWP30P140LVT U16411 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(N5833) );
  AOI22D1BWP30P140LVT U16412 ( .A1(n11749), .A2(
        inner_first_stage_data_reg[1023]), .B1(n11748), .B2(
        inner_first_stage_data_reg[991]), .ZN(n11759) );
  AOI22D1BWP30P140LVT U16413 ( .A1(n11751), .A2(
        inner_first_stage_data_reg[799]), .B1(n11750), .B2(
        inner_first_stage_data_reg[927]), .ZN(n11758) );
  AOI22D1BWP30P140LVT U16414 ( .A1(n11753), .A2(
        inner_first_stage_data_reg[959]), .B1(n11752), .B2(
        inner_first_stage_data_reg[895]), .ZN(n11757) );
  AOI22D1BWP30P140LVT U16415 ( .A1(n11755), .A2(
        inner_first_stage_data_reg[831]), .B1(n11754), .B2(
        inner_first_stage_data_reg[863]), .ZN(n11756) );
  ND4D1BWP30P140LVT U16416 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(N5834) );
  AOI22D1BWP30P140LVT U16417 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1088]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1152]), .ZN(n11763) );
  AOI22D1BWP30P140LVT U16418 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1120]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1024]), .ZN(n11762) );
  AOI22D1BWP30P140LVT U16419 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1216]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1248]), .ZN(n11761) );
  AOI22D1BWP30P140LVT U16420 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1184]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1056]), .ZN(n11760) );
  ND4D1BWP30P140LVT U16421 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(N7677) );
  AOI22D1BWP30P140LVT U16422 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1153]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1025]), .ZN(n11767) );
  AOI22D1BWP30P140LVT U16423 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1089]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1121]), .ZN(n11766) );
  AOI22D1BWP30P140LVT U16424 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1185]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1057]), .ZN(n11765) );
  AOI22D1BWP30P140LVT U16425 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1217]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1249]), .ZN(n11764) );
  ND4D1BWP30P140LVT U16426 ( .A1(n11767), .A2(n11766), .A3(n11765), .A4(n11764), .ZN(N7678) );
  AOI22D1BWP30P140LVT U16427 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1122]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1026]), .ZN(n11771) );
  AOI22D1BWP30P140LVT U16428 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1090]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1154]), .ZN(n11770) );
  AOI22D1BWP30P140LVT U16429 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1218]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1250]), .ZN(n11769) );
  AOI22D1BWP30P140LVT U16430 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1186]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1058]), .ZN(n11768) );
  ND4D1BWP30P140LVT U16431 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(N7679) );
  AOI22D1BWP30P140LVT U16432 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1155]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1027]), .ZN(n11775) );
  AOI22D1BWP30P140LVT U16433 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1091]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1123]), .ZN(n11774) );
  AOI22D1BWP30P140LVT U16434 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1219]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1059]), .ZN(n11773) );
  AOI22D1BWP30P140LVT U16435 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1251]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1187]), .ZN(n11772) );
  ND4D1BWP30P140LVT U16436 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(N7680) );
  AOI22D1BWP30P140LVT U16437 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1092]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1124]), .ZN(n11779) );
  AOI22D1BWP30P140LVT U16438 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1156]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1028]), .ZN(n11778) );
  AOI22D1BWP30P140LVT U16439 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1220]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1060]), .ZN(n11777) );
  AOI22D1BWP30P140LVT U16440 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1252]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1188]), .ZN(n11776) );
  ND4D1BWP30P140LVT U16441 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(N7681) );
  AOI22D1BWP30P140LVT U16442 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1093]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1125]), .ZN(n11783) );
  AOI22D1BWP30P140LVT U16443 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1157]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1029]), .ZN(n11782) );
  AOI22D1BWP30P140LVT U16444 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1221]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1189]), .ZN(n11781) );
  AOI22D1BWP30P140LVT U16445 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1253]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1061]), .ZN(n11780) );
  ND4D1BWP30P140LVT U16446 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(N7682) );
  AOI22D1BWP30P140LVT U16447 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1126]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1030]), .ZN(n11787) );
  AOI22D1BWP30P140LVT U16448 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1094]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1158]), .ZN(n11786) );
  AOI22D1BWP30P140LVT U16449 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1254]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1062]), .ZN(n11785) );
  AOI22D1BWP30P140LVT U16450 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1222]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1190]), .ZN(n11784) );
  ND4D1BWP30P140LVT U16451 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(N7683) );
  AOI22D1BWP30P140LVT U16452 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1095]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1159]), .ZN(n11791) );
  AOI22D1BWP30P140LVT U16453 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1127]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1031]), .ZN(n11790) );
  AOI22D1BWP30P140LVT U16454 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1223]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1255]), .ZN(n11789) );
  AOI22D1BWP30P140LVT U16455 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1191]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1063]), .ZN(n11788) );
  ND4D1BWP30P140LVT U16456 ( .A1(n11791), .A2(n11790), .A3(n11789), .A4(n11788), .ZN(N7684) );
  AOI22D1BWP30P140LVT U16457 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1160]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1032]), .ZN(n11795) );
  AOI22D1BWP30P140LVT U16458 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1096]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1128]), .ZN(n11794) );
  AOI22D1BWP30P140LVT U16459 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1192]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1064]), .ZN(n11793) );
  AOI22D1BWP30P140LVT U16460 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1224]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1256]), .ZN(n11792) );
  ND4D1BWP30P140LVT U16461 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(N7685) );
  AOI22D1BWP30P140LVT U16462 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1097]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1129]), .ZN(n11799) );
  AOI22D1BWP30P140LVT U16463 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1161]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1033]), .ZN(n11798) );
  AOI22D1BWP30P140LVT U16464 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1257]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1065]), .ZN(n11797) );
  AOI22D1BWP30P140LVT U16465 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1225]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1193]), .ZN(n11796) );
  ND4D1BWP30P140LVT U16466 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(N7686) );
  AOI22D1BWP30P140LVT U16467 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1098]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1130]), .ZN(n11803) );
  AOI22D1BWP30P140LVT U16468 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1162]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1034]), .ZN(n11802) );
  AOI22D1BWP30P140LVT U16469 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1258]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1066]), .ZN(n11801) );
  AOI22D1BWP30P140LVT U16470 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1226]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1194]), .ZN(n11800) );
  ND4D1BWP30P140LVT U16471 ( .A1(n11803), .A2(n11802), .A3(n11801), .A4(n11800), .ZN(N7687) );
  AOI22D1BWP30P140LVT U16472 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1131]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1035]), .ZN(n11807) );
  AOI22D1BWP30P140LVT U16473 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1099]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1163]), .ZN(n11806) );
  AOI22D1BWP30P140LVT U16474 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1259]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1067]), .ZN(n11805) );
  AOI22D1BWP30P140LVT U16475 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1227]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1195]), .ZN(n11804) );
  ND4D1BWP30P140LVT U16476 ( .A1(n11807), .A2(n11806), .A3(n11805), .A4(n11804), .ZN(N7688) );
  AOI22D1BWP30P140LVT U16477 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1164]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1132]), .ZN(n11811) );
  AOI22D1BWP30P140LVT U16478 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1100]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1036]), .ZN(n11810) );
  AOI22D1BWP30P140LVT U16479 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1228]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1196]), .ZN(n11809) );
  AOI22D1BWP30P140LVT U16480 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1260]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1068]), .ZN(n11808) );
  ND4D1BWP30P140LVT U16481 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(N7689) );
  AOI22D1BWP30P140LVT U16482 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1101]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1133]), .ZN(n11815) );
  AOI22D1BWP30P140LVT U16483 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1165]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1037]), .ZN(n11814) );
  AOI22D1BWP30P140LVT U16484 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1229]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1069]), .ZN(n11813) );
  AOI22D1BWP30P140LVT U16485 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1261]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1197]), .ZN(n11812) );
  ND4D1BWP30P140LVT U16486 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(N7690) );
  AOI22D1BWP30P140LVT U16487 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1102]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1134]), .ZN(n11819) );
  AOI22D1BWP30P140LVT U16488 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1166]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1038]), .ZN(n11818) );
  AOI22D1BWP30P140LVT U16489 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1230]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1070]), .ZN(n11817) );
  AOI22D1BWP30P140LVT U16490 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1262]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1198]), .ZN(n11816) );
  ND4D1BWP30P140LVT U16491 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(N7691) );
  AOI22D1BWP30P140LVT U16492 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1167]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1135]), .ZN(n11823) );
  AOI22D1BWP30P140LVT U16493 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1103]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1039]), .ZN(n11822) );
  AOI22D1BWP30P140LVT U16494 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1199]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1071]), .ZN(n11821) );
  AOI22D1BWP30P140LVT U16495 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1231]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1263]), .ZN(n11820) );
  ND4D1BWP30P140LVT U16496 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(N7692) );
  AOI22D1BWP30P140LVT U16497 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1168]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1136]), .ZN(n11827) );
  AOI22D1BWP30P140LVT U16498 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1104]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1040]), .ZN(n11826) );
  AOI22D1BWP30P140LVT U16499 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1232]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1072]), .ZN(n11825) );
  AOI22D1BWP30P140LVT U16500 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1264]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1200]), .ZN(n11824) );
  ND4D1BWP30P140LVT U16501 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(N7693) );
  AOI22D1BWP30P140LVT U16502 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1169]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1137]), .ZN(n11831) );
  AOI22D1BWP30P140LVT U16503 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1105]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1041]), .ZN(n11830) );
  AOI22D1BWP30P140LVT U16504 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1201]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1073]), .ZN(n11829) );
  AOI22D1BWP30P140LVT U16505 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1233]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1265]), .ZN(n11828) );
  ND4D1BWP30P140LVT U16506 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(N7694) );
  AOI22D1BWP30P140LVT U16507 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1170]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1042]), .ZN(n11835) );
  AOI22D1BWP30P140LVT U16508 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1106]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1138]), .ZN(n11834) );
  AOI22D1BWP30P140LVT U16509 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1234]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1266]), .ZN(n11833) );
  AOI22D1BWP30P140LVT U16510 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1202]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1074]), .ZN(n11832) );
  ND4D1BWP30P140LVT U16511 ( .A1(n11835), .A2(n11834), .A3(n11833), .A4(n11832), .ZN(N7695) );
  AOI22D1BWP30P140LVT U16512 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1107]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1171]), .ZN(n11839) );
  AOI22D1BWP30P140LVT U16513 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1139]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1043]), .ZN(n11838) );
  AOI22D1BWP30P140LVT U16514 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1235]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1267]), .ZN(n11837) );
  AOI22D1BWP30P140LVT U16515 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1203]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1075]), .ZN(n11836) );
  ND4D1BWP30P140LVT U16516 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(N7696) );
  AOI22D1BWP30P140LVT U16517 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1108]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1044]), .ZN(n11843) );
  AOI22D1BWP30P140LVT U16518 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1172]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1140]), .ZN(n11842) );
  AOI22D1BWP30P140LVT U16519 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1268]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1076]), .ZN(n11841) );
  AOI22D1BWP30P140LVT U16520 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1236]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1204]), .ZN(n11840) );
  ND4D1BWP30P140LVT U16521 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(N7697) );
  AOI22D1BWP30P140LVT U16522 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1109]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1141]), .ZN(n11847) );
  AOI22D1BWP30P140LVT U16523 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1173]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1045]), .ZN(n11846) );
  AOI22D1BWP30P140LVT U16524 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1205]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1077]), .ZN(n11845) );
  AOI22D1BWP30P140LVT U16525 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1237]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1269]), .ZN(n11844) );
  ND4D1BWP30P140LVT U16526 ( .A1(n11847), .A2(n11846), .A3(n11845), .A4(n11844), .ZN(N7698) );
  AOI22D1BWP30P140LVT U16527 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1142]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1046]), .ZN(n11851) );
  AOI22D1BWP30P140LVT U16528 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1110]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1174]), .ZN(n11850) );
  AOI22D1BWP30P140LVT U16529 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1238]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1078]), .ZN(n11849) );
  AOI22D1BWP30P140LVT U16530 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1270]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1206]), .ZN(n11848) );
  ND4D1BWP30P140LVT U16531 ( .A1(n11851), .A2(n11850), .A3(n11849), .A4(n11848), .ZN(N7699) );
  AOI22D1BWP30P140LVT U16532 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1111]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1175]), .ZN(n11855) );
  AOI22D1BWP30P140LVT U16533 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1143]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1047]), .ZN(n11854) );
  AOI22D1BWP30P140LVT U16534 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1271]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1207]), .ZN(n11853) );
  AOI22D1BWP30P140LVT U16535 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1239]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1079]), .ZN(n11852) );
  ND4D1BWP30P140LVT U16536 ( .A1(n11855), .A2(n11854), .A3(n11853), .A4(n11852), .ZN(N7700) );
  AOI22D1BWP30P140LVT U16537 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1144]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1048]), .ZN(n11859) );
  AOI22D1BWP30P140LVT U16538 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1112]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1176]), .ZN(n11858) );
  AOI22D1BWP30P140LVT U16539 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1272]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1208]), .ZN(n11857) );
  AOI22D1BWP30P140LVT U16540 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1240]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1080]), .ZN(n11856) );
  ND4D1BWP30P140LVT U16541 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(N7701) );
  AOI22D1BWP30P140LVT U16542 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1113]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1177]), .ZN(n11863) );
  AOI22D1BWP30P140LVT U16543 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1145]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1049]), .ZN(n11862) );
  AOI22D1BWP30P140LVT U16544 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1273]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1209]), .ZN(n11861) );
  AOI22D1BWP30P140LVT U16545 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1241]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1081]), .ZN(n11860) );
  ND4D1BWP30P140LVT U16546 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(N7702) );
  AOI22D1BWP30P140LVT U16547 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1146]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1050]), .ZN(n11867) );
  AOI22D1BWP30P140LVT U16548 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1114]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1178]), .ZN(n11866) );
  AOI22D1BWP30P140LVT U16549 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1242]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1082]), .ZN(n11865) );
  AOI22D1BWP30P140LVT U16550 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1274]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1210]), .ZN(n11864) );
  ND4D1BWP30P140LVT U16551 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(N7703) );
  AOI22D1BWP30P140LVT U16552 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1115]), .B1(n11887), .B2(
        inner_first_stage_data_reg[1179]), .ZN(n11871) );
  AOI22D1BWP30P140LVT U16553 ( .A1(n11884), .A2(
        inner_first_stage_data_reg[1147]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1051]), .ZN(n11870) );
  AOI22D1BWP30P140LVT U16554 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1243]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1275]), .ZN(n11869) );
  AOI22D1BWP30P140LVT U16555 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1211]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1083]), .ZN(n11868) );
  ND4D1BWP30P140LVT U16556 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(N7704) );
  AOI22D1BWP30P140LVT U16557 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1116]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1148]), .ZN(n11875) );
  AOI22D1BWP30P140LVT U16558 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1180]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1052]), .ZN(n11874) );
  AOI22D1BWP30P140LVT U16559 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1212]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1084]), .ZN(n11873) );
  AOI22D1BWP30P140LVT U16560 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1244]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1276]), .ZN(n11872) );
  ND4D1BWP30P140LVT U16561 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(N7705) );
  AOI22D1BWP30P140LVT U16562 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1117]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1053]), .ZN(n11879) );
  AOI22D1BWP30P140LVT U16563 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1181]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1149]), .ZN(n11878) );
  AOI22D1BWP30P140LVT U16564 ( .A1(n11888), .A2(
        inner_first_stage_data_reg[1277]), .B1(n11891), .B2(
        inner_first_stage_data_reg[1213]), .ZN(n11877) );
  AOI22D1BWP30P140LVT U16565 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1245]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1085]), .ZN(n11876) );
  ND4D1BWP30P140LVT U16566 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(N7706) );
  AOI22D1BWP30P140LVT U16567 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1182]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1150]), .ZN(n11883) );
  AOI22D1BWP30P140LVT U16568 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1118]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1054]), .ZN(n11882) );
  AOI22D1BWP30P140LVT U16569 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1246]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1278]), .ZN(n11881) );
  AOI22D1BWP30P140LVT U16570 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1214]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1086]), .ZN(n11880) );
  ND4D1BWP30P140LVT U16571 ( .A1(n11883), .A2(n11882), .A3(n11881), .A4(n11880), .ZN(N7707) );
  AOI22D1BWP30P140LVT U16572 ( .A1(n11885), .A2(
        inner_first_stage_data_reg[1119]), .B1(n11884), .B2(
        inner_first_stage_data_reg[1151]), .ZN(n11895) );
  AOI22D1BWP30P140LVT U16573 ( .A1(n11887), .A2(
        inner_first_stage_data_reg[1183]), .B1(n11886), .B2(
        inner_first_stage_data_reg[1055]), .ZN(n11894) );
  AOI22D1BWP30P140LVT U16574 ( .A1(n11889), .A2(
        inner_first_stage_data_reg[1247]), .B1(n11888), .B2(
        inner_first_stage_data_reg[1279]), .ZN(n11893) );
  AOI22D1BWP30P140LVT U16575 ( .A1(n11891), .A2(
        inner_first_stage_data_reg[1215]), .B1(n11890), .B2(
        inner_first_stage_data_reg[1087]), .ZN(n11892) );
  ND4D1BWP30P140LVT U16576 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(N7708) );
  AOI22D1BWP30P140LVT U16577 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1408]), .B1(n12025), .B2(
        inner_first_stage_data_reg[1376]), .ZN(n11899) );
  AOI22D1BWP30P140LVT U16578 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1312]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1440]), .ZN(n11898) );
  AOI22D1BWP30P140LVT U16579 ( .A1(n12024), .A2(
        inner_first_stage_data_reg[1344]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1280]), .ZN(n11897) );
  AOI22D1BWP30P140LVT U16580 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1504]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1472]), .ZN(n11896) );
  ND4D1BWP30P140LVT U16581 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(N8527) );
  AOI22D1BWP30P140LVT U16582 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1377]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1345]), .ZN(n11903) );
  AOI22D1BWP30P140LVT U16583 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1409]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1281]), .ZN(n11902) );
  AOI22D1BWP30P140LVT U16584 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1313]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1441]), .ZN(n11901) );
  AOI22D1BWP30P140LVT U16585 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1505]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1473]), .ZN(n11900) );
  ND4D1BWP30P140LVT U16586 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(N8528) );
  AOI22D1BWP30P140LVT U16587 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1314]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1282]), .ZN(n11907) );
  AOI22D1BWP30P140LVT U16588 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1410]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1442]), .ZN(n11906) );
  AOI22D1BWP30P140LVT U16589 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1378]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1346]), .ZN(n11905) );
  AOI22D1BWP30P140LVT U16590 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1506]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1474]), .ZN(n11904) );
  ND4D1BWP30P140LVT U16591 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(N8529) );
  AOI22D1BWP30P140LVT U16592 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1411]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1315]), .ZN(n11911) );
  AOI22D1BWP30P140LVT U16593 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1379]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1347]), .ZN(n11910) );
  AOI22D1BWP30P140LVT U16594 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1443]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1283]), .ZN(n11909) );
  AOI22D1BWP30P140LVT U16595 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1507]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1475]), .ZN(n11908) );
  ND4D1BWP30P140LVT U16596 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(N8530) );
  AOI22D1BWP30P140LVT U16597 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1412]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1284]), .ZN(n11915) );
  AOI22D1BWP30P140LVT U16598 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1316]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1348]), .ZN(n11914) );
  AOI22D1BWP30P140LVT U16599 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1380]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1444]), .ZN(n11913) );
  AOI22D1BWP30P140LVT U16600 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1508]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1476]), .ZN(n11912) );
  ND4D1BWP30P140LVT U16601 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(N8531) );
  AOI22D1BWP30P140LVT U16602 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1381]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1445]), .ZN(n11919) );
  AOI22D1BWP30P140LVT U16603 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1317]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1349]), .ZN(n11918) );
  AOI22D1BWP30P140LVT U16604 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1413]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1285]), .ZN(n11917) );
  AOI22D1BWP30P140LVT U16605 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1509]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1477]), .ZN(n11916) );
  ND4D1BWP30P140LVT U16606 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(N8532) );
  AOI22D1BWP30P140LVT U16607 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1382]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1286]), .ZN(n11923) );
  AOI22D1BWP30P140LVT U16608 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1414]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1350]), .ZN(n11922) );
  AOI22D1BWP30P140LVT U16609 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1318]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1446]), .ZN(n11921) );
  AOI22D1BWP30P140LVT U16610 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1510]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1478]), .ZN(n11920) );
  ND4D1BWP30P140LVT U16611 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(N8533) );
  AOI22D1BWP30P140LVT U16612 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1383]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1287]), .ZN(n11927) );
  AOI22D1BWP30P140LVT U16613 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1319]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1447]), .ZN(n11926) );
  AOI22D1BWP30P140LVT U16614 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1415]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1351]), .ZN(n11925) );
  AOI22D1BWP30P140LVT U16615 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1511]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1479]), .ZN(n11924) );
  ND4D1BWP30P140LVT U16616 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(N8534) );
  AOI22D1BWP30P140LVT U16617 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1320]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1448]), .ZN(n11931) );
  AOI22D1BWP30P140LVT U16618 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1416]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1288]), .ZN(n11930) );
  AOI22D1BWP30P140LVT U16619 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1384]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1352]), .ZN(n11929) );
  AOI22D1BWP30P140LVT U16620 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1512]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1480]), .ZN(n11928) );
  ND4D1BWP30P140LVT U16621 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(N8535) );
  AOI22D1BWP30P140LVT U16622 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1321]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1289]), .ZN(n11935) );
  AOI22D1BWP30P140LVT U16623 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1417]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1449]), .ZN(n11934) );
  AOI22D1BWP30P140LVT U16624 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1385]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1353]), .ZN(n11933) );
  AOI22D1BWP30P140LVT U16625 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1513]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1481]), .ZN(n11932) );
  ND4D1BWP30P140LVT U16626 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(N8536) );
  AOI22D1BWP30P140LVT U16627 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1450]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1290]), .ZN(n11939) );
  AOI22D1BWP30P140LVT U16628 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1418]), .B1(n12025), .B2(
        inner_first_stage_data_reg[1386]), .ZN(n11938) );
  AOI22D1BWP30P140LVT U16629 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1322]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1354]), .ZN(n11937) );
  AOI22D1BWP30P140LVT U16630 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1514]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1482]), .ZN(n11936) );
  ND4D1BWP30P140LVT U16631 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(N8537) );
  AOI22D1BWP30P140LVT U16632 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1387]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1323]), .ZN(n11943) );
  AOI22D1BWP30P140LVT U16633 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1451]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1291]), .ZN(n11942) );
  AOI22D1BWP30P140LVT U16634 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1419]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1355]), .ZN(n11941) );
  AOI22D1BWP30P140LVT U16635 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1515]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1483]), .ZN(n11940) );
  ND4D1BWP30P140LVT U16636 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(N8538) );
  AOI22D1BWP30P140LVT U16637 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1452]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1292]), .ZN(n11947) );
  AOI22D1BWP30P140LVT U16638 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1388]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1324]), .ZN(n11946) );
  AOI22D1BWP30P140LVT U16639 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1420]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1356]), .ZN(n11945) );
  AOI22D1BWP30P140LVT U16640 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1516]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1484]), .ZN(n11944) );
  ND4D1BWP30P140LVT U16641 ( .A1(n11947), .A2(n11946), .A3(n11945), .A4(n11944), .ZN(N8539) );
  AOI22D1BWP30P140LVT U16642 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1325]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1357]), .ZN(n11951) );
  AOI22D1BWP30P140LVT U16643 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1421]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1453]), .ZN(n11950) );
  AOI22D1BWP30P140LVT U16644 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1389]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1293]), .ZN(n11949) );
  AOI22D1BWP30P140LVT U16645 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1517]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1485]), .ZN(n11948) );
  ND4D1BWP30P140LVT U16646 ( .A1(n11951), .A2(n11950), .A3(n11949), .A4(n11948), .ZN(N8540) );
  AOI22D1BWP30P140LVT U16647 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1390]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1358]), .ZN(n11955) );
  AOI22D1BWP30P140LVT U16648 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1422]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1454]), .ZN(n11954) );
  AOI22D1BWP30P140LVT U16649 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1326]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1294]), .ZN(n11953) );
  AOI22D1BWP30P140LVT U16650 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1518]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1486]), .ZN(n11952) );
  ND4D1BWP30P140LVT U16651 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(N8541) );
  AOI22D1BWP30P140LVT U16652 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1391]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1455]), .ZN(n11959) );
  AOI22D1BWP30P140LVT U16653 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1423]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1295]), .ZN(n11958) );
  AOI22D1BWP30P140LVT U16654 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1327]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1359]), .ZN(n11957) );
  AOI22D1BWP30P140LVT U16655 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1519]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1487]), .ZN(n11956) );
  ND4D1BWP30P140LVT U16656 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(N8542) );
  AOI22D1BWP30P140LVT U16657 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1392]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1296]), .ZN(n11963) );
  AOI22D1BWP30P140LVT U16658 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1328]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1456]), .ZN(n11962) );
  AOI22D1BWP30P140LVT U16659 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1424]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1360]), .ZN(n11961) );
  AOI22D1BWP30P140LVT U16660 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1520]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1488]), .ZN(n11960) );
  ND4D1BWP30P140LVT U16661 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(N8543) );
  AOI22D1BWP30P140LVT U16662 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1393]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1457]), .ZN(n11967) );
  AOI22D1BWP30P140LVT U16663 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1329]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1297]), .ZN(n11966) );
  AOI22D1BWP30P140LVT U16664 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1425]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1361]), .ZN(n11965) );
  AOI22D1BWP30P140LVT U16665 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1521]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1489]), .ZN(n11964) );
  ND4D1BWP30P140LVT U16666 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(N8544) );
  AOI22D1BWP30P140LVT U16667 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1426]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1298]), .ZN(n11971) );
  AOI22D1BWP30P140LVT U16668 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1394]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1330]), .ZN(n11970) );
  AOI22D1BWP30P140LVT U16669 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1458]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1362]), .ZN(n11969) );
  AOI22D1BWP30P140LVT U16670 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1522]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1490]), .ZN(n11968) );
  ND4D1BWP30P140LVT U16671 ( .A1(n11971), .A2(n11970), .A3(n11969), .A4(n11968), .ZN(N8545) );
  AOI22D1BWP30P140LVT U16672 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1395]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1299]), .ZN(n11975) );
  AOI22D1BWP30P140LVT U16673 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1427]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1331]), .ZN(n11974) );
  AOI22D1BWP30P140LVT U16674 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1459]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1363]), .ZN(n11973) );
  AOI22D1BWP30P140LVT U16675 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1523]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1491]), .ZN(n11972) );
  ND4D1BWP30P140LVT U16676 ( .A1(n11975), .A2(n11974), .A3(n11973), .A4(n11972), .ZN(N8546) );
  AOI22D1BWP30P140LVT U16677 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1428]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1300]), .ZN(n11979) );
  AOI22D1BWP30P140LVT U16678 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1396]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1332]), .ZN(n11978) );
  AOI22D1BWP30P140LVT U16679 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1460]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1364]), .ZN(n11977) );
  AOI22D1BWP30P140LVT U16680 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1524]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1492]), .ZN(n11976) );
  ND4D1BWP30P140LVT U16681 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(N8547) );
  AOI22D1BWP30P140LVT U16682 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1461]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1301]), .ZN(n11983) );
  AOI22D1BWP30P140LVT U16683 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1397]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1365]), .ZN(n11982) );
  AOI22D1BWP30P140LVT U16684 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1429]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1333]), .ZN(n11981) );
  AOI22D1BWP30P140LVT U16685 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1525]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1493]), .ZN(n11980) );
  ND4D1BWP30P140LVT U16686 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(N8548) );
  AOI22D1BWP30P140LVT U16687 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1398]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1462]), .ZN(n11987) );
  AOI22D1BWP30P140LVT U16688 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1334]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1302]), .ZN(n11986) );
  AOI22D1BWP30P140LVT U16689 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1430]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1366]), .ZN(n11985) );
  AOI22D1BWP30P140LVT U16690 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1526]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1494]), .ZN(n11984) );
  ND4D1BWP30P140LVT U16691 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(N8549) );
  AOI22D1BWP30P140LVT U16692 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1335]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1367]), .ZN(n11991) );
  AOI22D1BWP30P140LVT U16693 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1399]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1303]), .ZN(n11990) );
  AOI22D1BWP30P140LVT U16694 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1431]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1463]), .ZN(n11989) );
  AOI22D1BWP30P140LVT U16695 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1527]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1495]), .ZN(n11988) );
  ND4D1BWP30P140LVT U16696 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(N8550) );
  AOI22D1BWP30P140LVT U16697 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1400]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1336]), .ZN(n11995) );
  AOI22D1BWP30P140LVT U16698 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1432]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1464]), .ZN(n11994) );
  AOI22D1BWP30P140LVT U16699 ( .A1(n12024), .A2(
        inner_first_stage_data_reg[1368]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1304]), .ZN(n11993) );
  AOI22D1BWP30P140LVT U16700 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1528]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1496]), .ZN(n11992) );
  ND4D1BWP30P140LVT U16701 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(N8551) );
  AOI22D1BWP30P140LVT U16702 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1465]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1305]), .ZN(n11999) );
  AOI22D1BWP30P140LVT U16703 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1433]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1369]), .ZN(n11998) );
  AOI22D1BWP30P140LVT U16704 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1401]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1337]), .ZN(n11997) );
  AOI22D1BWP30P140LVT U16705 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1529]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1497]), .ZN(n11996) );
  ND4D1BWP30P140LVT U16706 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(N8552) );
  AOI22D1BWP30P140LVT U16707 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1402]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1306]), .ZN(n12003) );
  AOI22D1BWP30P140LVT U16708 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1338]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1370]), .ZN(n12002) );
  AOI22D1BWP30P140LVT U16709 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1434]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1466]), .ZN(n12001) );
  AOI22D1BWP30P140LVT U16710 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1530]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1498]), .ZN(n12000) );
  ND4D1BWP30P140LVT U16711 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(N8553) );
  AOI22D1BWP30P140LVT U16712 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1435]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1467]), .ZN(n12007) );
  AOI22D1BWP30P140LVT U16713 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1403]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1307]), .ZN(n12006) );
  AOI22D1BWP30P140LVT U16714 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1339]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1371]), .ZN(n12005) );
  AOI22D1BWP30P140LVT U16715 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1531]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1499]), .ZN(n12004) );
  ND4D1BWP30P140LVT U16716 ( .A1(n12007), .A2(n12006), .A3(n12005), .A4(n12004), .ZN(N8554) );
  AOI22D1BWP30P140LVT U16717 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1404]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1308]), .ZN(n12011) );
  AOI22D1BWP30P140LVT U16718 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1436]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1468]), .ZN(n12010) );
  AOI22D1BWP30P140LVT U16719 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1340]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1372]), .ZN(n12009) );
  AOI22D1BWP30P140LVT U16720 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1532]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1500]), .ZN(n12008) );
  ND4D1BWP30P140LVT U16721 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(N8555) );
  AOI22D1BWP30P140LVT U16722 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1437]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1469]), .ZN(n12015) );
  AOI22D1BWP30P140LVT U16723 ( .A1(n12024), .A2(
        inner_first_stage_data_reg[1373]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1309]), .ZN(n12014) );
  AOI22D1BWP30P140LVT U16724 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1405]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1341]), .ZN(n12013) );
  AOI22D1BWP30P140LVT U16725 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1533]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1501]), .ZN(n12012) );
  ND4D1BWP30P140LVT U16726 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(N8556) );
  AOI22D1BWP30P140LVT U16727 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1406]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1374]), .ZN(n12019) );
  AOI22D1BWP30P140LVT U16728 ( .A1(n12020), .A2(
        inner_first_stage_data_reg[1470]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1310]), .ZN(n12018) );
  AOI22D1BWP30P140LVT U16729 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1438]), .B1(n12023), .B2(
        inner_first_stage_data_reg[1342]), .ZN(n12017) );
  AOI22D1BWP30P140LVT U16730 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1534]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1502]), .ZN(n12016) );
  ND4D1BWP30P140LVT U16731 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(N8557) );
  AOI22D1BWP30P140LVT U16732 ( .A1(n12021), .A2(
        inner_first_stage_data_reg[1439]), .B1(n12020), .B2(
        inner_first_stage_data_reg[1471]), .ZN(n12031) );
  AOI22D1BWP30P140LVT U16733 ( .A1(n12023), .A2(
        inner_first_stage_data_reg[1343]), .B1(n12022), .B2(
        inner_first_stage_data_reg[1311]), .ZN(n12030) );
  AOI22D1BWP30P140LVT U16734 ( .A1(n12025), .A2(
        inner_first_stage_data_reg[1407]), .B1(n12024), .B2(
        inner_first_stage_data_reg[1375]), .ZN(n12029) );
  AOI22D1BWP30P140LVT U16735 ( .A1(n12027), .A2(
        inner_first_stage_data_reg[1535]), .B1(n12026), .B2(
        inner_first_stage_data_reg[1503]), .ZN(n12028) );
  ND4D1BWP30P140LVT U16736 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(N8558) );
  AOI22D1BWP30P140LVT U16737 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1664]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1536]), .ZN(n12035) );
  AOI22D1BWP30P140LVT U16738 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1728]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1760]), .ZN(n12034) );
  AOI22D1BWP30P140LVT U16739 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1568]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1632]), .ZN(n12033) );
  AOI22D1BWP30P140LVT U16740 ( .A1(n12161), .A2(
        inner_first_stage_data_reg[1696]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1600]), .ZN(n12032) );
  ND4D1BWP30P140LVT U16741 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(N10401) );
  AOI22D1BWP30P140LVT U16742 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1665]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1537]), .ZN(n12039) );
  AOI22D1BWP30P140LVT U16743 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1633]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1601]), .ZN(n12038) );
  AOI22D1BWP30P140LVT U16744 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1729]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1569]), .ZN(n12037) );
  AOI22D1BWP30P140LVT U16745 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1761]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1697]), .ZN(n12036) );
  ND4D1BWP30P140LVT U16746 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(N10402) );
  AOI22D1BWP30P140LVT U16747 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1666]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1538]), .ZN(n12043) );
  AOI22D1BWP30P140LVT U16748 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1762]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1634]), .ZN(n12042) );
  AOI22D1BWP30P140LVT U16749 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1730]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1602]), .ZN(n12041) );
  AOI22D1BWP30P140LVT U16750 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1570]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1698]), .ZN(n12040) );
  ND4D1BWP30P140LVT U16751 ( .A1(n12043), .A2(n12042), .A3(n12041), .A4(n12040), .ZN(N10403) );
  AOI22D1BWP30P140LVT U16752 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1667]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1539]), .ZN(n12047) );
  AOI22D1BWP30P140LVT U16753 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1731]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1571]), .ZN(n12046) );
  AOI22D1BWP30P140LVT U16754 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1763]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1635]), .ZN(n12045) );
  AOI22D1BWP30P140LVT U16755 ( .A1(n12161), .A2(
        inner_first_stage_data_reg[1699]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1603]), .ZN(n12044) );
  ND4D1BWP30P140LVT U16756 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(N10404) );
  AOI22D1BWP30P140LVT U16757 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1668]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1540]), .ZN(n12051) );
  AOI22D1BWP30P140LVT U16758 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1764]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1636]), .ZN(n12050) );
  AOI22D1BWP30P140LVT U16759 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1732]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1604]), .ZN(n12049) );
  AOI22D1BWP30P140LVT U16760 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1572]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1700]), .ZN(n12048) );
  ND4D1BWP30P140LVT U16761 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(N10405) );
  AOI22D1BWP30P140LVT U16762 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1669]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1541]), .ZN(n12055) );
  AOI22D1BWP30P140LVT U16763 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1573]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1605]), .ZN(n12054) );
  AOI22D1BWP30P140LVT U16764 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1733]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1765]), .ZN(n12053) );
  AOI22D1BWP30P140LVT U16765 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1637]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1701]), .ZN(n12052) );
  ND4D1BWP30P140LVT U16766 ( .A1(n12055), .A2(n12054), .A3(n12053), .A4(n12052), .ZN(N10406) );
  AOI22D1BWP30P140LVT U16767 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1670]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1542]), .ZN(n12059) );
  AOI22D1BWP30P140LVT U16768 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1734]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1702]), .ZN(n12058) );
  AOI22D1BWP30P140LVT U16769 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1766]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1574]), .ZN(n12057) );
  AOI22D1BWP30P140LVT U16770 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1638]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1606]), .ZN(n12056) );
  ND4D1BWP30P140LVT U16771 ( .A1(n12059), .A2(n12058), .A3(n12057), .A4(n12056), .ZN(N10407) );
  AOI22D1BWP30P140LVT U16772 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1671]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1543]), .ZN(n12063) );
  AOI22D1BWP30P140LVT U16773 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1735]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1767]), .ZN(n12062) );
  AOI22D1BWP30P140LVT U16774 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1639]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1607]), .ZN(n12061) );
  AOI22D1BWP30P140LVT U16775 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1575]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1703]), .ZN(n12060) );
  ND4D1BWP30P140LVT U16776 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(N10408) );
  AOI22D1BWP30P140LVT U16777 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1672]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1544]), .ZN(n12067) );
  AOI22D1BWP30P140LVT U16778 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1640]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1608]), .ZN(n12066) );
  AOI22D1BWP30P140LVT U16779 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1576]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1704]), .ZN(n12065) );
  AOI22D1BWP30P140LVT U16780 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1736]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1768]), .ZN(n12064) );
  ND4D1BWP30P140LVT U16781 ( .A1(n12067), .A2(n12066), .A3(n12065), .A4(n12064), .ZN(N10409) );
  AOI22D1BWP30P140LVT U16782 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1673]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1545]), .ZN(n12071) );
  AOI22D1BWP30P140LVT U16783 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1737]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1705]), .ZN(n12070) );
  AOI22D1BWP30P140LVT U16784 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1769]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1577]), .ZN(n12069) );
  AOI22D1BWP30P140LVT U16785 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1641]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1609]), .ZN(n12068) );
  ND4D1BWP30P140LVT U16786 ( .A1(n12071), .A2(n12070), .A3(n12069), .A4(n12068), .ZN(N10410) );
  AOI22D1BWP30P140LVT U16787 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1674]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1546]), .ZN(n12075) );
  AOI22D1BWP30P140LVT U16788 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1738]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1706]), .ZN(n12074) );
  AOI22D1BWP30P140LVT U16789 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1770]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1642]), .ZN(n12073) );
  AOI22D1BWP30P140LVT U16790 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1578]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1610]), .ZN(n12072) );
  ND4D1BWP30P140LVT U16791 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(N10411) );
  AOI22D1BWP30P140LVT U16792 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1675]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1547]), .ZN(n12079) );
  AOI22D1BWP30P140LVT U16793 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1579]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1707]), .ZN(n12078) );
  AOI22D1BWP30P140LVT U16794 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1643]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1611]), .ZN(n12077) );
  AOI22D1BWP30P140LVT U16795 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1739]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1771]), .ZN(n12076) );
  ND4D1BWP30P140LVT U16796 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(N10412) );
  AOI22D1BWP30P140LVT U16797 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1676]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1548]), .ZN(n12083) );
  AOI22D1BWP30P140LVT U16798 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1740]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1708]), .ZN(n12082) );
  AOI22D1BWP30P140LVT U16799 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1772]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1612]), .ZN(n12081) );
  AOI22D1BWP30P140LVT U16800 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1580]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1644]), .ZN(n12080) );
  ND4D1BWP30P140LVT U16801 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(N10413) );
  AOI22D1BWP30P140LVT U16802 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1677]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1549]), .ZN(n12087) );
  AOI22D1BWP30P140LVT U16803 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1773]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1581]), .ZN(n12086) );
  AOI22D1BWP30P140LVT U16804 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1645]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1613]), .ZN(n12085) );
  AOI22D1BWP30P140LVT U16805 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1741]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1709]), .ZN(n12084) );
  ND4D1BWP30P140LVT U16806 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(N10414) );
  AOI22D1BWP30P140LVT U16807 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1678]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1550]), .ZN(n12091) );
  AOI22D1BWP30P140LVT U16808 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1774]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1614]), .ZN(n12090) );
  AOI22D1BWP30P140LVT U16809 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1742]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1710]), .ZN(n12089) );
  AOI22D1BWP30P140LVT U16810 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1582]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1646]), .ZN(n12088) );
  ND4D1BWP30P140LVT U16811 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(N10415) );
  AOI22D1BWP30P140LVT U16812 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1679]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1551]), .ZN(n12095) );
  AOI22D1BWP30P140LVT U16813 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1583]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1615]), .ZN(n12094) );
  AOI22D1BWP30P140LVT U16814 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1775]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1647]), .ZN(n12093) );
  AOI22D1BWP30P140LVT U16815 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1743]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1711]), .ZN(n12092) );
  ND4D1BWP30P140LVT U16816 ( .A1(n12095), .A2(n12094), .A3(n12093), .A4(n12092), .ZN(N10416) );
  AOI22D1BWP30P140LVT U16817 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1680]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1552]), .ZN(n12099) );
  AOI22D1BWP30P140LVT U16818 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1744]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1648]), .ZN(n12098) );
  AOI22D1BWP30P140LVT U16819 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1584]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1712]), .ZN(n12097) );
  AOI22D1BWP30P140LVT U16820 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1776]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1616]), .ZN(n12096) );
  ND4D1BWP30P140LVT U16821 ( .A1(n12099), .A2(n12098), .A3(n12097), .A4(n12096), .ZN(N10417) );
  AOI22D1BWP30P140LVT U16822 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1681]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1553]), .ZN(n12103) );
  AOI22D1BWP30P140LVT U16823 ( .A1(n12161), .A2(
        inner_first_stage_data_reg[1713]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1617]), .ZN(n12102) );
  AOI22D1BWP30P140LVT U16824 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1777]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1649]), .ZN(n12101) );
  AOI22D1BWP30P140LVT U16825 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1745]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1585]), .ZN(n12100) );
  ND4D1BWP30P140LVT U16826 ( .A1(n12103), .A2(n12102), .A3(n12101), .A4(n12100), .ZN(N10418) );
  AOI22D1BWP30P140LVT U16827 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1682]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1554]), .ZN(n12107) );
  AOI22D1BWP30P140LVT U16828 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1778]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1650]), .ZN(n12106) );
  AOI22D1BWP30P140LVT U16829 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1586]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1714]), .ZN(n12105) );
  AOI22D1BWP30P140LVT U16830 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1746]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1618]), .ZN(n12104) );
  ND4D1BWP30P140LVT U16831 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(N10419) );
  AOI22D1BWP30P140LVT U16832 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1683]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1555]), .ZN(n12111) );
  AOI22D1BWP30P140LVT U16833 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1779]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1715]), .ZN(n12110) );
  AOI22D1BWP30P140LVT U16834 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1587]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1619]), .ZN(n12109) );
  AOI22D1BWP30P140LVT U16835 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1747]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1651]), .ZN(n12108) );
  ND4D1BWP30P140LVT U16836 ( .A1(n12111), .A2(n12110), .A3(n12109), .A4(n12108), .ZN(N10420) );
  AOI22D1BWP30P140LVT U16837 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1684]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1556]), .ZN(n12115) );
  AOI22D1BWP30P140LVT U16838 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1588]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1652]), .ZN(n12114) );
  AOI22D1BWP30P140LVT U16839 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1748]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1780]), .ZN(n12113) );
  AOI22D1BWP30P140LVT U16840 ( .A1(n12161), .A2(
        inner_first_stage_data_reg[1716]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1620]), .ZN(n12112) );
  ND4D1BWP30P140LVT U16841 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(N10421) );
  AOI22D1BWP30P140LVT U16842 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1685]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1557]), .ZN(n12119) );
  AOI22D1BWP30P140LVT U16843 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1781]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1717]), .ZN(n12118) );
  AOI22D1BWP30P140LVT U16844 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1749]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1589]), .ZN(n12117) );
  AOI22D1BWP30P140LVT U16845 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1653]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1621]), .ZN(n12116) );
  ND4D1BWP30P140LVT U16846 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(N10422) );
  AOI22D1BWP30P140LVT U16847 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1686]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1558]), .ZN(n12123) );
  AOI22D1BWP30P140LVT U16848 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1750]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1622]), .ZN(n12122) );
  AOI22D1BWP30P140LVT U16849 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1782]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1718]), .ZN(n12121) );
  AOI22D1BWP30P140LVT U16850 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1590]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1654]), .ZN(n12120) );
  ND4D1BWP30P140LVT U16851 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(N10423) );
  AOI22D1BWP30P140LVT U16852 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1687]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1559]), .ZN(n12127) );
  AOI22D1BWP30P140LVT U16853 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1655]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1623]), .ZN(n12126) );
  AOI22D1BWP30P140LVT U16854 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1783]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1591]), .ZN(n12125) );
  AOI22D1BWP30P140LVT U16855 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1751]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1719]), .ZN(n12124) );
  ND4D1BWP30P140LVT U16856 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(N10424) );
  AOI22D1BWP30P140LVT U16857 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1688]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1560]), .ZN(n12131) );
  AOI22D1BWP30P140LVT U16858 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1752]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1784]), .ZN(n12130) );
  AOI22D1BWP30P140LVT U16859 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1656]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1624]), .ZN(n12129) );
  AOI22D1BWP30P140LVT U16860 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1592]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1720]), .ZN(n12128) );
  ND4D1BWP30P140LVT U16861 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(N10425) );
  AOI22D1BWP30P140LVT U16862 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1689]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1561]), .ZN(n12135) );
  AOI22D1BWP30P140LVT U16863 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1785]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1593]), .ZN(n12134) );
  AOI22D1BWP30P140LVT U16864 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1753]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1625]), .ZN(n12133) );
  AOI22D1BWP30P140LVT U16865 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1657]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1721]), .ZN(n12132) );
  ND4D1BWP30P140LVT U16866 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(N10426) );
  AOI22D1BWP30P140LVT U16867 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1690]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1562]), .ZN(n12139) );
  AOI22D1BWP30P140LVT U16868 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1754]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1786]), .ZN(n12138) );
  AOI22D1BWP30P140LVT U16869 ( .A1(n12161), .A2(
        inner_first_stage_data_reg[1722]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1626]), .ZN(n12137) );
  AOI22D1BWP30P140LVT U16870 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1594]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1658]), .ZN(n12136) );
  ND4D1BWP30P140LVT U16871 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(N10427) );
  AOI22D1BWP30P140LVT U16872 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1691]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1563]), .ZN(n12143) );
  AOI22D1BWP30P140LVT U16873 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1787]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1627]), .ZN(n12142) );
  AOI22D1BWP30P140LVT U16874 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1659]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1723]), .ZN(n12141) );
  AOI22D1BWP30P140LVT U16875 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1755]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1595]), .ZN(n12140) );
  ND4D1BWP30P140LVT U16876 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n12140), .ZN(N10428) );
  AOI22D1BWP30P140LVT U16877 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1692]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1564]), .ZN(n12147) );
  AOI22D1BWP30P140LVT U16878 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1596]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1724]), .ZN(n12146) );
  AOI22D1BWP30P140LVT U16879 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1788]), .B1(n12158), .B2(
        inner_first_stage_data_reg[1660]), .ZN(n12145) );
  AOI22D1BWP30P140LVT U16880 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1756]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1628]), .ZN(n12144) );
  ND4D1BWP30P140LVT U16881 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(N10429) );
  AOI22D1BWP30P140LVT U16882 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1693]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1565]), .ZN(n12151) );
  AOI22D1BWP30P140LVT U16883 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1757]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1725]), .ZN(n12150) );
  AOI22D1BWP30P140LVT U16884 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1789]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1597]), .ZN(n12149) );
  AOI22D1BWP30P140LVT U16885 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1661]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1629]), .ZN(n12148) );
  ND4D1BWP30P140LVT U16886 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(N10430) );
  AOI22D1BWP30P140LVT U16887 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1694]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1566]), .ZN(n12155) );
  AOI22D1BWP30P140LVT U16888 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1662]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1726]), .ZN(n12154) );
  AOI22D1BWP30P140LVT U16889 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1758]), .B1(n12162), .B2(
        inner_first_stage_data_reg[1598]), .ZN(n12153) );
  AOI22D1BWP30P140LVT U16890 ( .A1(n12159), .A2(
        inner_first_stage_data_reg[1790]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1630]), .ZN(n12152) );
  ND4D1BWP30P140LVT U16891 ( .A1(n12155), .A2(n12154), .A3(n12153), .A4(n12152), .ZN(N10431) );
  AOI22D1BWP30P140LVT U16892 ( .A1(n12156), .A2(
        inner_first_stage_data_reg[1695]), .B1(n7376), .B2(
        inner_first_stage_data_reg[1567]), .ZN(n12166) );
  AOI22D1BWP30P140LVT U16893 ( .A1(n12158), .A2(
        inner_first_stage_data_reg[1663]), .B1(n12157), .B2(
        inner_first_stage_data_reg[1631]), .ZN(n12165) );
  AOI22D1BWP30P140LVT U16894 ( .A1(n12160), .A2(
        inner_first_stage_data_reg[1759]), .B1(n12159), .B2(
        inner_first_stage_data_reg[1791]), .ZN(n12164) );
  AOI22D1BWP30P140LVT U16895 ( .A1(n12162), .A2(
        inner_first_stage_data_reg[1599]), .B1(n12161), .B2(
        inner_first_stage_data_reg[1727]), .ZN(n12163) );
  ND4D1BWP30P140LVT U16896 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(N10432) );
  AOI22D1BWP30P140LVT U16897 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1792]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1824]), .ZN(n12170) );
  AOI22D1BWP30P140LVT U16898 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1856]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1952]), .ZN(n12169) );
  AOI22D1BWP30P140LVT U16899 ( .A1(n12291), .A2(
        inner_first_stage_data_reg[1888]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1920]), .ZN(n12168) );
  AOI22D1BWP30P140LVT U16900 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2016]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1984]), .ZN(n12167) );
  ND4D1BWP30P140LVT U16901 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(N11251) );
  AOI22D1BWP30P140LVT U16902 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1857]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1921]), .ZN(n12174) );
  AOI22D1BWP30P140LVT U16903 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1825]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1889]), .ZN(n12173) );
  AOI22D1BWP30P140LVT U16904 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1793]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1953]), .ZN(n12172) );
  AOI22D1BWP30P140LVT U16905 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2017]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1985]), .ZN(n12171) );
  ND4D1BWP30P140LVT U16906 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(N11252) );
  AOI22D1BWP30P140LVT U16907 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1954]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1922]), .ZN(n12178) );
  AOI22D1BWP30P140LVT U16908 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1858]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1890]), .ZN(n12177) );
  AOI22D1BWP30P140LVT U16909 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1794]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1826]), .ZN(n12176) );
  AOI22D1BWP30P140LVT U16910 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2018]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1986]), .ZN(n12175) );
  ND4D1BWP30P140LVT U16911 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(N11253) );
  AOI22D1BWP30P140LVT U16912 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1859]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1955]), .ZN(n12182) );
  AOI22D1BWP30P140LVT U16913 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1795]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1827]), .ZN(n12181) );
  AOI22D1BWP30P140LVT U16914 ( .A1(n12291), .A2(
        inner_first_stage_data_reg[1891]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1923]), .ZN(n12180) );
  AOI22D1BWP30P140LVT U16915 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2019]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1987]), .ZN(n12179) );
  ND4D1BWP30P140LVT U16916 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(N11254) );
  AOI22D1BWP30P140LVT U16917 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1956]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1924]), .ZN(n12186) );
  AOI22D1BWP30P140LVT U16918 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1828]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1892]), .ZN(n12185) );
  AOI22D1BWP30P140LVT U16919 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1796]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1860]), .ZN(n12184) );
  AOI22D1BWP30P140LVT U16920 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2020]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1988]), .ZN(n12183) );
  ND4D1BWP30P140LVT U16921 ( .A1(n12186), .A2(n12185), .A3(n12184), .A4(n12183), .ZN(N11255) );
  AOI22D1BWP30P140LVT U16922 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1797]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1893]), .ZN(n12190) );
  AOI22D1BWP30P140LVT U16923 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1829]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1925]), .ZN(n12189) );
  AOI22D1BWP30P140LVT U16924 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1861]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1957]), .ZN(n12188) );
  AOI22D1BWP30P140LVT U16925 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2021]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1989]), .ZN(n12187) );
  ND4D1BWP30P140LVT U16926 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(N11256) );
  AOI22D1BWP30P140LVT U16927 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1958]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1926]), .ZN(n12194) );
  AOI22D1BWP30P140LVT U16928 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1830]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1862]), .ZN(n12193) );
  AOI22D1BWP30P140LVT U16929 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1798]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1894]), .ZN(n12192) );
  AOI22D1BWP30P140LVT U16930 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2022]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1990]), .ZN(n12191) );
  ND4D1BWP30P140LVT U16931 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(N11257) );
  AOI22D1BWP30P140LVT U16932 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1863]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1959]), .ZN(n12198) );
  AOI22D1BWP30P140LVT U16933 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1799]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1831]), .ZN(n12197) );
  AOI22D1BWP30P140LVT U16934 ( .A1(n12291), .A2(
        inner_first_stage_data_reg[1895]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1927]), .ZN(n12196) );
  AOI22D1BWP30P140LVT U16935 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2023]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1991]), .ZN(n12195) );
  ND4D1BWP30P140LVT U16936 ( .A1(n12198), .A2(n12197), .A3(n12196), .A4(n12195), .ZN(N11258) );
  AOI22D1BWP30P140LVT U16937 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1800]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1960]), .ZN(n12202) );
  AOI22D1BWP30P140LVT U16938 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1864]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1896]), .ZN(n12201) );
  AOI22D1BWP30P140LVT U16939 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1832]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1928]), .ZN(n12200) );
  AOI22D1BWP30P140LVT U16940 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2024]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1992]), .ZN(n12199) );
  ND4D1BWP30P140LVT U16941 ( .A1(n12202), .A2(n12201), .A3(n12200), .A4(n12199), .ZN(N11259) );
  AOI22D1BWP30P140LVT U16942 ( .A1(n12291), .A2(
        inner_first_stage_data_reg[1897]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1929]), .ZN(n12206) );
  AOI22D1BWP30P140LVT U16943 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1801]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1833]), .ZN(n12205) );
  AOI22D1BWP30P140LVT U16944 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1865]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1961]), .ZN(n12204) );
  AOI22D1BWP30P140LVT U16945 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2025]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1993]), .ZN(n12203) );
  ND4D1BWP30P140LVT U16946 ( .A1(n12206), .A2(n12205), .A3(n12204), .A4(n12203), .ZN(N11260) );
  AOI22D1BWP30P140LVT U16947 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1866]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1898]), .ZN(n12210) );
  AOI22D1BWP30P140LVT U16948 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1962]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1930]), .ZN(n12209) );
  AOI22D1BWP30P140LVT U16949 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1802]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1834]), .ZN(n12208) );
  AOI22D1BWP30P140LVT U16950 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2026]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1994]), .ZN(n12207) );
  ND4D1BWP30P140LVT U16951 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(N11261) );
  AOI22D1BWP30P140LVT U16952 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1803]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1963]), .ZN(n12214) );
  AOI22D1BWP30P140LVT U16953 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1835]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1931]), .ZN(n12213) );
  AOI22D1BWP30P140LVT U16954 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1867]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1899]), .ZN(n12212) );
  AOI22D1BWP30P140LVT U16955 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2027]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1995]), .ZN(n12211) );
  ND4D1BWP30P140LVT U16956 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(N11262) );
  AOI22D1BWP30P140LVT U16957 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1964]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1900]), .ZN(n12218) );
  AOI22D1BWP30P140LVT U16958 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1804]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1868]), .ZN(n12217) );
  AOI22D1BWP30P140LVT U16959 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1836]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1932]), .ZN(n12216) );
  AOI22D1BWP30P140LVT U16960 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2028]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1996]), .ZN(n12215) );
  ND4D1BWP30P140LVT U16961 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(N11263) );
  AOI22D1BWP30P140LVT U16962 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1965]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1901]), .ZN(n12222) );
  AOI22D1BWP30P140LVT U16963 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1837]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1869]), .ZN(n12221) );
  AOI22D1BWP30P140LVT U16964 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1805]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1933]), .ZN(n12220) );
  AOI22D1BWP30P140LVT U16965 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2029]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1997]), .ZN(n12219) );
  ND4D1BWP30P140LVT U16966 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(N11264) );
  AOI22D1BWP30P140LVT U16967 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1806]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1902]), .ZN(n12226) );
  AOI22D1BWP30P140LVT U16968 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1838]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1966]), .ZN(n12225) );
  AOI22D1BWP30P140LVT U16969 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1870]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1934]), .ZN(n12224) );
  AOI22D1BWP30P140LVT U16970 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2030]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1998]), .ZN(n12223) );
  ND4D1BWP30P140LVT U16971 ( .A1(n12226), .A2(n12225), .A3(n12224), .A4(n12223), .ZN(N11265) );
  AOI22D1BWP30P140LVT U16972 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1967]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1935]), .ZN(n12230) );
  AOI22D1BWP30P140LVT U16973 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1807]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1903]), .ZN(n12229) );
  AOI22D1BWP30P140LVT U16974 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1839]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1871]), .ZN(n12228) );
  AOI22D1BWP30P140LVT U16975 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2031]), .B1(n6211), .B2(
        inner_first_stage_data_reg[1999]), .ZN(n12227) );
  ND4D1BWP30P140LVT U16976 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(N11266) );
  AOI22D1BWP30P140LVT U16977 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1840]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1872]), .ZN(n12234) );
  AOI22D1BWP30P140LVT U16978 ( .A1(n12291), .A2(
        inner_first_stage_data_reg[1904]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1936]), .ZN(n12233) );
  AOI22D1BWP30P140LVT U16979 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1808]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1968]), .ZN(n12232) );
  AOI22D1BWP30P140LVT U16980 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2032]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2000]), .ZN(n12231) );
  ND4D1BWP30P140LVT U16981 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(N11267) );
  AOI22D1BWP30P140LVT U16982 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1841]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1873]), .ZN(n12238) );
  AOI22D1BWP30P140LVT U16983 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1969]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1937]), .ZN(n12237) );
  AOI22D1BWP30P140LVT U16984 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1809]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1905]), .ZN(n12236) );
  AOI22D1BWP30P140LVT U16985 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2033]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2001]), .ZN(n12235) );
  ND4D1BWP30P140LVT U16986 ( .A1(n12238), .A2(n12237), .A3(n12236), .A4(n12235), .ZN(N11268) );
  AOI22D1BWP30P140LVT U16987 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1810]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1842]), .ZN(n12242) );
  AOI22D1BWP30P140LVT U16988 ( .A1(n12291), .A2(
        inner_first_stage_data_reg[1906]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1938]), .ZN(n12241) );
  AOI22D1BWP30P140LVT U16989 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1874]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1970]), .ZN(n12240) );
  AOI22D1BWP30P140LVT U16990 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2034]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2002]), .ZN(n12239) );
  ND4D1BWP30P140LVT U16991 ( .A1(n12242), .A2(n12241), .A3(n12240), .A4(n12239), .ZN(N11269) );
  AOI22D1BWP30P140LVT U16992 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1843]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1907]), .ZN(n12246) );
  AOI22D1BWP30P140LVT U16993 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1811]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1939]), .ZN(n12245) );
  AOI22D1BWP30P140LVT U16994 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1875]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1971]), .ZN(n12244) );
  AOI22D1BWP30P140LVT U16995 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2035]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2003]), .ZN(n12243) );
  ND4D1BWP30P140LVT U16996 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(N11270) );
  AOI22D1BWP30P140LVT U16997 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1812]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1844]), .ZN(n12250) );
  AOI22D1BWP30P140LVT U16998 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1876]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1908]), .ZN(n12249) );
  AOI22D1BWP30P140LVT U16999 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1972]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1940]), .ZN(n12248) );
  AOI22D1BWP30P140LVT U17000 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2036]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2004]), .ZN(n12247) );
  ND4D1BWP30P140LVT U17001 ( .A1(n12250), .A2(n12249), .A3(n12248), .A4(n12247), .ZN(N11271) );
  AOI22D1BWP30P140LVT U17002 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1813]), .B1(n12296), .B2(
        inner_first_stage_data_reg[1845]), .ZN(n12254) );
  AOI22D1BWP30P140LVT U17003 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1973]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1941]), .ZN(n12253) );
  AOI22D1BWP30P140LVT U17004 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1877]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1909]), .ZN(n12252) );
  AOI22D1BWP30P140LVT U17005 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2037]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2005]), .ZN(n12251) );
  ND4D1BWP30P140LVT U17006 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(N11272) );
  AOI22D1BWP30P140LVT U17007 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1814]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1910]), .ZN(n12258) );
  AOI22D1BWP30P140LVT U17008 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1846]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1942]), .ZN(n12257) );
  AOI22D1BWP30P140LVT U17009 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1878]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1974]), .ZN(n12256) );
  AOI22D1BWP30P140LVT U17010 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2038]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2006]), .ZN(n12255) );
  ND4D1BWP30P140LVT U17011 ( .A1(n12258), .A2(n12257), .A3(n12256), .A4(n12255), .ZN(N11273) );
  AOI22D1BWP30P140LVT U17012 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1847]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1879]), .ZN(n12262) );
  AOI22D1BWP30P140LVT U17013 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1975]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1943]), .ZN(n12261) );
  AOI22D1BWP30P140LVT U17014 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1815]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1911]), .ZN(n12260) );
  AOI22D1BWP30P140LVT U17015 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2039]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2007]), .ZN(n12259) );
  ND4D1BWP30P140LVT U17016 ( .A1(n12262), .A2(n12261), .A3(n12260), .A4(n12259), .ZN(N11274) );
  AOI22D1BWP30P140LVT U17017 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1880]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1976]), .ZN(n12266) );
  AOI22D1BWP30P140LVT U17018 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1848]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1944]), .ZN(n12265) );
  AOI22D1BWP30P140LVT U17019 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1816]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1912]), .ZN(n12264) );
  AOI22D1BWP30P140LVT U17020 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2040]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2008]), .ZN(n12263) );
  ND4D1BWP30P140LVT U17021 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(N11275) );
  AOI22D1BWP30P140LVT U17022 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1817]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1977]), .ZN(n12270) );
  AOI22D1BWP30P140LVT U17023 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1881]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1913]), .ZN(n12269) );
  AOI22D1BWP30P140LVT U17024 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1849]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1945]), .ZN(n12268) );
  AOI22D1BWP30P140LVT U17025 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2041]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2009]), .ZN(n12267) );
  ND4D1BWP30P140LVT U17026 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(N11276) );
  AOI22D1BWP30P140LVT U17027 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1978]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1914]), .ZN(n12274) );
  AOI22D1BWP30P140LVT U17028 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1850]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1882]), .ZN(n12273) );
  AOI22D1BWP30P140LVT U17029 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1818]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1946]), .ZN(n12272) );
  AOI22D1BWP30P140LVT U17030 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2042]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2010]), .ZN(n12271) );
  ND4D1BWP30P140LVT U17031 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(N11277) );
  AOI22D1BWP30P140LVT U17032 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1819]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1947]), .ZN(n12278) );
  AOI22D1BWP30P140LVT U17033 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1851]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1883]), .ZN(n12277) );
  AOI22D1BWP30P140LVT U17034 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1979]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1915]), .ZN(n12276) );
  AOI22D1BWP30P140LVT U17035 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2043]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2011]), .ZN(n12275) );
  ND4D1BWP30P140LVT U17036 ( .A1(n12278), .A2(n12277), .A3(n12276), .A4(n12275), .ZN(N11278) );
  AOI22D1BWP30P140LVT U17037 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1820]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1948]), .ZN(n12282) );
  AOI22D1BWP30P140LVT U17038 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1852]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1884]), .ZN(n12281) );
  AOI22D1BWP30P140LVT U17039 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1980]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1916]), .ZN(n12280) );
  AOI22D1BWP30P140LVT U17040 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2044]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2012]), .ZN(n12279) );
  ND4D1BWP30P140LVT U17041 ( .A1(n12282), .A2(n12281), .A3(n12280), .A4(n12279), .ZN(N11279) );
  AOI22D1BWP30P140LVT U17042 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1821]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1917]), .ZN(n12286) );
  AOI22D1BWP30P140LVT U17043 ( .A1(n12293), .A2(
        inner_first_stage_data_reg[1885]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1981]), .ZN(n12285) );
  AOI22D1BWP30P140LVT U17044 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1853]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1949]), .ZN(n12284) );
  AOI22D1BWP30P140LVT U17045 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2045]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2013]), .ZN(n12283) );
  ND4D1BWP30P140LVT U17046 ( .A1(n12286), .A2(n12285), .A3(n12284), .A4(n12283), .ZN(N11280) );
  AOI22D1BWP30P140LVT U17047 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1854]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1886]), .ZN(n12290) );
  AOI22D1BWP30P140LVT U17048 ( .A1(n12291), .A2(
        inner_first_stage_data_reg[1918]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1950]), .ZN(n12289) );
  AOI22D1BWP30P140LVT U17049 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1822]), .B1(n12292), .B2(
        inner_first_stage_data_reg[1982]), .ZN(n12288) );
  AOI22D1BWP30P140LVT U17050 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2046]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2014]), .ZN(n12287) );
  ND4D1BWP30P140LVT U17051 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(N11281) );
  AOI22D1BWP30P140LVT U17052 ( .A1(n12292), .A2(
        inner_first_stage_data_reg[1983]), .B1(n12291), .B2(
        inner_first_stage_data_reg[1919]), .ZN(n12301) );
  AOI22D1BWP30P140LVT U17053 ( .A1(n12294), .A2(
        inner_first_stage_data_reg[1823]), .B1(n12293), .B2(
        inner_first_stage_data_reg[1887]), .ZN(n12300) );
  AOI22D1BWP30P140LVT U17054 ( .A1(n12296), .A2(
        inner_first_stage_data_reg[1855]), .B1(n12295), .B2(
        inner_first_stage_data_reg[1951]), .ZN(n12299) );
  AOI22D1BWP30P140LVT U17055 ( .A1(n12297), .A2(
        inner_first_stage_data_reg[2047]), .B1(n6211), .B2(
        inner_first_stage_data_reg[2015]), .ZN(n12298) );
  ND4D1BWP30P140LVT U17056 ( .A1(n12301), .A2(n12300), .A3(n12299), .A4(n12298), .ZN(N11282) );
endmodule

