
module crossbar_one_hot_comb_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA32 ( 
        i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [31:0] i_valid;
  input [1023:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [255:0] i_cmd;
  input i_en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205;

  INVD2BWP30P140LVT U3 ( .I(n3961), .ZN(n3348) );
  NR3D1P5BWP30P140LVT U4 ( .A1(n5444), .A2(n1985), .A3(n1987), .ZN(n1986) );
  INR3D1BWP30P140LVT U5 ( .A1(i_cmd[212]), .B1(n5461), .B2(n1987), .ZN(n2638)
         );
  INR3D1BWP30P140LVT U6 ( .A1(i_cmd[220]), .B1(n5457), .B2(n1987), .ZN(n2639)
         );
  CKBD1BWP30P140LVT U7 ( .I(n615), .Z(n1264) );
  CKBD1BWP30P140LVT U8 ( .I(n606), .Z(n1254) );
  CKBD1BWP30P140LVT U9 ( .I(n4105), .Z(n4721) );
  INVD1BWP30P140LVT U10 ( .I(n75), .ZN(n1924) );
  INVD1BWP30P140LVT U11 ( .I(n69), .ZN(n1912) );
  NR3D1P5BWP30P140LVT U12 ( .A1(n5473), .A2(n4072), .A3(n4071), .ZN(n4073) );
  INVD2BWP30P140LVT U13 ( .I(n1241), .ZN(n37) );
  INVD2BWP30P140LVT U14 ( .I(n1), .ZN(n2) );
  INVD1BWP30P140LVT U15 ( .I(n3856), .ZN(n4021) );
  INVD3BWP30P140LVT U16 ( .I(n3984), .ZN(n4020) );
  INVD3BWP30P140LVT U17 ( .I(n4046), .ZN(n4006) );
  INVD1P5BWP30P140LVT U18 ( .I(n3878), .ZN(n3347) );
  INR3D1BWP30P140LVT U19 ( .A1(i_cmd[204]), .B1(n5459), .B2(n1987), .ZN(n2635)
         );
  NR3D1P5BWP30P140LVT U20 ( .A1(n5455), .A2(n1988), .A3(n1990), .ZN(n1989) );
  NR3D1P5BWP30P140LVT U21 ( .A1(n5455), .A2(n1305), .A3(n1308), .ZN(n1944) );
  INR3D1BWP30P140LVT U22 ( .A1(i_cmd[209]), .B1(n5461), .B2(n619), .ZN(n600)
         );
  INR3D1BWP30P140LVT U23 ( .A1(i_cmd[217]), .B1(n619), .B2(n5457), .ZN(n617)
         );
  NR3D1P5BWP30P140LVT U24 ( .A1(n126), .A2(n619), .A3(n5444), .ZN(n1253) );
  INR3D2BWP30P140LVT U25 ( .A1(i_cmd[19]), .B1(n5451), .B2(n1298), .ZN(n1925)
         );
  INR3D2BWP30P140LVT U26 ( .A1(i_cmd[27]), .B1(n5446), .B2(n1298), .ZN(n1936)
         );
  NR3D1P5BWP30P140LVT U27 ( .A1(n5450), .A2(n1970), .A3(n1969), .ZN(n2624) );
  CKBD1BWP30P140LVT U28 ( .I(n1243), .Z(n117) );
  AN3D1BWP30P140LVT U29 ( .A1(i_valid[13]), .A2(i_cmd[109]), .A3(n2680), .Z(
        n3303) );
  INVD1BWP30P140LVT U30 ( .I(n44), .ZN(n4025) );
  CKBD1BWP30P140LVT U31 ( .I(n1235), .Z(n25) );
  NR3D1P5BWP30P140LVT U32 ( .A1(n5477), .A2(n2681), .A3(n2682), .ZN(n3331) );
  NR3D1P5BWP30P140LVT U33 ( .A1(n5477), .A2(n129), .A3(n5480), .ZN(n6181) );
  NR3D1P5BWP30P140LVT U34 ( .A1(n5450), .A2(n196), .A3(n579), .ZN(n5398) );
  NR3D1P5BWP30P140LVT U35 ( .A1(n5473), .A2(n5472), .A3(n5489), .ZN(n5474) );
  NR3D1P5BWP30P140LVT U36 ( .A1(n114), .A2(n5457), .A3(n2670), .ZN(n113) );
  NR3D1P5BWP30P140LVT U37 ( .A1(n5493), .A2(n2652), .A3(n2651), .ZN(n2935) );
  INVD3BWP30P140LVT U38 ( .I(n3267), .ZN(n3329) );
  INVD1BWP30P140LVT U39 ( .I(n26), .ZN(n3301) );
  INVD1BWP30P140LVT U40 ( .I(n3246), .ZN(n3330) );
  NR3D1P5BWP30P140LVT U41 ( .A1(n5476), .A2(n130), .A3(n3370), .ZN(n4022) );
  ND3D1BWP30P140LVT U42 ( .A1(n420), .A2(n419), .A3(n418), .ZN(n1987) );
  NR3D1P5BWP30P140LVT U43 ( .A1(n5444), .A2(n3364), .A3(n3363), .ZN(n4027) );
  INR3D1BWP30P140LVT U44 ( .A1(i_cmd[202]), .B1(n5459), .B2(n3363), .ZN(n4024)
         );
  INR3D2BWP30P140LVT U45 ( .A1(i_cmd[63]), .B1(n5471), .B2(n5495), .ZN(n6160)
         );
  NR3D1P5BWP30P140LVT U46 ( .A1(n5493), .A2(n122), .A3(n5495), .ZN(n6190) );
  INVD0P7BWP30P140LVT U47 ( .I(n3982), .ZN(n3447) );
  NR3D0P7BWP30P140LVT U48 ( .A1(n5470), .A2(n1286), .A3(n1299), .ZN(n1934) );
  ND3D2BWP30P140LVT U49 ( .A1(n550), .A2(n549), .A3(n551), .ZN(n619) );
  INR3D1BWP30P140LVT U50 ( .A1(i_cmd[155]), .B1(n5478), .B2(n1296), .ZN(n1910)
         );
  INR3D1BWP30P140LVT U51 ( .A1(i_cmd[17]), .B1(n590), .B2(n5451), .ZN(n1229)
         );
  ND3D3BWP30P140LVT U52 ( .A1(n562), .A2(n561), .A3(n560), .ZN(n620) );
  OR3D1BWP30P140LVT U53 ( .A1(n277), .A2(n276), .A3(n275), .Z(n5495) );
  NR3D1P5BWP30P140LVT U54 ( .A1(n5444), .A2(n2671), .A3(n2670), .ZN(n3307) );
  ND3OPTPAD4BWP30P140LVT U55 ( .A1(n82), .A2(n460), .A3(n463), .ZN(n1299) );
  NR2OPTPAD1BWP30P140LVT U56 ( .A1(n407), .A2(n406), .ZN(n415) );
  ND3D1BWP30P140LVT U57 ( .A1(n513), .A2(n521), .A3(n505), .ZN(n3362) );
  ND3D2BWP30P140LVT U58 ( .A1(n371), .A2(n368), .A3(n369), .ZN(n2670) );
  ND3D1BWP30P140LVT U59 ( .A1(n473), .A2(n455), .A3(n456), .ZN(n1298) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n367), .A2(n60), .Z(n371) );
  IND4D1BWP30P140LVT U61 ( .A1(n365), .B1(n364), .B2(n363), .B3(n362), .ZN(
        n2667) );
  INR2D2BWP30P140LVT U62 ( .A1(n118), .B1(n453), .ZN(n473) );
  NR3OPTPAD2BWP30P140LVT U63 ( .A1(n13), .A2(n559), .A3(n555), .ZN(n568) );
  CKND2D2BWP30P140LVT U64 ( .A1(n452), .A2(n451), .ZN(n453) );
  NR2OPTPAD1BWP30P140LVT U65 ( .A1(n358), .A2(n357), .ZN(n367) );
  NR2D1BWP30P140LVT U66 ( .A1(n426), .A2(n547), .ZN(n412) );
  NR2OPTPAD1BWP30P140LVT U67 ( .A1(n472), .A2(n449), .ZN(n451) );
  INVD1BWP30P140LVT U68 ( .I(n460), .ZN(n86) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n376), .A2(i_en), .Z(n358) );
  INVD1BWP30P140LVT U70 ( .I(n81), .ZN(n449) );
  NR2D2BWP30P140LVT U71 ( .A1(n553), .A2(n549), .ZN(n565) );
  IND2D1BWP30P140LVT U72 ( .A1(n186), .B1(n185), .ZN(n213) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n462), .A2(i_en), .Z(n461) );
  NR2D1BWP30P140LVT U74 ( .A1(n501), .A2(n503), .ZN(n514) );
  NR2D1BWP30P140LVT U75 ( .A1(n547), .A2(n261), .ZN(n262) );
  NR2D1BWP30P140LVT U76 ( .A1(n547), .A2(n259), .ZN(n263) );
  INR2D1BWP30P140LVT U77 ( .A1(n375), .B1(n547), .ZN(n355) );
  NR2OPTIBD6BWP30P140LVT U78 ( .A1(n545), .A2(n547), .ZN(n562) );
  NR2D1BWP30P140LVT U79 ( .A1(n465), .A2(n467), .ZN(n460) );
  NR2D1BWP30P140LVT U80 ( .A1(n547), .A2(n268), .ZN(n281) );
  INR2D1BWP30P140LVT U81 ( .A1(i_en), .B1(n468), .ZN(n465) );
  MUX2D0BWP30P140LVT U82 ( .I0(n250), .I1(n145), .S(i_cmd[199]), .Z(n280) );
  MUX2D0BWP30P140LVT U83 ( .I0(n337), .I1(n149), .S(i_cmd[197]), .Z(n372) );
  MUX2D0BWP30P140LVT U84 ( .I0(n248), .I1(n144), .S(i_cmd[167]), .Z(n268) );
  NR2D1BWP30P140LVT U85 ( .A1(n511), .A2(n497), .ZN(n507) );
  INR2D1BWP30P140LVT U86 ( .A1(i_en), .B1(n464), .ZN(n467) );
  NR2D1BWP30P140LVT U87 ( .A1(n86), .A2(n461), .ZN(n452) );
  INR3D2BWP30P140LVT U88 ( .A1(i_cmd[11]), .B1(n5442), .B2(n1298), .ZN(n1914)
         );
  BUFFD2BWP30P140LVT U89 ( .I(n616), .Z(n5) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n366), .A2(i_en), .Z(n360) );
  INVD2BWP30P140LVT U91 ( .I(n3288), .ZN(n3) );
  CKBD1BWP30P140LVT U92 ( .I(n2655), .Z(n3318) );
  INR3D2BWP30P140LVT U93 ( .A1(i_cmd[205]), .B1(n5459), .B2(n2670), .ZN(n3304)
         );
  INR3D2BWP30P140LVT U94 ( .A1(i_cmd[213]), .B1(n5461), .B2(n2670), .ZN(n3316)
         );
  INR3D2BWP30P140LVT U95 ( .A1(i_cmd[55]), .B1(n5495), .B2(n5494), .ZN(n6189)
         );
  INR3D2BWP30P140LVT U96 ( .A1(i_cmd[47]), .B1(n5495), .B2(n5487), .ZN(n5488)
         );
  ND3D1BWP30P140LVT U97 ( .A1(n569), .A2(n11), .A3(n567), .ZN(n590) );
  INVD1BWP30P140LVT U98 ( .I(n1278), .ZN(n1) );
  INVD1BWP30P140LVT U99 ( .I(n117), .ZN(n4) );
  INR3D2BWP30P140LVT U100 ( .A1(i_cmd[18]), .B1(n5451), .B2(n3362), .ZN(n4028)
         );
  INR2D1BWP30P140LVT U101 ( .A1(n415), .B1(n414), .ZN(n418) );
  INVD2BWP30P140LVT U102 ( .I(n451), .ZN(n457) );
  NR2OPTPAD4BWP30P140LVT U103 ( .A1(n546), .A2(n562), .ZN(n558) );
  INVD1BWP30P140LVT U104 ( .I(n507), .ZN(n517) );
  NR2OPTPAD1BWP30P140LVT U105 ( .A1(n281), .A2(n267), .ZN(n285) );
  IND2D1BWP30P140LVT U106 ( .A1(n471), .B1(i_en), .ZN(n81) );
  ND2D1BWP30P140LVT U107 ( .A1(n149), .A2(n336), .ZN(n337) );
  OR3D1BWP30P140LVT U108 ( .A1(i_cmd[83]), .A2(i_cmd[91]), .A3(i_cmd[75]), .Z(
        n445) );
  OR3D1BWP30P140LVT U109 ( .A1(i_cmd[139]), .A2(i_cmd[155]), .A3(i_cmd[147]), 
        .Z(n431) );
  AN4D0BWP30P140LVT U110 ( .A1(n1424), .A2(n1423), .A3(n1422), .A4(n1421), .Z(
        n47) );
  AN4D0BWP30P140LVT U111 ( .A1(n1420), .A2(n1419), .A3(n1418), .A4(n1417), .Z(
        n49) );
  AN4D0BWP30P140LVT U112 ( .A1(n1597), .A2(n1596), .A3(n1595), .A4(n1594), .Z(
        n62) );
  AN4D0BWP30P140LVT U113 ( .A1(n1605), .A2(n1604), .A3(n1603), .A4(n1602), .Z(
        n64) );
  AN4D0BWP30P140LVT U114 ( .A1(n1609), .A2(n1608), .A3(n1607), .A4(n1606), .Z(
        n1610) );
  AN4D0BWP30P140LVT U115 ( .A1(n1428), .A2(n1427), .A3(n1426), .A4(n1425), .Z(
        n48) );
  AN4D0BWP30P140LVT U116 ( .A1(n1601), .A2(n1600), .A3(n1599), .A4(n1598), .Z(
        n63) );
  NR3D1P5BWP30P140LVT U117 ( .A1(n5476), .A2(n139), .A3(n1287), .ZN(n1279) );
  OR3D1BWP30P140LVT U118 ( .A1(n70), .A2(n5481), .A3(n1296), .Z(n69) );
  NR3D1P5BWP30P140LVT U119 ( .A1(n5497), .A2(n1292), .A3(n1295), .ZN(n1293) );
  NR3D1P5BWP30P140LVT U120 ( .A1(n5477), .A2(n4103), .A3(n4102), .ZN(n4722) );
  ND3D2BWP30P140LVT U121 ( .A1(n501), .A2(n500), .A3(n502), .ZN(n3363) );
  NR3D1P5BWP30P140LVT U122 ( .A1(n5493), .A2(n123), .A3(n572), .ZN(n5399) );
  NR3D1P5BWP30P140LVT U123 ( .A1(n5493), .A2(n1958), .A3(n1980), .ZN(n2600) );
  NR3D1P5BWP30P140LVT U124 ( .A1(n5477), .A2(n125), .A3(n1975), .ZN(n2601) );
  INVD1BWP30P140LVT U125 ( .I(n2651), .ZN(n2677) );
  ND3D2BWP30P140LVT U126 ( .A1(n545), .A2(n546), .A3(n560), .ZN(n607) );
  OR3D1BWP30P140LVT U127 ( .A1(n5490), .A2(n2669), .A3(n2668), .Z(n26) );
  NR3D1P5BWP30P140LVT U128 ( .A1(n5450), .A2(n131), .A3(n3362), .ZN(n4038) );
  NR2D1BWP30P140LVT U129 ( .A1(n499), .A2(n498), .ZN(n502) );
  NR3D1P5BWP30P140LVT U130 ( .A1(n5477), .A2(n124), .A3(n578), .ZN(n5414) );
  NR3D1P5BWP30P140LVT U131 ( .A1(n5450), .A2(n2649), .A3(n2656), .ZN(n3319) );
  INR3D2BWP30P140LVT U132 ( .A1(i_cmd[26]), .B1(n5446), .B2(n3362), .ZN(n4026)
         );
  NR3D1P5BWP30P140LVT U133 ( .A1(n5450), .A2(n134), .A3(n4107), .ZN(n4097) );
  NR2D1BWP30P140LVT U134 ( .A1(n450), .A2(n454), .ZN(n470) );
  NR3D1P5BWP30P140LVT U135 ( .A1(n5490), .A2(n3374), .A3(n3381), .ZN(n4048) );
  NR3D1P5BWP30P140LVT U136 ( .A1(n5477), .A2(n3380), .A3(n3384), .ZN(n4052) );
  NR3D1P5BWP30P140LVT U137 ( .A1(n5470), .A2(n3382), .A3(n3381), .ZN(n3383) );
  NR3D1P5BWP30P140LVT U138 ( .A1(n5470), .A2(n4065), .A3(n4071), .ZN(n4066) );
  NR2D1BWP30P140LVT U139 ( .A1(n266), .A2(n265), .ZN(n279) );
  NR3D1P5BWP30P140LVT U140 ( .A1(n5486), .A2(n4069), .A3(n4071), .ZN(n4070) );
  NR3D1P5BWP30P140LVT U141 ( .A1(n5490), .A2(n4067), .A3(n4071), .ZN(n4068) );
  IND3D2BWP30P140LVT U142 ( .A1(n270), .B1(n269), .B2(n283), .ZN(n5453) );
  IND2D2BWP30P140LVT U143 ( .A1(n182), .B1(n211), .ZN(n183) );
  NR3D1P5BWP30P140LVT U144 ( .A1(n522), .A2(n506), .A3(n517), .ZN(n513) );
  INR3D1BWP30P140LVT U145 ( .A1(n331), .B1(n319), .B2(n332), .ZN(n326) );
  INVD1BWP30P140LVT U146 ( .I(n374), .ZN(n356) );
  INR2D2BWP30P140LVT U147 ( .A1(n285), .B1(n284), .ZN(n269) );
  NR2OPTPAD2BWP30P140LVT U148 ( .A1(n475), .A2(n455), .ZN(n459) );
  NR2OPTPAD2BWP30P140LVT U149 ( .A1(n379), .A2(n355), .ZN(n362) );
  INVD4BWP30P140LVT U150 ( .I(n12), .ZN(n455) );
  NR2D3BWP30P140LVT U151 ( .A1(n373), .A2(n368), .ZN(n359) );
  ND2D1BWP30P140LVT U152 ( .A1(i_en), .A2(n329), .ZN(n310) );
  ND2D1BWP30P140LVT U153 ( .A1(i_en), .A2(n424), .ZN(n404) );
  INVD1BWP30P140LVT U154 ( .I(n454), .ZN(n118) );
  ND2D1BWP30P140LVT U155 ( .A1(i_en), .A2(n352), .ZN(n361) );
  INVD1BWP30P140LVT U156 ( .I(n366), .ZN(n60) );
  INVD1BWP30P140LVT U157 ( .I(n518), .ZN(n516) );
  IND2D2BWP30P140LVT U158 ( .A1(n474), .B1(i_en), .ZN(n12) );
  ND2D1BWP30P140LVT U159 ( .A1(i_en), .A2(n277), .ZN(n274) );
  ND2D1BWP30P140LVT U160 ( .A1(n414), .A2(i_en), .ZN(n409) );
  AN4D0BWP30P140LVT U161 ( .A1(n198), .A2(n197), .A3(n187), .A4(n195), .Z(n189) );
  ND4D1BWP30P140LVT U162 ( .A1(n2669), .A2(n2664), .A3(n2650), .A4(n2665), 
        .ZN(n366) );
  OR3D1BWP30P140LVT U163 ( .A1(i_cmd[142]), .A2(i_cmd[158]), .A3(i_cmd[150]), 
        .Z(n299) );
  OR3D1BWP30P140LVT U164 ( .A1(i_cmd[214]), .A2(i_cmd[206]), .A3(i_cmd[222]), 
        .Z(n290) );
  OR3D1BWP30P140LVT U165 ( .A1(i_cmd[84]), .A2(i_cmd[92]), .A3(i_cmd[76]), .Z(
        n385) );
  OR3D1BWP30P140LVT U166 ( .A1(i_cmd[182]), .A2(i_cmd[190]), .A3(i_cmd[174]), 
        .Z(n287) );
  OR3D1BWP30P140LVT U167 ( .A1(i_cmd[180]), .A2(i_cmd[188]), .A3(i_cmd[172]), 
        .Z(n392) );
  OR3D1BWP30P140LVT U168 ( .A1(i_cmd[212]), .A2(i_cmd[204]), .A3(i_cmd[220]), 
        .Z(n395) );
  OR3D1BWP30P140LVT U169 ( .A1(i_cmd[112]), .A2(i_cmd[120]), .A3(i_cmd[104]), 
        .Z(n175) );
  OR3D1BWP30P140LVT U170 ( .A1(i_cmd[24]), .A2(i_cmd[8]), .A3(i_cmd[16]), .Z(
        n160) );
  OR3D1BWP30P140LVT U171 ( .A1(i_cmd[208]), .A2(i_cmd[200]), .A3(i_cmd[216]), 
        .Z(n168) );
  INR3D2BWP30P140LVT U172 ( .A1(i_cmd[9]), .B1(n5442), .B2(n590), .ZN(n1232)
         );
  INR3D2BWP30P140LVT U173 ( .A1(i_cmd[9]), .B1(n5442), .B2(n590), .ZN(n103) );
  ND3D1BWP30P140LVT U174 ( .A1(n558), .A2(n555), .A3(n554), .ZN(n616) );
  INVD2BWP30P140LVT U175 ( .I(n228), .ZN(n5411) );
  INVD2BWP30P140LVT U176 ( .I(n5264), .ZN(n5428) );
  IND3D4BWP30P140LVT U177 ( .A1(n409), .B1(n408), .B2(n415), .ZN(n1978) );
  NR3D1P5BWP30P140LVT U178 ( .A1(n5493), .A2(n141), .A3(n4112), .ZN(n4108) );
  NR2OPTPAD1BWP30P140LVT U179 ( .A1(n308), .A2(n321), .ZN(n327) );
  OA211D1BWP30P140LVT U180 ( .A1(n583), .A2(i_cmd[129]), .B(n6), .C(i_en), .Z(
        n559) );
  AO21D1BWP30P140LVT U181 ( .A1(n543), .A2(n544), .B(n582), .Z(n6) );
  NR2D3BWP30P140LVT U182 ( .A1(n219), .A2(n193), .ZN(n211) );
  NR3D1P5BWP30P140LVT U183 ( .A1(n5444), .A2(n221), .A3(n571), .ZN(n5407) );
  INVD2BWP30P140LVT U184 ( .I(n558), .ZN(n13) );
  CKBD1BWP30P140LVT U185 ( .I(n3311), .Z(n7) );
  BUFFD3BWP30P140LVT U186 ( .I(n618), .Z(n1244) );
  MAOI22D1BWP30P140LVT U187 ( .A1(n1231), .A2(i_data_bus[972]), .B1(n4), .B2(
        n8), .ZN(n855) );
  INVD1BWP30P140LVT U188 ( .I(i_data_bus[108]), .ZN(n8) );
  IND4D1BWP30P140LVT U189 ( .A1(n9), .B1(n672), .B2(n671), .B3(n670), .ZN(n688) );
  AO22D1BWP30P140LVT U190 ( .A1(n1241), .A2(i_data_bus[515]), .B1(n1229), .B2(
        i_data_bus[67]), .Z(n9) );
  ND3OPTPAD2BWP30P140LVT U191 ( .A1(n566), .A2(n565), .A3(n564), .ZN(n10) );
  INR3D8BWP30P140LVT U192 ( .A1(n459), .B1(n458), .B2(n457), .ZN(n463) );
  ND3D2BWP30P140LVT U193 ( .A1(i_valid[14]), .A2(i_cmd[117]), .A3(n2680), .ZN(
        n3246) );
  AOI22D1BWP30P140LVT U194 ( .A1(i_data_bus[155]), .A2(n2935), .B1(
        i_data_bus[475]), .B2(n3330), .ZN(n3228) );
  NR3D0P7BWP30P140LVT U195 ( .A1(n13), .A2(n559), .A3(n555), .ZN(n11) );
  INR3D4BWP30P140LVT U196 ( .A1(i_cmd[153]), .B1(n595), .B2(n5478), .ZN(n1240)
         );
  MAOI22D1BWP30P140LVT U197 ( .A1(i_data_bus[928]), .A2(n1242), .B1(n14), .B2(
        n37), .ZN(n587) );
  INVD1BWP30P140LVT U198 ( .I(i_data_bus[512]), .ZN(n14) );
  MAOI22D1BWP30P140LVT U199 ( .A1(n1231), .A2(i_data_bus[988]), .B1(n37), .B2(
        n15), .ZN(n1172) );
  INVD1BWP30P140LVT U200 ( .I(i_data_bus[540]), .ZN(n15) );
  MAOI22D1BWP30P140LVT U201 ( .A1(n594), .A2(i_data_bus[921]), .B1(n30), .B2(
        n16), .ZN(n1111) );
  INVD1BWP30P140LVT U202 ( .I(i_data_bus[569]), .ZN(n16) );
  INVD1BWP30P140LVT U203 ( .I(n1233), .ZN(n30) );
  MAOI22D1BWP30P140LVT U204 ( .A1(n1231), .A2(i_data_bus[962]), .B1(n32), .B2(
        n17), .ZN(n652) );
  INVD1BWP30P140LVT U205 ( .I(i_data_bus[66]), .ZN(n17) );
  INVD1BWP30P140LVT U206 ( .I(n1229), .ZN(n32) );
  MAOI22D1BWP30P140LVT U207 ( .A1(n594), .A2(i_data_bus[905]), .B1(n32), .B2(
        n18), .ZN(n791) );
  INVD1BWP30P140LVT U208 ( .I(i_data_bus[73]), .ZN(n18) );
  INVD1BWP30P140LVT U209 ( .I(n1234), .ZN(n23) );
  INR3D4BWP30P140LVT U210 ( .A1(i_cmd[145]), .B1(n595), .B2(n5481), .ZN(n1234)
         );
  MAOI22D1BWP30P140LVT U211 ( .A1(n594), .A2(i_data_bus[903]), .B1(n37), .B2(
        n19), .ZN(n751) );
  INVD1BWP30P140LVT U212 ( .I(i_data_bus[519]), .ZN(n19) );
  MAOI22D1BWP30P140LVT U213 ( .A1(n1231), .A2(i_data_bus[968]), .B1(n20), .B2(
        n21), .ZN(n772) );
  INVD1BWP30P140LVT U214 ( .I(n25), .ZN(n20) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[8]), .ZN(n21) );
  MAOI22D1BWP30P140LVT U216 ( .A1(n1242), .A2(i_data_bus[958]), .B1(n37), .B2(
        n22), .ZN(n1211) );
  INVD1BWP30P140LVT U217 ( .I(i_data_bus[542]), .ZN(n22) );
  MAOI22D1BWP30P140LVT U218 ( .A1(n594), .A2(i_data_bus[911]), .B1(n23), .B2(
        n24), .ZN(n911) );
  INVD1BWP30P140LVT U219 ( .I(i_data_bus[591]), .ZN(n24) );
  MAOI22D1BWP30P140LVT U220 ( .A1(n1242), .A2(i_data_bus[951]), .B1(n4), .B2(
        n27), .ZN(n1069) );
  INVD1BWP30P140LVT U221 ( .I(i_data_bus[119]), .ZN(n27) );
  MAOI22D1BWP30P140LVT U222 ( .A1(n1231), .A2(i_data_bus[973]), .B1(n30), .B2(
        n28), .ZN(n870) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[557]), .ZN(n28) );
  INR3D4BWP30P140LVT U224 ( .A1(i_cmd[137]), .B1(n5479), .B2(n595), .ZN(n1233)
         );
  MAOI22D1BWP30P140LVT U225 ( .A1(n1242), .A2(i_data_bus[933]), .B1(n4), .B2(
        n29), .ZN(n709) );
  INVD1BWP30P140LVT U226 ( .I(i_data_bus[101]), .ZN(n29) );
  ND3OPTPAD2BWP30P140LVT U227 ( .A1(n564), .A2(n565), .A3(n566), .ZN(n592) );
  MAOI22D1BWP30P140LVT U228 ( .A1(n594), .A2(i_data_bus[927]), .B1(n30), .B2(
        n31), .ZN(n1237) );
  INVD1BWP30P140LVT U229 ( .I(i_data_bus[575]), .ZN(n31) );
  MAOI22D1BWP30P140LVT U230 ( .A1(n594), .A2(i_data_bus[913]), .B1(n32), .B2(
        n33), .ZN(n950) );
  INVD1BWP30P140LVT U231 ( .I(i_data_bus[81]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U232 ( .A1(n6095), .A2(n3961), .B1(i_data_bus[412]), 
        .B2(n4022), .ZN(n3967) );
  INVD1BWP30P140LVT U233 ( .I(n4022), .ZN(n4007) );
  MAOI22D1BWP30P140LVT U234 ( .A1(n1231), .A2(i_data_bus[971]), .B1(n4), .B2(
        n34), .ZN(n829) );
  INVD1BWP30P140LVT U235 ( .I(i_data_bus[107]), .ZN(n34) );
  MAOI22D1BWP30P140LVT U236 ( .A1(n1231), .A2(i_data_bus[967]), .B1(n4), .B2(
        n35), .ZN(n749) );
  INVD1BWP30P140LVT U237 ( .I(i_data_bus[103]), .ZN(n35) );
  MAOI22D1BWP30P140LVT U238 ( .A1(n594), .A2(i_data_bus[922]), .B1(n37), .B2(
        n36), .ZN(n1129) );
  INVD1BWP30P140LVT U239 ( .I(i_data_bus[538]), .ZN(n36) );
  BUFFD2BWP30P140LVT U240 ( .I(n584), .Z(n1241) );
  MAOI22D1BWP30P140LVT U241 ( .A1(n594), .A2(i_data_bus[908]), .B1(n37), .B2(
        n38), .ZN(n849) );
  INVD1BWP30P140LVT U242 ( .I(i_data_bus[524]), .ZN(n38) );
  NR2D2BWP30P140LVT U243 ( .A1(n547), .A2(n280), .ZN(n267) );
  INR3D2BWP30P140LVT U244 ( .A1(n521), .B1(n505), .B2(n522), .ZN(n508) );
  INR2D4BWP30P140LVT U245 ( .A1(n514), .B1(n515), .ZN(n521) );
  INVD1BWP30P140LVT U246 ( .I(n3930), .ZN(n42) );
  MAOI22D1BWP30P140LVT U247 ( .A1(i_data_bus[86]), .A2(n4028), .B1(n39), .B2(
        n41), .ZN(n3830) );
  INVD1BWP30P140LVT U248 ( .I(i_data_bus[118]), .ZN(n39) );
  INVD1BWP30P140LVT U249 ( .I(n4026), .ZN(n41) );
  MAOI22D1BWP30P140LVT U250 ( .A1(i_data_bus[64]), .A2(n4028), .B1(n40), .B2(
        n41), .ZN(n3368) );
  INVD1BWP30P140LVT U251 ( .I(i_data_bus[96]), .ZN(n40) );
  INR2D4BWP30P140LVT U252 ( .A1(n359), .B1(n360), .ZN(n378) );
  IND4D1BWP30P140LVT U253 ( .A1(n42), .B1(n3929), .B2(n3928), .B3(n3927), .ZN(
        o_data_bus[90]) );
  MAOI22D1BWP30P140LVT U254 ( .A1(i_data_bus[74]), .A2(n4028), .B1(n43), .B2(
        n44), .ZN(n3584) );
  INVD1BWP30P140LVT U255 ( .I(i_data_bus[42]), .ZN(n43) );
  IND4D1BWP30P140LVT U256 ( .A1(n1433), .B1(n47), .B2(n48), .B3(n49), .ZN(
        o_data_bus[102]) );
  OR3D1BWP30P140LVT U257 ( .A1(n45), .A2(n5442), .A3(n3362), .Z(n44) );
  INVD1BWP30P140LVT U258 ( .I(i_cmd[10]), .ZN(n45) );
  MAOI22D1BWP30P140LVT U259 ( .A1(i_data_bus[85]), .A2(n1925), .B1(n46), .B2(
        n56), .ZN(n1716) );
  INVD1BWP30P140LVT U260 ( .I(i_data_bus[629]), .ZN(n46) );
  INVD1BWP30P140LVT U261 ( .I(n1910), .ZN(n56) );
  MAOI22D1BWP30P140LVT U262 ( .A1(i_data_bus[73]), .A2(n1925), .B1(n50), .B2(
        n80), .ZN(n1477) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[521]), .ZN(n50) );
  NR3D1P5BWP30P140LVT U264 ( .A1(n5477), .A2(n1284), .A3(n1296), .ZN(n1927) );
  INVD1BWP30P140LVT U265 ( .I(n1927), .ZN(n80) );
  MAOI22D1BWP30P140LVT U266 ( .A1(i_data_bus[108]), .A2(n1936), .B1(n51), .B2(
        n74), .ZN(n1541) );
  INVD1BWP30P140LVT U267 ( .I(i_data_bus[972]), .ZN(n51) );
  INVD1BWP30P140LVT U268 ( .I(n1923), .ZN(n74) );
  MAOI22D1BWP30P140LVT U269 ( .A1(i_data_bus[36]), .A2(n1914), .B1(n52), .B2(
        n75), .ZN(n1380) );
  INVD1BWP30P140LVT U270 ( .I(i_data_bus[548]), .ZN(n52) );
  OR3D1BWP30P140LVT U271 ( .A1(n76), .A2(n5479), .A3(n1296), .Z(n75) );
  MAOI22D1BWP30P140LVT U272 ( .A1(i_data_bus[86]), .A2(n1925), .B1(n53), .B2(
        n69), .ZN(n1737) );
  INVD1BWP30P140LVT U273 ( .I(i_data_bus[598]), .ZN(n53) );
  MAOI22D1BWP30P140LVT U274 ( .A1(i_data_bus[72]), .A2(n1925), .B1(n54), .B2(
        n72), .ZN(n1463) );
  INVD1BWP30P140LVT U275 ( .I(i_data_bus[904]), .ZN(n54) );
  INVD2BWP30P140LVT U276 ( .I(n128), .ZN(n72) );
  MAOI22D1BWP30P140LVT U277 ( .A1(i_data_bus[44]), .A2(n1914), .B1(n55), .B2(
        n56), .ZN(n1543) );
  INVD1BWP30P140LVT U278 ( .I(i_data_bus[620]), .ZN(n55) );
  MAOI22D1BWP30P140LVT U279 ( .A1(i_data_bus[71]), .A2(n1925), .B1(n57), .B2(
        n74), .ZN(n1443) );
  INVD1BWP30P140LVT U280 ( .I(i_data_bus[967]), .ZN(n57) );
  NR3D0P7BWP30P140LVT U281 ( .A1(n5470), .A2(n2664), .A3(n2668), .ZN(n58) );
  NR3D0P7BWP30P140LVT U282 ( .A1(n5470), .A2(n2664), .A3(n2668), .ZN(n59) );
  ND3D2BWP30P140LVT U283 ( .A1(n360), .A2(n359), .A3(n367), .ZN(n2668) );
  IND4D1BWP30P140LVT U284 ( .A1(n61), .B1(n1793), .B2(n1792), .B3(n1791), .ZN(
        n1809) );
  AO22D1BWP30P140LVT U285 ( .A1(i_data_bus[281]), .A2(n1293), .B1(
        i_data_bus[249]), .B2(n1911), .Z(n61) );
  ND4D1BWP30P140LVT U286 ( .A1(n62), .A2(n63), .A3(n64), .A4(n1610), .ZN(
        o_data_bus[111]) );
  MAOI22D1BWP30P140LVT U287 ( .A1(i_data_bus[34]), .A2(n1914), .B1(n65), .B2(
        n74), .ZN(n1345) );
  INVD1BWP30P140LVT U288 ( .I(i_data_bus[962]), .ZN(n65) );
  MAOI22D1BWP30P140LVT U289 ( .A1(i_data_bus[75]), .A2(n1925), .B1(n93), .B2(
        n74), .ZN(n1522) );
  INVD1BWP30P140LVT U290 ( .I(i_data_bus[971]), .ZN(n93) );
  NR3D1P5BWP30P140LVT U291 ( .A1(n5490), .A2(n1285), .A3(n1299), .ZN(n1923) );
  MAOI22D1BWP30P140LVT U292 ( .A1(i_data_bus[40]), .A2(n1914), .B1(n66), .B2(
        n75), .ZN(n1462) );
  INVD1BWP30P140LVT U293 ( .I(i_data_bus[552]), .ZN(n66) );
  MAOI22D1BWP30P140LVT U294 ( .A1(i_data_bus[109]), .A2(n1936), .B1(n67), .B2(
        n72), .ZN(n1559) );
  INVD1BWP30P140LVT U295 ( .I(i_data_bus[909]), .ZN(n67) );
  MAOI22D1BWP30P140LVT U296 ( .A1(i_data_bus[112]), .A2(n1936), .B1(n68), .B2(
        n72), .ZN(n1612) );
  INVD1BWP30P140LVT U297 ( .I(i_data_bus[912]), .ZN(n68) );
  INVD1BWP30P140LVT U298 ( .I(i_cmd[147]), .ZN(n70) );
  MAOI22D1BWP30P140LVT U299 ( .A1(i_data_bus[41]), .A2(n1914), .B1(n71), .B2(
        n72), .ZN(n1475) );
  INVD1BWP30P140LVT U300 ( .I(i_data_bus[905]), .ZN(n71) );
  MAOI22D1BWP30P140LVT U301 ( .A1(i_data_bus[68]), .A2(n1925), .B1(n73), .B2(
        n74), .ZN(n1378) );
  INVD1BWP30P140LVT U302 ( .I(i_data_bus[964]), .ZN(n73) );
  INVD1BWP30P140LVT U303 ( .I(i_cmd[139]), .ZN(n76) );
  INVD1BWP30P140LVT U304 ( .I(n3043), .ZN(n90) );
  MAOI22D1BWP30P140LVT U305 ( .A1(i_data_bus[87]), .A2(n1925), .B1(n77), .B2(
        n78), .ZN(n1752) );
  INVD1BWP30P140LVT U306 ( .I(i_data_bus[1015]), .ZN(n77) );
  INVD1BWP30P140LVT U307 ( .I(n1934), .ZN(n78) );
  MAOI22D1BWP30P140LVT U308 ( .A1(i_data_bus[82]), .A2(n1925), .B1(n79), .B2(
        n80), .ZN(n1652) );
  INVD1BWP30P140LVT U309 ( .I(i_data_bus[530]), .ZN(n79) );
  CKAN2D1BWP30P140LVT U310 ( .A1(n462), .A2(i_en), .Z(n82) );
  INVD1BWP30P140LVT U311 ( .I(n3307), .ZN(n112) );
  AOI22D1BWP30P140LVT U312 ( .A1(i_data_bus[306]), .A2(n3322), .B1(
        i_data_bus[786]), .B2(n3307), .ZN(n3043) );
  MAOI22D1BWP30P140LVT U313 ( .A1(i_data_bus[849]), .A2(n3316), .B1(n83), .B2(
        n84), .ZN(n3019) );
  INVD1BWP30P140LVT U314 ( .I(i_data_bus[49]), .ZN(n83) );
  INVD1BWP30P140LVT U315 ( .I(n3305), .ZN(n84) );
  MAOI22D1BWP30P140LVT U316 ( .A1(i_data_bus[837]), .A2(n3316), .B1(n85), .B2(
        n101), .ZN(n2778) );
  INVD1BWP30P140LVT U317 ( .I(i_data_bus[677]), .ZN(n85) );
  INVD1BWP30P140LVT U318 ( .I(n2653), .ZN(n101) );
  MAOI22D1BWP30P140LVT U319 ( .A1(i_data_bus[845]), .A2(n3316), .B1(n87), .B2(
        n88), .ZN(n2943) );
  INVD1BWP30P140LVT U320 ( .I(i_data_bus[269]), .ZN(n87) );
  INVD1BWP30P140LVT U321 ( .I(n3318), .ZN(n88) );
  MAOI22D1BWP30P140LVT U322 ( .A1(i_data_bus[863]), .A2(n3316), .B1(n89), .B2(
        n92), .ZN(n3326) );
  INVD1BWP30P140LVT U323 ( .I(i_data_bus[95]), .ZN(n89) );
  INVD1BWP30P140LVT U324 ( .I(n3317), .ZN(n92) );
  IND4D1BWP30P140LVT U325 ( .A1(n90), .B1(n3042), .B2(n3041), .B3(n3040), .ZN(
        n3051) );
  MAOI22D1BWP30P140LVT U326 ( .A1(i_data_bus[844]), .A2(n3316), .B1(n91), .B2(
        n92), .ZN(n2917) );
  INVD1BWP30P140LVT U327 ( .I(i_data_bus[76]), .ZN(n91) );
  MAOI22D1BWP30P140LVT U328 ( .A1(i_data_bus[843]), .A2(n3316), .B1(n93), .B2(
        n26), .ZN(n2901) );
  MAOI22D1BWP30P140LVT U329 ( .A1(i_data_bus[854]), .A2(n3316), .B1(n94), .B2(
        n101), .ZN(n3123) );
  INVD1BWP30P140LVT U330 ( .I(i_data_bus[694]), .ZN(n94) );
  MAOI22D1BWP30P140LVT U331 ( .A1(i_data_bus[846]), .A2(n3316), .B1(n95), .B2(
        n96), .ZN(n2957) );
  INVD1BWP30P140LVT U332 ( .I(i_data_bus[814]), .ZN(n95) );
  INVD1BWP30P140LVT U333 ( .I(n3304), .ZN(n96) );
  MAOI22D1BWP30P140LVT U334 ( .A1(i_data_bus[842]), .A2(n3316), .B1(n97), .B2(
        n112), .ZN(n2876) );
  INVD1BWP30P140LVT U335 ( .I(i_data_bus[778]), .ZN(n97) );
  MAOI22D1BWP30P140LVT U336 ( .A1(i_data_bus[857]), .A2(n3316), .B1(n98), .B2(
        n99), .ZN(n3179) );
  INVD1BWP30P140LVT U337 ( .I(i_data_bus[313]), .ZN(n98) );
  INVD1BWP30P140LVT U338 ( .I(n3322), .ZN(n99) );
  MAOI22D1BWP30P140LVT U339 ( .A1(i_data_bus[836]), .A2(n3316), .B1(n100), 
        .B2(n101), .ZN(n2756) );
  INVD1BWP30P140LVT U340 ( .I(i_data_bus[676]), .ZN(n100) );
  IND4D1BWP30P140LVT U341 ( .A1(n102), .B1(n3055), .B2(n3054), .B3(n3053), 
        .ZN(o_data_bus[178]) );
  INVD1BWP30P140LVT U342 ( .I(n3056), .ZN(n102) );
  MAOI22D1BWP30P140LVT U343 ( .A1(i_data_bus[859]), .A2(n3316), .B1(n3939), 
        .B2(n104), .ZN(n3218) );
  INVD1BWP30P140LVT U344 ( .I(n3321), .ZN(n104) );
  MAOI22D1BWP30P140LVT U345 ( .A1(i_data_bus[833]), .A2(n3316), .B1(n105), 
        .B2(n26), .ZN(n2695) );
  INVD1BWP30P140LVT U346 ( .I(i_data_bus[961]), .ZN(n105) );
  MAOI22D1BWP30P140LVT U347 ( .A1(i_data_bus[848]), .A2(n3316), .B1(n106), 
        .B2(n112), .ZN(n3001) );
  INVD1BWP30P140LVT U348 ( .I(i_data_bus[784]), .ZN(n106) );
  MAOI22D1BWP30P140LVT U349 ( .A1(i_data_bus[856]), .A2(n3316), .B1(n107), 
        .B2(n108), .ZN(n3158) );
  INVD1BWP30P140LVT U350 ( .I(i_data_bus[1016]), .ZN(n107) );
  INVD1BWP30P140LVT U351 ( .I(n58), .ZN(n108) );
  MAOI22D1BWP30P140LVT U352 ( .A1(i_data_bus[835]), .A2(n3316), .B1(n109), 
        .B2(n110), .ZN(n2735) );
  INVD1BWP30P140LVT U353 ( .I(i_data_bus[99]), .ZN(n109) );
  INVD1BWP30P140LVT U354 ( .I(n3308), .ZN(n110) );
  MAOI22D1BWP30P140LVT U355 ( .A1(i_data_bus[841]), .A2(n3316), .B1(n111), 
        .B2(n112), .ZN(n2859) );
  INVD1BWP30P140LVT U356 ( .I(i_data_bus[777]), .ZN(n111) );
  INVD1BWP30P140LVT U357 ( .I(i_cmd[221]), .ZN(n114) );
  MAOI22D1BWP30P140LVT U358 ( .A1(i_data_bus[855]), .A2(n3316), .B1(n115), 
        .B2(n116), .ZN(n3142) );
  INVD1BWP30P140LVT U359 ( .I(i_data_bus[759]), .ZN(n115) );
  INVD1BWP30P140LVT U360 ( .I(n2659), .ZN(n116) );
  NR2OPTPAD1BWP30P140LVT U361 ( .A1(n427), .A2(n412), .ZN(n402) );
  INR3D2BWP30P140LVT U362 ( .A1(i_cmd[218]), .B1(n5457), .B2(n3363), .ZN(n4039) );
  INR3D2BWP30P140LVT U363 ( .A1(i_cmd[210]), .B1(n5461), .B2(n3363), .ZN(n4036) );
  NR2D4BWP30P140LVT U364 ( .A1(n561), .A2(n547), .ZN(n546) );
  INVD15BWP30P140LVT U365 ( .I(i_en), .ZN(n547) );
  INR3D2BWP30P140LVT U366 ( .A1(i_cmd[201]), .B1(n619), .B2(n5459), .ZN(n1256)
         );
  NR2D1BWP30P140LVT U367 ( .A1(n547), .A2(n369), .ZN(n373) );
  INVD1BWP30P140LVT U368 ( .I(i_valid[16]), .ZN(n5477) );
  OR3D1BWP30P140LVT U369 ( .A1(i_cmd[176]), .A2(i_cmd[184]), .A3(i_cmd[168]), 
        .Z(n206) );
  INVD1BWP30P140LVT U370 ( .I(i_valid[12]), .ZN(n5476) );
  INVD1BWP30P140LVT U371 ( .I(i_valid[8]), .ZN(n5497) );
  INVD1BWP30P140LVT U372 ( .I(i_valid[0]), .ZN(n5450) );
  INVD1BWP30P140LVT U373 ( .I(i_valid[4]), .ZN(n5493) );
  INVD1BWP30P140LVT U374 ( .I(i_valid[24]), .ZN(n5444) );
  INVD1BWP30P140LVT U375 ( .I(i_valid[20]), .ZN(n5455) );
  ND2D1BWP30P140LVT U376 ( .A1(n124), .A2(n163), .ZN(n164) );
  ND2D1BWP30P140LVT U377 ( .A1(i_en), .A2(n209), .ZN(n181) );
  AOI21D1BWP30P140LVT U378 ( .A1(i_cmd[192]), .A2(n168), .B(n170), .ZN(n204)
         );
  NR2D1BWP30P140LVT U379 ( .A1(n190), .A2(n547), .ZN(n205) );
  NR2D1BWP30P140LVT U380 ( .A1(n547), .A2(n500), .ZN(n503) );
  ND2D1BWP30P140LVT U381 ( .A1(n143), .A2(n348), .ZN(n349) );
  ND2D1BWP30P140LVT U382 ( .A1(n148), .A2(n334), .ZN(n335) );
  ND2D1BWP30P140LVT U383 ( .A1(n144), .A2(n247), .ZN(n248) );
  ND2D1BWP30P140LVT U384 ( .A1(n145), .A2(n249), .ZN(n250) );
  IND2D1BWP30P140LVT U385 ( .A1(n284), .B1(n283), .ZN(n265) );
  ND3D2BWP30P140LVT U386 ( .A1(n512), .A2(n511), .A3(n510), .ZN(n3370) );
  INVD1BWP30P140LVT U387 ( .I(i_cmd[233]), .ZN(n540) );
  INVD1BWP30P140LVT U388 ( .I(i_cmd[228]), .ZN(n400) );
  INVD1BWP30P140LVT U389 ( .I(i_cmd[238]), .ZN(n306) );
  INVD1BWP30P140LVT U390 ( .I(i_cmd[232]), .ZN(n166) );
  INVD1BWP30P140LVT U391 ( .I(n3370), .ZN(n3373) );
  INVD1BWP30P140LVT U392 ( .I(i_valid[19]), .ZN(n5478) );
  INVD1BWP30P140LVT U393 ( .I(i_valid[18]), .ZN(n5481) );
  INVD1BWP30P140LVT U394 ( .I(i_valid[17]), .ZN(n5479) );
  ND2D1BWP30P140LVT U395 ( .A1(n181), .A2(n208), .ZN(n184) );
  OR3D1BWP30P140LVT U396 ( .A1(i_cmd[80]), .A2(i_cmd[88]), .A3(i_cmd[72]), .Z(
        n224) );
  ND2D1BWP30P140LVT U397 ( .A1(n133), .A2(n443), .ZN(n444) );
  ND2D1BWP30P140LVT U398 ( .A1(n125), .A2(n381), .ZN(n382) );
  IND2D1BWP30P140LVT U399 ( .A1(n423), .B1(n404), .ZN(n407) );
  ND2D1BWP30P140LVT U400 ( .A1(n402), .A2(n401), .ZN(n406) );
  ND2OPTIBD1BWP30P140LVT U401 ( .A1(n408), .A2(n409), .ZN(n403) );
  ND2OPTIBD1BWP30P140LVT U402 ( .A1(n323), .A2(n310), .ZN(n314) );
  MUX2D0BWP30P140LVT U403 ( .I0(n258), .I1(n146), .S(i_cmd[231]), .Z(n261) );
  ND2D1BWP30P140LVT U404 ( .A1(n146), .A2(n257), .ZN(n258) );
  INVD1BWP30P140LVT U405 ( .I(n282), .ZN(n266) );
  ND2D1BWP30P140LVT U406 ( .A1(n274), .A2(n276), .ZN(n264) );
  ND2D1BWP30P140LVT U407 ( .A1(n122), .A2(n245), .ZN(n246) );
  ND2D1BWP30P140LVT U408 ( .A1(n269), .A2(n270), .ZN(n272) );
  NR2D1BWP30P140LVT U409 ( .A1(n263), .A2(n262), .ZN(n271) );
  INVD1BWP30P140LVT U410 ( .I(i_valid[14]), .ZN(n4083) );
  INVD1BWP30P140LVT U411 ( .I(i_valid[13]), .ZN(n4085) );
  INVD1BWP30P140LVT U412 ( .I(i_valid[15]), .ZN(n4110) );
  CKBD1BWP30P140LVT U413 ( .I(n605), .Z(n1255) );
  NR3D1P5BWP30P140LVT U414 ( .A1(n608), .A2(n5), .A3(n5493), .ZN(n1263) );
  NR3D0P7BWP30P140LVT U415 ( .A1(n121), .A2(n590), .A3(n5450), .ZN(n1235) );
  NR3D0P7BWP30P140LVT U416 ( .A1(n593), .A2(n592), .A3(n5473), .ZN(n594) );
  NR3D0P7BWP30P140LVT U417 ( .A1(n591), .A2(n10), .A3(n5490), .ZN(n1231) );
  NR3D0P7BWP30P140LVT U418 ( .A1(n5470), .A2(n581), .A3(n10), .ZN(n1230) );
  NR3OPTPAD2BWP30P140LVT U419 ( .A1(n621), .A2(n620), .A3(n5497), .ZN(n1246)
         );
  NR3D0P7BWP30P140LVT U420 ( .A1(n585), .A2(n592), .A3(n5486), .ZN(n1242) );
  INR3D0BWP30P140LVT U421 ( .A1(i_cmd[25]), .B1(n590), .B2(n5446), .ZN(n1243)
         );
  CKBD1BWP30P140LVT U422 ( .I(n3376), .Z(n4051) );
  CKBD1BWP30P140LVT U423 ( .I(n3350), .Z(n4040) );
  NR3D0P7BWP30P140LVT U424 ( .A1(n5450), .A2(n138), .A3(n1298), .ZN(n1278) );
  NR3D0P7BWP30P140LVT U425 ( .A1(n5473), .A2(n1297), .A3(n1299), .ZN(n128) );
  NR3D0P7BWP30P140LVT U426 ( .A1(n5486), .A2(n1300), .A3(n1299), .ZN(n127) );
  AN3D1BWP30P140LVT U427 ( .A1(i_valid[7]), .A2(i_cmd[59]), .A3(n1294), .Z(
        n1911) );
  AN3D1BWP30P140LVT U428 ( .A1(i_valid[5]), .A2(i_cmd[43]), .A3(n1294), .Z(
        n1915) );
  AN3D1BWP30P140LVT U429 ( .A1(i_valid[6]), .A2(i_cmd[51]), .A3(n1294), .Z(
        n1916) );
  AN3D1BWP30P140LVT U430 ( .A1(i_cmd[12]), .A2(i_valid[1]), .A3(n1976), .Z(
        n2628) );
  AN3D1BWP30P140LVT U431 ( .A1(i_cmd[28]), .A2(i_valid[3]), .A3(n1976), .Z(
        n2623) );
  INVD1BWP30P140LVT U432 ( .I(n1976), .ZN(n1969) );
  CKBD1BWP30P140LVT U433 ( .I(n1964), .Z(n2606) );
  AN3D1BWP30P140LVT U434 ( .A1(i_cmd[20]), .A2(i_valid[2]), .A3(n1976), .Z(
        n2602) );
  CKBD1BWP30P140LVT U435 ( .I(n1965), .Z(n2614) );
  INVD1BWP30P140LVT U436 ( .I(i_valid[9]), .ZN(n4095) );
  INVD1BWP30P140LVT U437 ( .I(i_valid[11]), .ZN(n4074) );
  INVD1BWP30P140LVT U438 ( .I(i_valid[10]), .ZN(n4084) );
  ND3D1BWP30P140LVT U439 ( .A1(i_valid[15]), .A2(i_cmd[125]), .A3(n2680), .ZN(
        n3267) );
  INVD1BWP30P140LVT U440 ( .I(n2679), .ZN(n3288) );
  CKBD1BWP30P140LVT U441 ( .I(n4082), .Z(n4731) );
  INVD1BWP30P140LVT U442 ( .I(i_valid[28]), .ZN(n5473) );
  INVD1BWP30P140LVT U443 ( .I(i_valid[6]), .ZN(n5494) );
  INVD1BWP30P140LVT U444 ( .I(i_valid[5]), .ZN(n5487) );
  INVD1BWP30P140LVT U445 ( .I(i_valid[27]), .ZN(n5457) );
  INVD1BWP30P140LVT U446 ( .I(i_valid[22]), .ZN(n5448) );
  INVD1BWP30P140LVT U447 ( .I(i_valid[31]), .ZN(n5470) );
  INVD1BWP30P140LVT U448 ( .I(i_valid[26]), .ZN(n5461) );
  INVD1BWP30P140LVT U449 ( .I(i_valid[25]), .ZN(n5459) );
  INVD1BWP30P140LVT U450 ( .I(i_valid[3]), .ZN(n5446) );
  INVD1BWP30P140LVT U451 ( .I(i_valid[2]), .ZN(n5451) );
  INVD1BWP30P140LVT U452 ( .I(i_valid[29]), .ZN(n5486) );
  INVD1BWP30P140LVT U453 ( .I(i_valid[30]), .ZN(n5490) );
  INVD1BWP30P140LVT U454 ( .I(i_valid[7]), .ZN(n5471) );
  INVD1BWP30P140LVT U455 ( .I(i_valid[1]), .ZN(n5442) );
  INVD1BWP30P140LVT U456 ( .I(i_valid[23]), .ZN(n5458) );
  INVD1BWP30P140LVT U457 ( .I(i_valid[21]), .ZN(n5463) );
  ND2D1BWP30P140LVT U458 ( .A1(n160), .A2(n161), .ZN(n162) );
  ND2D1BWP30P140LVT U459 ( .A1(i_en), .A2(n180), .ZN(n208) );
  ND2D1BWP30P140LVT U460 ( .A1(n123), .A2(n173), .ZN(n174) );
  NR2D1BWP30P140LVT U461 ( .A1(n220), .A2(n547), .ZN(n193) );
  NR2D1BWP30P140LVT U462 ( .A1(n191), .A2(n205), .ZN(n185) );
  NR2D1BWP30P140LVT U463 ( .A1(n189), .A2(n547), .ZN(n186) );
  NR2D1BWP30P140LVT U464 ( .A1(n184), .A2(n213), .ZN(n192) );
  NR2D1BWP30P140LVT U465 ( .A1(n194), .A2(n547), .ZN(n219) );
  NR2D1BWP30P140LVT U466 ( .A1(n550), .A2(n547), .ZN(n553) );
  NR2D1BWP30P140LVT U467 ( .A1(n552), .A2(n547), .ZN(n549) );
  INR2D1BWP30P140LVT U468 ( .A1(n556), .B1(n559), .ZN(n554) );
  MUX2D0BWP30P140LVT U469 ( .I0(n533), .I1(n153), .S(i_cmd[33]), .Z(n557) );
  ND2D1BWP30P140LVT U470 ( .A1(n153), .A2(n532), .ZN(n533) );
  INR2D1BWP30P140LVT U471 ( .A1(n565), .B1(n566), .ZN(n567) );
  CKAN2D1BWP30P140LVT U472 ( .A1(n548), .A2(i_en), .Z(n566) );
  MUX2D0BWP30P140LVT U473 ( .I0(n480), .I1(n152), .S(i_cmd[194]), .Z(n504) );
  ND2D1BWP30P140LVT U474 ( .A1(n152), .A2(n479), .ZN(n480) );
  CKAN2D1BWP30P140LVT U475 ( .A1(n499), .A2(i_en), .Z(n515) );
  ND2D1BWP30P140LVT U476 ( .A1(n131), .A2(n486), .ZN(n487) );
  ND2D1BWP30P140LVT U477 ( .A1(n159), .A2(n491), .ZN(n492) );
  NR2D1BWP30P140LVT U478 ( .A1(n512), .A2(n547), .ZN(n497) );
  MUX2D0BWP30P140LVT U479 ( .I0(n482), .I1(n154), .S(i_cmd[162]), .Z(n500) );
  ND2D1BWP30P140LVT U480 ( .A1(n154), .A2(n481), .ZN(n482) );
  NR2D1BWP30P140LVT U481 ( .A1(n496), .A2(n547), .ZN(n511) );
  INR2D2BWP30P140LVT U482 ( .A1(n508), .B1(n519), .ZN(n510) );
  MUX2D0BWP30P140LVT U483 ( .I0(n437), .I1(n150), .S(i_cmd[163]), .Z(n468) );
  ND2D1BWP30P140LVT U484 ( .A1(n150), .A2(n436), .ZN(n437) );
  MUX2D0BWP30P140LVT U485 ( .I0(n439), .I1(n151), .S(i_cmd[195]), .Z(n464) );
  ND2D1BWP30P140LVT U486 ( .A1(n151), .A2(n438), .ZN(n439) );
  NR2D1BWP30P140LVT U487 ( .A1(n448), .A2(n547), .ZN(n472) );
  NR2D1BWP30P140LVT U488 ( .A1(n456), .A2(n547), .ZN(n475) );
  NR2D1BWP30P140LVT U489 ( .A1(n416), .A2(n547), .ZN(n419) );
  NR2D1BWP30P140LVT U490 ( .A1(n420), .A2(n547), .ZN(n417) );
  NR2D1BWP30P140LVT U491 ( .A1(n417), .A2(n419), .ZN(n408) );
  NR2D1BWP30P140LVT U492 ( .A1(n413), .A2(n547), .ZN(n427) );
  ND2D1BWP30P140LVT U493 ( .A1(n158), .A2(n390), .ZN(n391) );
  ND2D1BWP30P140LVT U494 ( .A1(i_en), .A2(n410), .ZN(n401) );
  NR2D1BWP30P140LVT U495 ( .A1(n407), .A2(n403), .ZN(n411) );
  ND2D1BWP30P140LVT U496 ( .A1(n156), .A2(n388), .ZN(n389) );
  NR2D1BWP30P140LVT U497 ( .A1(n406), .A2(n403), .ZN(n422) );
  AOI21D1BWP30P140LVT U498 ( .A1(i_cmd[5]), .A2(n136), .B(n342), .ZN(n376) );
  ND2OPTIBD1BWP30P140LVT U499 ( .A1(n353), .A2(n361), .ZN(n374) );
  AOI211OPTREPBD2BWP30P140LVT U500 ( .A1(n345), .A2(n2681), .B(n344), .C(n547), 
        .ZN(n379) );
  ND2D1BWP30P140LVT U501 ( .A1(n155), .A2(n350), .ZN(n351) );
  ND2D1BWP30P140LVT U502 ( .A1(n157), .A2(n346), .ZN(n347) );
  ND2D1BWP30P140LVT U503 ( .A1(i_en), .A2(n365), .ZN(n353) );
  CKAN2D1BWP30P140LVT U504 ( .A1(n309), .A2(i_en), .Z(n328) );
  AOI21D1BWP30P140LVT U505 ( .A1(i_cmd[6]), .A2(n134), .B(n303), .ZN(n329) );
  NR2D1BWP30P140LVT U506 ( .A1(n313), .A2(n547), .ZN(n332) );
  MUX2D0BWP30P140LVT U507 ( .I0(n296), .I1(n132), .S(i_cmd[102]), .Z(n311) );
  ND2D1BWP30P140LVT U508 ( .A1(n132), .A2(n295), .ZN(n296) );
  NR2D1BWP30P140LVT U509 ( .A1(n319), .A2(n314), .ZN(n330) );
  NR2D1BWP30P140LVT U510 ( .A1(n307), .A2(n547), .ZN(n321) );
  NR2D1BWP30P140LVT U511 ( .A1(n322), .A2(n547), .ZN(n308) );
  MUX2D0BWP30P140LVT U512 ( .I0(n294), .I1(n147), .S(i_cmd[70]), .Z(n316) );
  ND2D1BWP30P140LVT U513 ( .A1(n147), .A2(n293), .ZN(n294) );
  NR2D1BWP30P140LVT U514 ( .A1(n312), .A2(n315), .ZN(n331) );
  NR2D1BWP30P140LVT U515 ( .A1(n317), .A2(n547), .ZN(n319) );
  NR2D1BWP30P140LVT U516 ( .A1(n332), .A2(n314), .ZN(n318) );
  INR2D1BWP30P140LVT U517 ( .A1(n327), .B1(n328), .ZN(n323) );
  INVD1BWP30P140LVT U518 ( .I(n310), .ZN(n324) );
  MUX2D0BWP30P140LVT U519 ( .I0(n242), .I1(n135), .S(i_cmd[71]), .Z(n259) );
  ND2D1BWP30P140LVT U520 ( .A1(n135), .A2(n241), .ZN(n242) );
  NR2D1BWP30P140LVT U521 ( .A1(n264), .A2(n272), .ZN(n260) );
  ND2D1BWP30P140LVT U522 ( .A1(i_en), .A2(n266), .ZN(n270) );
  ND2D1BWP30P140LVT U523 ( .A1(n142), .A2(n243), .ZN(n244) );
  ND2D1BWP30P140LVT U524 ( .A1(i_en), .A2(n273), .ZN(n276) );
  IND2D1BWP30P140LVT U525 ( .A1(n272), .B1(n271), .ZN(n275) );
  INVD1BWP30P140LVT U526 ( .I(n4911), .ZN(n5423) );
  AN3D1BWP30P140LVT U527 ( .A1(i_valid[22]), .A2(i_cmd[176]), .A3(n576), .Z(
        n5424) );
  INVD1BWP30P140LVT U528 ( .I(n5220), .ZN(n5422) );
  AN3D1BWP30P140LVT U529 ( .A1(i_valid[20]), .A2(n207), .A3(n576), .Z(n5426)
         );
  AN3D1BWP30P140LVT U530 ( .A1(i_valid[23]), .A2(i_cmd[184]), .A3(n576), .Z(
        n5412) );
  INVD1BWP30P140LVT U531 ( .I(n5351), .ZN(n5394) );
  AN3D1BWP30P140LVT U532 ( .A1(i_valid[21]), .A2(i_cmd[168]), .A3(n576), .Z(
        n5393) );
  INVD1BWP30P140LVT U533 ( .I(n3327), .ZN(n2678) );
  AN3D1BWP30P140LVT U534 ( .A1(i_cmd[61]), .A2(i_valid[7]), .A3(n2677), .Z(
        n3328) );
  INVD1BWP30P140LVT U535 ( .I(n3125), .ZN(n2676) );
  CKBD1BWP30P140LVT U536 ( .I(n2658), .Z(n3302) );
  INVD1BWP30P140LVT U537 ( .I(n119), .ZN(n6192) );
  INVD1BWP30P140LVT U538 ( .I(n6116), .ZN(n6188) );
  INVD1BWP30P140LVT U539 ( .I(n5920), .ZN(n6193) );
  INVD1BWP30P140LVT U540 ( .I(n5898), .ZN(n6174) );
  CKBD1BWP30P140LVT U541 ( .I(n5445), .Z(n6165) );
  INVD1BWP30P140LVT U542 ( .I(n6094), .ZN(n6178) );
  INVD1BWP30P140LVT U543 ( .I(n5728), .ZN(n6187) );
  CKBD1BWP30P140LVT U544 ( .I(n5456), .Z(n6156) );
  AN3D1BWP30P140LVT U545 ( .A1(n194), .A2(n218), .A3(n193), .Z(n577) );
  AN3D1BWP30P140LVT U546 ( .A1(n496), .A2(n510), .A3(n497), .Z(n3371) );
  ND3D1BWP30P140LVT U547 ( .A1(n475), .A2(n474), .A3(n473), .ZN(n1296) );
  INR3D0BWP30P140LVT U548 ( .A1(n422), .B1(n405), .B2(n404), .ZN(n1976) );
  INVD1BWP30P140LVT U549 ( .I(n5496), .ZN(n5468) );
  INVD1BWP30P140LVT U550 ( .I(n5492), .ZN(n5475) );
  AN4D0BWP30P140LVT U551 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .Z(
        n3394) );
  AN4D0BWP30P140LVT U552 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .Z(
        n3414) );
  AN4D0BWP30P140LVT U553 ( .A1(n3420), .A2(n3419), .A3(n3418), .A4(n3417), .Z(
        n3435) );
  AN4D0BWP30P140LVT U554 ( .A1(n3441), .A2(n3440), .A3(n3439), .A4(n3438), .Z(
        n3457) );
  AN4D0BWP30P140LVT U555 ( .A1(n3463), .A2(n3462), .A3(n3461), .A4(n3460), .Z(
        n3478) );
  AN4D0BWP30P140LVT U556 ( .A1(n3481), .A2(n3483), .A3(n3482), .A4(n3484), .Z(
        n3498) );
  AN4D0BWP30P140LVT U557 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .Z(
        n3518) );
  AN4D0BWP30P140LVT U558 ( .A1(n3524), .A2(n3523), .A3(n3522), .A4(n3521), .Z(
        n3539) );
  AN4D0BWP30P140LVT U559 ( .A1(n3545), .A2(n3544), .A3(n3543), .A4(n3542), .Z(
        n3559) );
  AN4D0BWP30P140LVT U560 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .Z(
        n3580) );
  AN4D0BWP30P140LVT U561 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .Z(
        n3600) );
  AN4D0BWP30P140LVT U562 ( .A1(n3606), .A2(n3605), .A3(n3604), .A4(n3603), .Z(
        n3620) );
  AN4D0BWP30P140LVT U563 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .Z(
        n3640) );
  AN4D0BWP30P140LVT U564 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .Z(
        n3660) );
  AN4D0BWP30P140LVT U565 ( .A1(n3666), .A2(n3665), .A3(n3664), .A4(n3663), .Z(
        n3681) );
  AN4D0BWP30P140LVT U566 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .Z(
        n3702) );
  AN4D0BWP30P140LVT U567 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .Z(
        n3723) );
  AN4D0BWP30P140LVT U568 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .Z(
        n3743) );
  AN4D0BWP30P140LVT U569 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .Z(
        n3763) );
  AN4D0BWP30P140LVT U570 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .Z(
        n3783) );
  AN4D0BWP30P140LVT U571 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .Z(
        n3804) );
  AN4D0BWP30P140LVT U572 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .Z(
        n3825) );
  AN4D0BWP30P140LVT U573 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .Z(
        n3845) );
  AN4D0BWP30P140LVT U574 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .Z(
        n3866) );
  AN4D0BWP30P140LVT U575 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .Z(
        n3888) );
  AN4D0BWP30P140LVT U576 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .Z(
        n3908) );
  AN4D0BWP30P140LVT U577 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .Z(
        n3928) );
  AN4D0BWP30P140LVT U578 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .Z(
        n3949) );
  AN4D0BWP30P140LVT U579 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .Z(
        n3971) );
  AN4D0BWP30P140LVT U580 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .Z(
        n3995) );
  AN4D0BWP30P140LVT U581 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .Z(
        n4017) );
  AN4D0BWP30P140LVT U582 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .Z(
        n4062) );
  NR3D1P5BWP30P140LVT U583 ( .A1(n5473), .A2(n3377), .A3(n3381), .ZN(n3378) );
  NR3D1P5BWP30P140LVT U584 ( .A1(n5493), .A2(n3354), .A3(n3365), .ZN(n3355) );
  INVD1BWP30P140LVT U585 ( .I(n120), .ZN(n6143) );
  INVD1BWP30P140LVT U586 ( .I(n5488), .ZN(n6175) );
  INVD1BWP30P140LVT U587 ( .I(n222), .ZN(n5408) );
  INR3D2BWP30P140LVT U588 ( .A1(i_cmd[112]), .B1(n574), .B2(n4083), .ZN(n222)
         );
  OR3D1BWP30P140LVT U589 ( .A1(n5476), .A2(n142), .A3(n5475), .Z(n119) );
  OR3D1BWP30P140LVT U590 ( .A1(n5497), .A2(n135), .A3(n5496), .Z(n120) );
  INR3D2BWP30P140LVT U591 ( .A1(i_cmd[189]), .B1(n5458), .B2(n2666), .ZN(n2659) );
  INR3D2BWP30P140LVT U592 ( .A1(i_cmd[214]), .B1(n5461), .B2(n4106), .ZN(n4096) );
  INR3D2BWP30P140LVT U593 ( .A1(i_cmd[173]), .B1(n5463), .B2(n2666), .ZN(n2653) );
  INR3D2BWP30P140LVT U594 ( .A1(i_cmd[178]), .B1(n5448), .B2(n3361), .ZN(n3360) );
  INR3D2BWP30P140LVT U595 ( .A1(i_cmd[206]), .B1(n5459), .B2(n4106), .ZN(n4076) );
  INR3D2BWP30P140LVT U596 ( .A1(i_cmd[174]), .B1(n5463), .B2(n4093), .ZN(n4075) );
  INR3D2BWP30P140LVT U597 ( .A1(i_cmd[58]), .B1(n5471), .B2(n3365), .ZN(n3352)
         );
  INR3D2BWP30P140LVT U598 ( .A1(i_cmd[50]), .B1(n5494), .B2(n3365), .ZN(n3351)
         );
  INR3D2BWP30P140LVT U599 ( .A1(i_cmd[186]), .B1(n5458), .B2(n3361), .ZN(n3353) );
  INR3D2BWP30P140LVT U600 ( .A1(i_cmd[190]), .B1(n5458), .B2(n4093), .ZN(n4088) );
  INR3D2BWP30P140LVT U601 ( .A1(i_cmd[126]), .B1(n4110), .B2(n4109), .ZN(n4111) );
  INVD1BWP30P140LVT U602 ( .I(n2935), .ZN(n3044) );
  INVD1BWP30P140LVT U603 ( .I(n223), .ZN(n5308) );
  INR3D2BWP30P140LVT U604 ( .A1(i_cmd[120]), .B1(n574), .B2(n4110), .ZN(n223)
         );
  INVD1BWP30P140LVT U605 ( .I(n227), .ZN(n228) );
  OR3D1BWP30P140LVT U606 ( .A1(i_cmd[25]), .A2(i_cmd[9]), .A3(i_cmd[17]), .Z(
        n121) );
  OR3D1BWP30P140LVT U607 ( .A1(i_cmd[63]), .A2(i_cmd[55]), .A3(i_cmd[47]), .Z(
        n122) );
  OR3D1BWP30P140LVT U608 ( .A1(i_cmd[48]), .A2(i_cmd[56]), .A3(i_cmd[40]), .Z(
        n123) );
  OR3D1BWP30P140LVT U609 ( .A1(i_cmd[136]), .A2(i_cmd[152]), .A3(i_cmd[144]), 
        .Z(n124) );
  OR3D1BWP30P140LVT U610 ( .A1(i_cmd[140]), .A2(i_cmd[156]), .A3(i_cmd[148]), 
        .Z(n125) );
  OR3D1BWP30P140LVT U611 ( .A1(i_cmd[209]), .A2(i_cmd[201]), .A3(i_cmd[217]), 
        .Z(n126) );
  OR3D1BWP30P140LVT U612 ( .A1(i_cmd[151]), .A2(i_cmd[143]), .A3(i_cmd[159]), 
        .Z(n129) );
  OR3D1BWP30P140LVT U613 ( .A1(i_cmd[114]), .A2(i_cmd[122]), .A3(i_cmd[106]), 
        .Z(n130) );
  OR3D1BWP30P140LVT U614 ( .A1(i_cmd[26]), .A2(i_cmd[10]), .A3(i_cmd[18]), .Z(
        n131) );
  OR3D1BWP30P140LVT U615 ( .A1(i_cmd[118]), .A2(i_cmd[126]), .A3(i_cmd[110]), 
        .Z(n132) );
  OR3D1BWP30P140LVT U616 ( .A1(i_cmd[51]), .A2(i_cmd[59]), .A3(i_cmd[43]), .Z(
        n133) );
  OR3D1BWP30P140LVT U617 ( .A1(i_cmd[30]), .A2(i_cmd[14]), .A3(i_cmd[22]), .Z(
        n134) );
  OR3D1BWP30P140LVT U618 ( .A1(i_cmd[87]), .A2(i_cmd[95]), .A3(i_cmd[79]), .Z(
        n135) );
  OR3D1BWP30P140LVT U619 ( .A1(i_cmd[29]), .A2(i_cmd[13]), .A3(i_cmd[21]), .Z(
        n136) );
  OR3D1BWP30P140LVT U620 ( .A1(i_cmd[177]), .A2(i_cmd[185]), .A3(i_cmd[169]), 
        .Z(n137) );
  OR3D1BWP30P140LVT U621 ( .A1(i_cmd[27]), .A2(i_cmd[11]), .A3(i_cmd[19]), .Z(
        n138) );
  OR3D1BWP30P140LVT U622 ( .A1(i_cmd[107]), .A2(i_cmd[115]), .A3(i_cmd[123]), 
        .Z(n139) );
  OR3D1BWP30P140LVT U623 ( .A1(i_cmd[116]), .A2(i_cmd[124]), .A3(i_cmd[108]), 
        .Z(n140) );
  OR3D1BWP30P140LVT U624 ( .A1(i_cmd[54]), .A2(i_cmd[62]), .A3(i_cmd[46]), .Z(
        n141) );
  OR3D1BWP30P140LVT U625 ( .A1(i_cmd[127]), .A2(i_cmd[111]), .A3(i_cmd[119]), 
        .Z(n142) );
  OR3D1BWP30P140LVT U626 ( .A1(i_cmd[117]), .A2(i_cmd[125]), .A3(i_cmd[109]), 
        .Z(n143) );
  OR3D1BWP30P140LVT U627 ( .A1(i_cmd[191]), .A2(i_cmd[183]), .A3(i_cmd[175]), 
        .Z(n144) );
  OR3D1BWP30P140LVT U628 ( .A1(i_cmd[223]), .A2(i_cmd[215]), .A3(i_cmd[207]), 
        .Z(n145) );
  OR3D1BWP30P140LVT U629 ( .A1(i_cmd[247]), .A2(i_cmd[239]), .A3(i_cmd[255]), 
        .Z(n146) );
  OR3D1BWP30P140LVT U630 ( .A1(i_cmd[86]), .A2(i_cmd[94]), .A3(i_cmd[78]), .Z(
        n147) );
  OR3D1BWP30P140LVT U631 ( .A1(i_cmd[181]), .A2(i_cmd[189]), .A3(i_cmd[173]), 
        .Z(n148) );
  OR3D1BWP30P140LVT U632 ( .A1(i_cmd[213]), .A2(i_cmd[205]), .A3(i_cmd[221]), 
        .Z(n149) );
  OR3D1BWP30P140LVT U633 ( .A1(i_cmd[179]), .A2(i_cmd[187]), .A3(i_cmd[171]), 
        .Z(n150) );
  OR3D1BWP30P140LVT U634 ( .A1(i_cmd[211]), .A2(i_cmd[203]), .A3(i_cmd[219]), 
        .Z(n151) );
  OR3D1BWP30P140LVT U635 ( .A1(i_cmd[210]), .A2(i_cmd[202]), .A3(i_cmd[218]), 
        .Z(n152) );
  OR3D1BWP30P140LVT U636 ( .A1(i_cmd[49]), .A2(i_cmd[57]), .A3(i_cmd[41]), .Z(
        n153) );
  OR3D1BWP30P140LVT U637 ( .A1(i_cmd[178]), .A2(i_cmd[186]), .A3(i_cmd[170]), 
        .Z(n154) );
  OR3D1BWP30P140LVT U638 ( .A1(i_cmd[85]), .A2(i_cmd[93]), .A3(i_cmd[77]), .Z(
        n155) );
  OR3D1BWP30P140LVT U639 ( .A1(i_cmd[52]), .A2(i_cmd[60]), .A3(i_cmd[44]), .Z(
        n156) );
  OR3D1BWP30P140LVT U640 ( .A1(i_cmd[53]), .A2(i_cmd[61]), .A3(i_cmd[45]), .Z(
        n157) );
  OR3D1BWP30P140LVT U641 ( .A1(i_cmd[28]), .A2(i_cmd[12]), .A3(i_cmd[20]), .Z(
        n158) );
  OR3D1BWP30P140LVT U642 ( .A1(i_cmd[50]), .A2(i_cmd[58]), .A3(i_cmd[42]), .Z(
        n159) );
  MAOI222D1BWP30P140LVT U643 ( .A(i_cmd[24]), .B(i_cmd[8]), .C(i_cmd[16]), 
        .ZN(n161) );
  MUX2NUD1BWP30P140LVT U644 ( .I0(n162), .I1(n160), .S(i_cmd[0]), .ZN(n209) );
  MAOI222D1BWP30P140LVT U645 ( .A(i_cmd[136]), .B(i_cmd[152]), .C(i_cmd[144]), 
        .ZN(n163) );
  MUX2NUD1BWP30P140LVT U646 ( .I0(n164), .I1(n124), .S(i_cmd[128]), .ZN(n180)
         );
  OR4D1BWP30P140LVT U647 ( .A1(i_cmd[224]), .A2(i_cmd[240]), .A3(i_cmd[248]), 
        .A4(n166), .Z(n198) );
  INVD1BWP30P140LVT U648 ( .I(i_cmd[248]), .ZN(n165) );
  IND4D1BWP30P140LVT U649 ( .A1(i_cmd[224]), .B1(i_cmd[240]), .B2(n165), .B3(
        n166), .ZN(n197) );
  IND4D1BWP30P140LVT U650 ( .A1(i_cmd[240]), .B1(i_cmd[224]), .B2(n165), .B3(
        n166), .ZN(n187) );
  NR2D1BWP30P140LVT U651 ( .A1(i_cmd[224]), .A2(i_cmd[240]), .ZN(n167) );
  ND3D1BWP30P140LVT U652 ( .A1(i_cmd[248]), .A2(n167), .A3(n166), .ZN(n195) );
  MAOI222D1BWP30P140LVT U653 ( .A(i_cmd[208]), .B(i_cmd[200]), .C(i_cmd[216]), 
        .ZN(n169) );
  AOI21D1BWP30P140LVT U654 ( .A1(n168), .A2(n169), .B(i_cmd[192]), .ZN(n170)
         );
  CKAN2D1BWP30P140LVT U655 ( .A1(n204), .A2(i_en), .Z(n191) );
  MAOI222D1BWP30P140LVT U656 ( .A(i_cmd[176]), .B(i_cmd[184]), .C(i_cmd[168]), 
        .ZN(n171) );
  AOI21D1BWP30P140LVT U657 ( .A1(n206), .A2(n171), .B(i_cmd[160]), .ZN(n172)
         );
  AO21D1BWP30P140LVT U658 ( .A1(i_cmd[160]), .A2(n206), .B(n172), .Z(n190) );
  MAOI222D1BWP30P140LVT U659 ( .A(i_cmd[48]), .B(i_cmd[56]), .C(i_cmd[40]), 
        .ZN(n173) );
  MUX2NUD1BWP30P140LVT U660 ( .I0(n174), .I1(n123), .S(i_cmd[32]), .ZN(n210)
         );
  INR2D1BWP30P140LVT U661 ( .A1(n210), .B1(n547), .ZN(n182) );
  MAOI222D1BWP30P140LVT U662 ( .A(i_cmd[112]), .B(i_cmd[120]), .C(i_cmd[104]), 
        .ZN(n176) );
  AOI21D1BWP30P140LVT U663 ( .A1(n175), .A2(n176), .B(i_cmd[96]), .ZN(n177) );
  AO21D1BWP30P140LVT U664 ( .A1(i_cmd[96]), .A2(n175), .B(n177), .Z(n194) );
  MAOI222D1BWP30P140LVT U665 ( .A(i_cmd[80]), .B(i_cmd[88]), .C(i_cmd[72]), 
        .ZN(n178) );
  AOI21D1BWP30P140LVT U666 ( .A1(n224), .A2(n178), .B(i_cmd[64]), .ZN(n179) );
  AO21D1BWP30P140LVT U667 ( .A1(i_cmd[64]), .A2(n224), .B(n179), .Z(n220) );
  OR4D1BWP30P140LVT U668 ( .A1(n181), .A2(n180), .A3(n213), .A4(n183), .Z(n579) );
  INR3D2BWP30P140LVT U669 ( .A1(i_cmd[8]), .B1(n5442), .B2(n579), .ZN(n5395)
         );
  ND3D1BWP30P140LVT U670 ( .A1(n192), .A2(n182), .A3(n211), .ZN(n572) );
  INR3D2BWP30P140LVT U671 ( .A1(i_cmd[56]), .B1(n5471), .B2(n572), .ZN(n5401)
         );
  AO22D1BWP30P140LVT U672 ( .A1(i_data_bus[59]), .A2(n5395), .B1(
        i_data_bus[251]), .B2(n5401), .Z(n240) );
  NR2D3BWP30P140LVT U673 ( .A1(n184), .A2(n183), .ZN(n188) );
  ND3OPTPAD2BWP30P140LVT U674 ( .A1(n186), .A2(n185), .A3(n188), .ZN(n573) );
  NR3D0P7BWP30P140LVT U675 ( .A1(n5473), .A2(n187), .A3(n573), .ZN(n5389) );
  AOI22D1BWP30P140LVT U676 ( .A1(i_data_bus[923]), .A2(n5389), .B1(
        i_data_bus[155]), .B2(n5399), .ZN(n239) );
  ND2OPTIBD1BWP30P140LVT U677 ( .A1(n189), .A2(n188), .ZN(n203) );
  IND3D1BWP30P140LVT U678 ( .A1(n203), .B1(n191), .B2(n190), .ZN(n571) );
  INR3D2BWP30P140LVT U679 ( .A1(i_cmd[200]), .B1(n5459), .B2(n571), .ZN(n5427)
         );
  INR2D1BWP30P140LVT U680 ( .A1(n192), .B1(n210), .ZN(n218) );
  ND3D1BWP30P140LVT U681 ( .A1(i_valid[9]), .A2(i_cmd[72]), .A3(n577), .ZN(
        n5264) );
  AOI22D1BWP30P140LVT U682 ( .A1(i_data_bus[827]), .A2(n5427), .B1(
        i_data_bus[315]), .B2(n5428), .ZN(n238) );
  INR3D2BWP30P140LVT U683 ( .A1(i_cmd[24]), .B1(n5446), .B2(n579), .ZN(n5402)
         );
  INR3D2BWP30P140LVT U684 ( .A1(i_cmd[40]), .B1(n5487), .B2(n572), .ZN(n5391)
         );
  AO22D1BWP30P140LVT U685 ( .A1(i_data_bus[123]), .A2(n5402), .B1(
        i_data_bus[187]), .B2(n5391), .Z(n202) );
  NR3D0P7BWP30P140LVT U686 ( .A1(n5470), .A2(n195), .A3(n573), .ZN(n5396) );
  INVD1BWP30P140LVT U687 ( .I(i_cmd[0]), .ZN(n196) );
  AOI22D1BWP30P140LVT U688 ( .A1(i_data_bus[1019]), .A2(n5396), .B1(
        i_data_bus[27]), .B2(n5398), .ZN(n201) );
  INR3D2BWP30P140LVT U689 ( .A1(i_cmd[16]), .B1(n5451), .B2(n579), .ZN(n5390)
         );
  INR3D2BWP30P140LVT U690 ( .A1(i_cmd[48]), .B1(n5494), .B2(n572), .ZN(n5400)
         );
  AOI22D1BWP30P140LVT U691 ( .A1(i_data_bus[91]), .A2(n5390), .B1(
        i_data_bus[219]), .B2(n5400), .ZN(n200) );
  NR3D0P7BWP30P140LVT U692 ( .A1(n5490), .A2(n197), .A3(n573), .ZN(n5392) );
  NR3D0P7BWP30P140LVT U693 ( .A1(n5486), .A2(n198), .A3(n573), .ZN(n5397) );
  AOI22D1BWP30P140LVT U694 ( .A1(i_data_bus[987]), .A2(n5392), .B1(
        i_data_bus[955]), .B2(n5397), .ZN(n199) );
  IND4D1BWP30P140LVT U695 ( .A1(n202), .B1(n201), .B2(n200), .B3(n199), .ZN(
        n236) );
  INVD1BWP30P140LVT U696 ( .I(i_data_bus[379]), .ZN(n3939) );
  ND3D1BWP30P140LVT U697 ( .A1(i_valid[11]), .A2(i_cmd[88]), .A3(n577), .ZN(
        n4911) );
  INR3D2BWP30P140LVT U698 ( .A1(i_cmd[216]), .B1(n5457), .B2(n571), .ZN(n5410)
         );
  MOAI22D1BWP30P140LVT U699 ( .A1(n3939), .A2(n4911), .B1(i_data_bus[891]), 
        .B2(n5410), .ZN(n235) );
  INR3D0BWP30P140LVT U700 ( .A1(n205), .B1(n204), .B2(n203), .ZN(n576) );
  INVD1BWP30P140LVT U701 ( .I(n206), .ZN(n207) );
  AOI22D1BWP30P140LVT U702 ( .A1(i_data_bus[731]), .A2(n5424), .B1(
        i_data_bus[667]), .B2(n5426), .ZN(n217) );
  ND3D1BWP30P140LVT U703 ( .A1(i_valid[10]), .A2(i_cmd[80]), .A3(n577), .ZN(
        n5220) );
  AOI22D1BWP30P140LVT U704 ( .A1(i_data_bus[763]), .A2(n5412), .B1(
        i_data_bus[347]), .B2(n5422), .ZN(n216) );
  INR4D0BWP30P140LVT U705 ( .A1(n211), .B1(n210), .B2(n209), .B3(n208), .ZN(
        n212) );
  IND2D1BWP30P140LVT U706 ( .A1(n213), .B1(n212), .ZN(n578) );
  INR3D2BWP30P140LVT U707 ( .A1(i_cmd[136]), .B1(n5479), .B2(n578), .ZN(n5417)
         );
  INR3D2BWP30P140LVT U708 ( .A1(i_cmd[152]), .B1(n5478), .B2(n578), .ZN(n5416)
         );
  AOI22D1BWP30P140LVT U709 ( .A1(i_data_bus[571]), .A2(n5417), .B1(
        i_data_bus[635]), .B2(n5416), .ZN(n215) );
  INR3D2BWP30P140LVT U710 ( .A1(i_cmd[144]), .B1(n5481), .B2(n578), .ZN(n5415)
         );
  AOI22D1BWP30P140LVT U711 ( .A1(i_data_bus[603]), .A2(n5415), .B1(
        i_data_bus[539]), .B2(n5414), .ZN(n214) );
  ND4D1BWP30P140LVT U712 ( .A1(n217), .A2(n216), .A3(n215), .A4(n214), .ZN(
        n234) );
  ND3D1BWP30P140LVT U713 ( .A1(n220), .A2(n219), .A3(n218), .ZN(n574) );
  INR3D2BWP30P140LVT U714 ( .A1(i_cmd[104]), .B1(n4085), .B2(n574), .ZN(n5413)
         );
  AOI22D1BWP30P140LVT U715 ( .A1(i_data_bus[443]), .A2(n5413), .B1(
        i_data_bus[699]), .B2(n5393), .ZN(n232) );
  INVD1BWP30P140LVT U716 ( .I(i_cmd[192]), .ZN(n221) );
  AOI22D1BWP30P140LVT U717 ( .A1(i_data_bus[795]), .A2(n5407), .B1(
        i_data_bus[475]), .B2(n222), .ZN(n231) );
  INVD1BWP30P140LVT U718 ( .I(n224), .ZN(n225) );
  ND3D1BWP30P140LVT U719 ( .A1(i_valid[8]), .A2(n225), .A3(n577), .ZN(n5351)
         );
  AOI22D1BWP30P140LVT U720 ( .A1(i_data_bus[507]), .A2(n223), .B1(
        i_data_bus[283]), .B2(n5394), .ZN(n230) );
  INVD1BWP30P140LVT U721 ( .I(i_cmd[96]), .ZN(n226) );
  NR3D0P7BWP30P140LVT U722 ( .A1(n5476), .A2(n226), .A3(n574), .ZN(n227) );
  INR3D2BWP30P140LVT U723 ( .A1(i_cmd[208]), .B1(n5461), .B2(n571), .ZN(n5425)
         );
  AOI22D1BWP30P140LVT U724 ( .A1(i_data_bus[411]), .A2(n5411), .B1(
        i_data_bus[859]), .B2(n5425), .ZN(n229) );
  ND4D1BWP30P140LVT U725 ( .A1(n232), .A2(n231), .A3(n230), .A4(n229), .ZN(
        n233) );
  NR4D0BWP30P140LVT U726 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .ZN(
        n237) );
  IND4D1BWP30P140LVT U727 ( .A1(n240), .B1(n239), .B2(n238), .B3(n237), .ZN(
        o_data_bus[27]) );
  MAOI222D1BWP30P140LVT U728 ( .A(i_cmd[87]), .B(i_cmd[95]), .C(i_cmd[79]), 
        .ZN(n241) );
  MAOI222D1BWP30P140LVT U729 ( .A(i_cmd[127]), .B(i_cmd[111]), .C(i_cmd[119]), 
        .ZN(n243) );
  MUX2NUD1BWP30P140LVT U730 ( .I0(n244), .I1(n142), .S(i_cmd[103]), .ZN(n277)
         );
  MAOI222D1BWP30P140LVT U731 ( .A(i_cmd[63]), .B(i_cmd[55]), .C(i_cmd[47]), 
        .ZN(n245) );
  MUX2NUD1BWP30P140LVT U732 ( .I0(n246), .I1(n122), .S(i_cmd[39]), .ZN(n273)
         );
  MAOI222D1BWP30P140LVT U733 ( .A(i_cmd[191]), .B(i_cmd[183]), .C(i_cmd[175]), 
        .ZN(n247) );
  MAOI222D1BWP30P140LVT U734 ( .A(i_cmd[223]), .B(i_cmd[215]), .C(i_cmd[207]), 
        .ZN(n249) );
  MAOI222D1BWP30P140LVT U735 ( .A(i_cmd[151]), .B(i_cmd[143]), .C(i_cmd[159]), 
        .ZN(n251) );
  AOI21D1BWP30P140LVT U736 ( .A1(n251), .A2(n129), .B(i_cmd[135]), .ZN(n252)
         );
  AOI211D1BWP30P140LVT U737 ( .A1(i_cmd[135]), .A2(n129), .B(n547), .C(n252), 
        .ZN(n284) );
  INVD1BWP30P140LVT U738 ( .I(i_cmd[7]), .ZN(n5449) );
  NR2D1BWP30P140LVT U739 ( .A1(i_cmd[31]), .A2(n5449), .ZN(n256) );
  INVD1BWP30P140LVT U740 ( .I(i_cmd[31]), .ZN(n5447) );
  NR2D1BWP30P140LVT U741 ( .A1(i_cmd[7]), .A2(n5447), .ZN(n255) );
  INVD1BWP30P140LVT U742 ( .I(i_cmd[15]), .ZN(n5441) );
  INVD1BWP30P140LVT U743 ( .I(i_cmd[23]), .ZN(n5452) );
  AOI22D1BWP30P140LVT U744 ( .A1(i_cmd[23]), .A2(i_cmd[15]), .B1(n5441), .B2(
        n5452), .ZN(n254) );
  OAI22D1BWP30P140LVT U745 ( .A1(i_cmd[23]), .A2(i_cmd[15]), .B1(i_cmd[31]), 
        .B2(i_cmd[7]), .ZN(n253) );
  OAI31D1BWP30P140LVT U746 ( .A1(n256), .A2(n255), .A3(n254), .B(n253), .ZN(
        n282) );
  MAOI222D1BWP30P140LVT U747 ( .A(i_cmd[247]), .B(i_cmd[239]), .C(i_cmd[255]), 
        .ZN(n257) );
  ND3D1BWP30P140LVT U748 ( .A1(n259), .A2(n260), .A3(n262), .ZN(n5489) );
  ND3D1BWP30P140LVT U749 ( .A1(n263), .A2(n261), .A3(n260), .ZN(n5496) );
  INR2D2BWP30P140LVT U750 ( .A1(n271), .B1(n264), .ZN(n283) );
  ND3D1BWP30P140LVT U751 ( .A1(n268), .A2(n267), .A3(n279), .ZN(n5460) );
  NR3D0P7BWP30P140LVT U752 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n5492) );
  ND4D1BWP30P140LVT U753 ( .A1(n5460), .A2(n5453), .A3(n5475), .A4(n5495), 
        .ZN(n278) );
  INR3D0BWP30P140LVT U754 ( .A1(n5489), .B1(n5468), .B2(n278), .ZN(n286) );
  ND3D1BWP30P140LVT U755 ( .A1(n281), .A2(n280), .A3(n279), .ZN(n5462) );
  ND4D1BWP30P140LVT U756 ( .A1(n285), .A2(n284), .A3(n283), .A4(n282), .ZN(
        n5480) );
  ND3D1BWP30P140LVT U757 ( .A1(n286), .A2(n5462), .A3(n5480), .ZN(o_valid[7])
         );
  MAOI222D1BWP30P140LVT U758 ( .A(i_cmd[182]), .B(i_cmd[190]), .C(i_cmd[174]), 
        .ZN(n288) );
  AOI21D1BWP30P140LVT U759 ( .A1(n287), .A2(n288), .B(i_cmd[166]), .ZN(n289)
         );
  AO21D1BWP30P140LVT U760 ( .A1(i_cmd[166]), .A2(n287), .B(n289), .Z(n322) );
  MAOI222D1BWP30P140LVT U761 ( .A(i_cmd[214]), .B(i_cmd[206]), .C(i_cmd[222]), 
        .ZN(n291) );
  AOI21D1BWP30P140LVT U762 ( .A1(n290), .A2(n291), .B(i_cmd[198]), .ZN(n292)
         );
  AO21D1BWP30P140LVT U763 ( .A1(i_cmd[198]), .A2(n290), .B(n292), .Z(n307) );
  MAOI222D1BWP30P140LVT U764 ( .A(i_cmd[86]), .B(i_cmd[94]), .C(i_cmd[78]), 
        .ZN(n293) );
  NR2OPTPAD1BWP30P140LVT U765 ( .A1(n547), .A2(n316), .ZN(n312) );
  MAOI222D1BWP30P140LVT U766 ( .A(i_cmd[118]), .B(i_cmd[126]), .C(i_cmd[110]), 
        .ZN(n295) );
  NR2OPTPAD1BWP30P140LVT U767 ( .A1(n547), .A2(n311), .ZN(n315) );
  MAOI222D1BWP30P140LVT U768 ( .A(i_cmd[54]), .B(i_cmd[62]), .C(i_cmd[46]), 
        .ZN(n297) );
  AOI21D1BWP30P140LVT U769 ( .A1(n141), .A2(n297), .B(i_cmd[38]), .ZN(n298) );
  AO21D1BWP30P140LVT U770 ( .A1(i_cmd[38]), .A2(n141), .B(n298), .Z(n317) );
  MAOI222D1BWP30P140LVT U771 ( .A(i_cmd[142]), .B(i_cmd[158]), .C(i_cmd[150]), 
        .ZN(n300) );
  AOI21D1BWP30P140LVT U772 ( .A1(n299), .A2(n300), .B(i_cmd[134]), .ZN(n301)
         );
  AO21D1BWP30P140LVT U773 ( .A1(i_cmd[134]), .A2(n299), .B(n301), .Z(n313) );
  MAOI222D1BWP30P140LVT U774 ( .A(i_cmd[30]), .B(i_cmd[14]), .C(i_cmd[22]), 
        .ZN(n302) );
  AOI21D1BWP30P140LVT U775 ( .A1(n134), .A2(n302), .B(i_cmd[6]), .ZN(n303) );
  INVD1BWP30P140LVT U776 ( .I(i_cmd[254]), .ZN(n305) );
  IND4D1BWP30P140LVT U777 ( .A1(i_cmd[230]), .B1(i_cmd[246]), .B2(n306), .B3(
        n305), .ZN(n4067) );
  NR2D1BWP30P140LVT U778 ( .A1(i_cmd[230]), .A2(i_cmd[246]), .ZN(n304) );
  ND3D1BWP30P140LVT U779 ( .A1(i_cmd[254]), .A2(n304), .A3(n306), .ZN(n4065)
         );
  OR4D1BWP30P140LVT U780 ( .A1(i_cmd[230]), .A2(i_cmd[246]), .A3(i_cmd[254]), 
        .A4(n306), .Z(n4069) );
  IND4D1BWP30P140LVT U781 ( .A1(i_cmd[246]), .B1(i_cmd[230]), .B2(n306), .B3(
        n305), .ZN(n4072) );
  ND4D1BWP30P140LVT U782 ( .A1(n4067), .A2(n4065), .A3(n4069), .A4(n4072), 
        .ZN(n309) );
  INR3D0BWP30P140LVT U783 ( .A1(n326), .B1(n324), .B2(n309), .ZN(n320) );
  ND3D1BWP30P140LVT U784 ( .A1(n308), .A2(n307), .A3(n320), .ZN(n4093) );
  ND4D1BWP30P140LVT U785 ( .A1(n313), .A2(n312), .A3(n311), .A4(n330), .ZN(
        n4094) );
  ND4D1BWP30P140LVT U786 ( .A1(n317), .A2(n316), .A3(n315), .A4(n318), .ZN(
        n4109) );
  ND3D1BWP30P140LVT U787 ( .A1(n319), .A2(n331), .A3(n318), .ZN(n4112) );
  ND4D1BWP30P140LVT U788 ( .A1(n4093), .A2(n4094), .A3(n4109), .A4(n4112), 
        .ZN(n325) );
  ND3D1BWP30P140LVT U789 ( .A1(n322), .A2(n321), .A3(n320), .ZN(n4106) );
  ND3D1BWP30P140LVT U790 ( .A1(n326), .A2(n324), .A3(n323), .ZN(n4107) );
  IND3D1BWP30P140LVT U791 ( .A1(n325), .B1(n4106), .B2(n4107), .ZN(n333) );
  IND4D1BWP30P140LVT U792 ( .A1(n329), .B1(n328), .B2(n327), .B3(n326), .ZN(
        n4071) );
  ND3D1BWP30P140LVT U793 ( .A1(n332), .A2(n331), .A3(n330), .ZN(n4102) );
  IND3D1BWP30P140LVT U794 ( .A1(n333), .B1(n4071), .B2(n4102), .ZN(o_valid[6])
         );
  MAOI222D1BWP30P140LVT U795 ( .A(i_cmd[181]), .B(i_cmd[189]), .C(i_cmd[173]), 
        .ZN(n334) );
  MUX2D1BWP30P140LVT U796 ( .I0(n335), .I1(n148), .S(i_cmd[165]), .Z(n369) );
  MAOI222D1BWP30P140LVT U797 ( .A(i_cmd[213]), .B(i_cmd[205]), .C(i_cmd[221]), 
        .ZN(n336) );
  NR2D2BWP30P140LVT U798 ( .A1(n547), .A2(n372), .ZN(n368) );
  INVD1BWP30P140LVT U799 ( .I(i_cmd[253]), .ZN(n338) );
  INVD1BWP30P140LVT U800 ( .I(i_cmd[237]), .ZN(n340) );
  INVD1BWP30P140LVT U801 ( .I(i_cmd[229]), .ZN(n339) );
  ND4D1BWP30P140LVT U802 ( .A1(n338), .A2(n340), .A3(n339), .A4(i_cmd[245]), 
        .ZN(n2669) );
  OR4D1BWP30P140LVT U803 ( .A1(i_cmd[245]), .A2(i_cmd[229]), .A3(i_cmd[237]), 
        .A4(n338), .Z(n2664) );
  OR4D1BWP30P140LVT U804 ( .A1(i_cmd[245]), .A2(i_cmd[253]), .A3(i_cmd[237]), 
        .A4(n339), .Z(n2650) );
  OR4D1BWP30P140LVT U805 ( .A1(i_cmd[245]), .A2(i_cmd[253]), .A3(i_cmd[229]), 
        .A4(n340), .Z(n2665) );
  MAOI222D1BWP30P140LVT U806 ( .A(i_cmd[29]), .B(i_cmd[13]), .C(i_cmd[21]), 
        .ZN(n341) );
  AOI21D1BWP30P140LVT U807 ( .A1(n136), .A2(n341), .B(i_cmd[5]), .ZN(n342) );
  INR2D2BWP30P140LVT U808 ( .A1(n378), .B1(n358), .ZN(n363) );
  NR3D0P7BWP30P140LVT U809 ( .A1(i_cmd[141]), .A2(i_cmd[157]), .A3(i_cmd[149]), 
        .ZN(n345) );
  INVD1BWP30P140LVT U810 ( .I(i_cmd[133]), .ZN(n2681) );
  MAOI222D1BWP30P140LVT U811 ( .A(i_cmd[141]), .B(i_cmd[157]), .C(i_cmd[149]), 
        .ZN(n343) );
  AOI21D1BWP30P140LVT U812 ( .A1(n343), .A2(n2681), .B(n345), .ZN(n344) );
  INR2D1BWP30P140LVT U813 ( .A1(n363), .B1(n379), .ZN(n354) );
  MAOI222D1BWP30P140LVT U814 ( .A(i_cmd[53]), .B(i_cmd[61]), .C(i_cmd[45]), 
        .ZN(n346) );
  MUX2NUD1BWP30P140LVT U815 ( .I0(n347), .I1(n157), .S(i_cmd[37]), .ZN(n375)
         );
  MAOI222D1BWP30P140LVT U816 ( .A(i_cmd[117]), .B(i_cmd[125]), .C(i_cmd[109]), 
        .ZN(n348) );
  MUX2NUD1BWP30P140LVT U817 ( .I0(n349), .I1(n143), .S(i_cmd[101]), .ZN(n365)
         );
  MAOI222D1BWP30P140LVT U818 ( .A(i_cmd[85]), .B(i_cmd[93]), .C(i_cmd[77]), 
        .ZN(n350) );
  MUX2NUD1BWP30P140LVT U819 ( .I0(n351), .I1(n155), .S(i_cmd[69]), .ZN(n352)
         );
  ND3D1BWP30P140LVT U820 ( .A1(n354), .A2(n355), .A3(n356), .ZN(n2651) );
  INR4D1BWP30P140LVT U821 ( .A1(n354), .B1(n375), .B2(n353), .B3(n352), .ZN(
        n2680) );
  ND2OPTIBD2BWP30P140LVT U822 ( .A1(n356), .A2(n362), .ZN(n357) );
  IND3D1BWP30P140LVT U823 ( .A1(n357), .B1(n358), .B2(n378), .ZN(n2656) );
  INVD1BWP30P140LVT U824 ( .I(n361), .ZN(n364) );
  ND4D1BWP30P140LVT U825 ( .A1(n2656), .A2(n2668), .A3(n2667), .A4(n2670), 
        .ZN(n370) );
  NR3D0P7BWP30P140LVT U826 ( .A1(n2677), .A2(n2680), .A3(n370), .ZN(n380) );
  ND3D1BWP30P140LVT U827 ( .A1(n373), .A2(n372), .A3(n371), .ZN(n2666) );
  NR3D0P7BWP30P140LVT U828 ( .A1(n376), .A2(n375), .A3(n374), .ZN(n377) );
  ND3D1BWP30P140LVT U829 ( .A1(n379), .A2(n378), .A3(n377), .ZN(n2682) );
  ND3D1BWP30P140LVT U830 ( .A1(n380), .A2(n2666), .A3(n2682), .ZN(o_valid[5])
         );
  MAOI222D1BWP30P140LVT U831 ( .A(i_cmd[140]), .B(i_cmd[156]), .C(i_cmd[148]), 
        .ZN(n381) );
  MUX2NUD1BWP30P140LVT U832 ( .I0(n382), .I1(n125), .S(i_cmd[132]), .ZN(n410)
         );
  MAOI222D1BWP30P140LVT U833 ( .A(i_cmd[116]), .B(i_cmd[124]), .C(i_cmd[108]), 
        .ZN(n383) );
  AOI21D1BWP30P140LVT U834 ( .A1(n140), .A2(n383), .B(i_cmd[100]), .ZN(n384)
         );
  AO21D1BWP30P140LVT U835 ( .A1(i_cmd[100]), .A2(n140), .B(n384), .Z(n413) );
  MAOI222D1BWP30P140LVT U836 ( .A(i_cmd[84]), .B(i_cmd[92]), .C(i_cmd[76]), 
        .ZN(n386) );
  AOI21D1BWP30P140LVT U837 ( .A1(n385), .A2(n386), .B(i_cmd[68]), .ZN(n387) );
  AO21D1BWP30P140LVT U838 ( .A1(i_cmd[68]), .A2(n385), .B(n387), .Z(n426) );
  MAOI222D1BWP30P140LVT U839 ( .A(i_cmd[52]), .B(i_cmd[60]), .C(i_cmd[44]), 
        .ZN(n388) );
  MUX2NUD1BWP30P140LVT U840 ( .I0(n389), .I1(n156), .S(i_cmd[36]), .ZN(n405)
         );
  INR2D1BWP30P140LVT U841 ( .A1(n405), .B1(n547), .ZN(n423) );
  MAOI222D1BWP30P140LVT U842 ( .A(i_cmd[28]), .B(i_cmd[12]), .C(i_cmd[20]), 
        .ZN(n390) );
  MUX2NUD1BWP30P140LVT U843 ( .I0(n391), .I1(n158), .S(i_cmd[4]), .ZN(n424) );
  MAOI222D1BWP30P140LVT U844 ( .A(i_cmd[180]), .B(i_cmd[188]), .C(i_cmd[172]), 
        .ZN(n393) );
  AOI21D1BWP30P140LVT U845 ( .A1(n392), .A2(n393), .B(i_cmd[164]), .ZN(n394)
         );
  AO21D1BWP30P140LVT U846 ( .A1(i_cmd[164]), .A2(n392), .B(n394), .Z(n420) );
  MAOI222D1BWP30P140LVT U847 ( .A(i_cmd[212]), .B(i_cmd[204]), .C(i_cmd[220]), 
        .ZN(n396) );
  AOI21D1BWP30P140LVT U848 ( .A1(n395), .A2(n396), .B(i_cmd[196]), .ZN(n397)
         );
  AO21D1BWP30P140LVT U849 ( .A1(i_cmd[196]), .A2(n395), .B(n397), .Z(n416) );
  NR2D1BWP30P140LVT U850 ( .A1(i_cmd[252]), .A2(i_cmd[236]), .ZN(n398) );
  ND3D1BWP30P140LVT U851 ( .A1(n398), .A2(i_cmd[244]), .A3(n400), .ZN(n1957)
         );
  INVD1BWP30P140LVT U852 ( .I(i_cmd[244]), .ZN(n399) );
  IND4D1BWP30P140LVT U853 ( .A1(i_cmd[252]), .B1(i_cmd[236]), .B2(n400), .B3(
        n399), .ZN(n1968) );
  OR4D1BWP30P140LVT U854 ( .A1(i_cmd[252]), .A2(i_cmd[236]), .A3(i_cmd[244]), 
        .A4(n400), .Z(n1979) );
  IND4D1BWP30P140LVT U855 ( .A1(i_cmd[236]), .B1(i_cmd[252]), .B2(n400), .B3(
        n399), .ZN(n1967) );
  ND4D1BWP30P140LVT U856 ( .A1(n1957), .A2(n1968), .A3(n1979), .A4(n1967), 
        .ZN(n414) );
  IND3D1BWP30P140LVT U857 ( .A1(n401), .B1(n402), .B2(n411), .ZN(n1975) );
  INR2D1BWP30P140LVT U858 ( .A1(n411), .B1(n410), .ZN(n425) );
  ND3D1BWP30P140LVT U859 ( .A1(n413), .A2(n412), .A3(n425), .ZN(n1977) );
  ND3D1BWP30P140LVT U860 ( .A1(n417), .A2(n416), .A3(n418), .ZN(n1990) );
  ND4D1BWP30P140LVT U861 ( .A1(n1978), .A2(n1977), .A3(n1990), .A4(n1987), 
        .ZN(n421) );
  INR3D0BWP30P140LVT U862 ( .A1(n1975), .B1(n1976), .B2(n421), .ZN(n428) );
  IND3D1BWP30P140LVT U863 ( .A1(n424), .B1(n423), .B2(n422), .ZN(n1980) );
  ND3D1BWP30P140LVT U864 ( .A1(n427), .A2(n426), .A3(n425), .ZN(n1966) );
  ND3D1BWP30P140LVT U865 ( .A1(n428), .A2(n1980), .A3(n1966), .ZN(o_valid[4])
         );
  MAOI222D1BWP30P140LVT U866 ( .A(i_cmd[107]), .B(i_cmd[115]), .C(i_cmd[123]), 
        .ZN(n429) );
  AOI21D1BWP30P140LVT U867 ( .A1(n139), .A2(n429), .B(i_cmd[99]), .ZN(n430) );
  AO21D1BWP30P140LVT U868 ( .A1(i_cmd[99]), .A2(n139), .B(n430), .Z(n448) );
  MAOI222D1BWP30P140LVT U869 ( .A(i_cmd[139]), .B(i_cmd[155]), .C(i_cmd[147]), 
        .ZN(n432) );
  AOI21D1BWP30P140LVT U870 ( .A1(n431), .A2(n432), .B(i_cmd[131]), .ZN(n433)
         );
  AO21D1BWP30P140LVT U871 ( .A1(i_cmd[131]), .A2(n431), .B(n433), .Z(n456) );
  MAOI222D1BWP30P140LVT U872 ( .A(i_cmd[27]), .B(i_cmd[11]), .C(i_cmd[19]), 
        .ZN(n434) );
  AOI21D1BWP30P140LVT U873 ( .A1(n138), .A2(n434), .B(i_cmd[3]), .ZN(n435) );
  AO21D1BWP30P140LVT U874 ( .A1(i_cmd[3]), .A2(n138), .B(n435), .Z(n474) );
  MAOI222D1BWP30P140LVT U875 ( .A(i_cmd[179]), .B(i_cmd[187]), .C(i_cmd[171]), 
        .ZN(n436) );
  MAOI222D1BWP30P140LVT U876 ( .A(i_cmd[211]), .B(i_cmd[203]), .C(i_cmd[219]), 
        .ZN(n438) );
  INVD1BWP30P140LVT U877 ( .I(i_cmd[227]), .ZN(n441) );
  INVD1BWP30P140LVT U878 ( .I(i_cmd[243]), .ZN(n442) );
  INVD1BWP30P140LVT U879 ( .I(i_cmd[235]), .ZN(n440) );
  ND4D1BWP30P140LVT U880 ( .A1(n441), .A2(n442), .A3(n440), .A4(i_cmd[251]), 
        .ZN(n1286) );
  OR4D1BWP30P140LVT U881 ( .A1(i_cmd[251]), .A2(i_cmd[227]), .A3(i_cmd[243]), 
        .A4(n440), .Z(n1300) );
  OR4D1BWP30P140LVT U882 ( .A1(i_cmd[251]), .A2(i_cmd[235]), .A3(i_cmd[243]), 
        .A4(n441), .Z(n1297) );
  OR4D1BWP30P140LVT U883 ( .A1(i_cmd[251]), .A2(i_cmd[227]), .A3(i_cmd[235]), 
        .A4(n442), .Z(n1285) );
  ND4D1BWP30P140LVT U884 ( .A1(n1286), .A2(n1300), .A3(n1297), .A4(n1285), 
        .ZN(n462) );
  ND2OPTIBD1BWP30P140LVT U885 ( .A1(n459), .A2(n452), .ZN(n450) );
  MAOI222D1BWP30P140LVT U886 ( .A(i_cmd[51]), .B(i_cmd[59]), .C(i_cmd[43]), 
        .ZN(n443) );
  MUX2NUD1BWP30P140LVT U887 ( .I0(n444), .I1(n133), .S(i_cmd[35]), .ZN(n454)
         );
  MAOI222D1BWP30P140LVT U888 ( .A(i_cmd[83]), .B(i_cmd[91]), .C(i_cmd[75]), 
        .ZN(n446) );
  AOI21D1BWP30P140LVT U889 ( .A1(n445), .A2(n446), .B(i_cmd[67]), .ZN(n447) );
  AO21D1BWP30P140LVT U890 ( .A1(i_cmd[67]), .A2(n445), .B(n447), .Z(n471) );
  ND3D1BWP30P140LVT U891 ( .A1(n448), .A2(n470), .A3(n449), .ZN(n1295) );
  CKAN2D1BWP30P140LVT U892 ( .A1(n454), .A2(i_en), .Z(n458) );
  INR3D0BWP30P140LVT U893 ( .A1(n458), .B1(n450), .B2(n457), .ZN(n1294) );
  INR2D1BWP30P140LVT U894 ( .A1(n463), .B1(n462), .ZN(n466) );
  ND3D1BWP30P140LVT U895 ( .A1(n465), .A2(n464), .A3(n466), .ZN(n1308) );
  ND3D1BWP30P140LVT U896 ( .A1(n468), .A2(n467), .A3(n466), .ZN(n1306) );
  ND4D1BWP30P140LVT U897 ( .A1(n1298), .A2(n1299), .A3(n1308), .A4(n1306), 
        .ZN(n469) );
  INR3D0BWP30P140LVT U898 ( .A1(n1295), .B1(n1294), .B2(n469), .ZN(n476) );
  ND3D1BWP30P140LVT U899 ( .A1(n472), .A2(n471), .A3(n470), .ZN(n1287) );
  ND3D1BWP30P140LVT U900 ( .A1(n476), .A2(n1287), .A3(n1296), .ZN(o_valid[3])
         );
  MAOI222D1BWP30P140LVT U901 ( .A(i_cmd[114]), .B(i_cmd[122]), .C(i_cmd[106]), 
        .ZN(n477) );
  AOI21D1BWP30P140LVT U902 ( .A1(n130), .A2(n477), .B(i_cmd[98]), .ZN(n478) );
  AO21D1BWP30P140LVT U903 ( .A1(i_cmd[98]), .A2(n130), .B(n478), .Z(n496) );
  MAOI222D1BWP30P140LVT U904 ( .A(i_cmd[210]), .B(i_cmd[202]), .C(i_cmd[218]), 
        .ZN(n479) );
  NR2OPTPAD1BWP30P140LVT U905 ( .A1(n547), .A2(n504), .ZN(n501) );
  MAOI222D1BWP30P140LVT U906 ( .A(i_cmd[178]), .B(i_cmd[186]), .C(i_cmd[170]), 
        .ZN(n481) );
  INVD1BWP30P140LVT U907 ( .I(i_cmd[250]), .ZN(n485) );
  INVD1BWP30P140LVT U908 ( .I(i_cmd[234]), .ZN(n484) );
  INVD1BWP30P140LVT U909 ( .I(i_cmd[242]), .ZN(n483) );
  ND4D1BWP30P140LVT U910 ( .A1(n485), .A2(n484), .A3(n483), .A4(i_cmd[226]), 
        .ZN(n3377) );
  OR4D1BWP30P140LVT U911 ( .A1(i_cmd[226]), .A2(i_cmd[250]), .A3(i_cmd[234]), 
        .A4(n483), .Z(n3374) );
  OR4D1BWP30P140LVT U912 ( .A1(i_cmd[226]), .A2(i_cmd[250]), .A3(i_cmd[242]), 
        .A4(n484), .Z(n3375) );
  OR4D1BWP30P140LVT U913 ( .A1(i_cmd[226]), .A2(i_cmd[242]), .A3(i_cmd[234]), 
        .A4(n485), .Z(n3382) );
  ND4D1BWP30P140LVT U914 ( .A1(n3377), .A2(n3374), .A3(n3375), .A4(n3382), 
        .ZN(n499) );
  MAOI222D1BWP30P140LVT U915 ( .A(i_cmd[26]), .B(i_cmd[10]), .C(i_cmd[18]), 
        .ZN(n486) );
  MUX2NUD1BWP30P140LVT U916 ( .I0(n487), .I1(n131), .S(i_cmd[2]), .ZN(n518) );
  NR2OPTPAD1BWP30P140LVT U917 ( .A1(n547), .A2(n516), .ZN(n505) );
  NR3D0P7BWP30P140LVT U918 ( .A1(i_cmd[138]), .A2(i_cmd[154]), .A3(i_cmd[146]), 
        .ZN(n3379) );
  INVD1BWP30P140LVT U919 ( .I(i_cmd[130]), .ZN(n490) );
  MAOI222D1BWP30P140LVT U920 ( .A(i_cmd[138]), .B(i_cmd[154]), .C(i_cmd[146]), 
        .ZN(n488) );
  AOI21D1BWP30P140LVT U921 ( .A1(n488), .A2(n490), .B(n3379), .ZN(n489) );
  AOI211D1BWP30P140LVT U922 ( .A1(n3379), .A2(n490), .B(n489), .C(n547), .ZN(
        n522) );
  MAOI222D1BWP30P140LVT U923 ( .A(i_cmd[50]), .B(i_cmd[58]), .C(i_cmd[42]), 
        .ZN(n491) );
  MUX2NUD1BWP30P140LVT U924 ( .I0(n492), .I1(n159), .S(i_cmd[34]), .ZN(n519)
         );
  OR3D1BWP30P140LVT U925 ( .A1(i_cmd[82]), .A2(i_cmd[90]), .A3(i_cmd[74]), .Z(
        n495) );
  MAOI222D1BWP30P140LVT U926 ( .A(i_cmd[82]), .B(i_cmd[90]), .C(i_cmd[74]), 
        .ZN(n493) );
  AOI21D1BWP30P140LVT U927 ( .A1(n495), .A2(n493), .B(i_cmd[66]), .ZN(n494) );
  AO21D1BWP30P140LVT U928 ( .A1(i_cmd[66]), .A2(n495), .B(n494), .Z(n512) );
  INR2D1BWP30P140LVT U929 ( .A1(n519), .B1(n547), .ZN(n506) );
  IND2D1BWP30P140LVT U930 ( .A1(n505), .B1(n513), .ZN(n498) );
  ND3D1BWP30P140LVT U931 ( .A1(n504), .A2(n503), .A3(n502), .ZN(n3361) );
  ND3D1BWP30P140LVT U932 ( .A1(n508), .A2(n507), .A3(n506), .ZN(n3365) );
  ND4D1BWP30P140LVT U933 ( .A1(n3363), .A2(n3361), .A3(n3362), .A4(n3365), 
        .ZN(n509) );
  NR2D1BWP30P140LVT U934 ( .A1(n3371), .A2(n509), .ZN(n523) );
  ND4D1BWP30P140LVT U935 ( .A1(n516), .A2(n515), .A3(n514), .A4(n513), .ZN(
        n3381) );
  NR3D0P7BWP30P140LVT U936 ( .A1(n519), .A2(n518), .A3(n517), .ZN(n520) );
  ND3D1BWP30P140LVT U937 ( .A1(n522), .A2(n521), .A3(n520), .ZN(n3384) );
  ND4D1BWP30P140LVT U938 ( .A1(n523), .A2(n3370), .A3(n3381), .A4(n3384), .ZN(
        o_valid[2]) );
  NR3D0P7BWP30P140LVT U939 ( .A1(i_cmd[81]), .A2(i_cmd[73]), .A3(i_cmd[89]), 
        .ZN(n524) );
  INVD1BWP30P140LVT U940 ( .I(n524), .ZN(n527) );
  MAOI222D1BWP30P140LVT U941 ( .A(i_cmd[81]), .B(i_cmd[73]), .C(i_cmd[89]), 
        .ZN(n525) );
  AOI21D1BWP30P140LVT U942 ( .A1(n527), .A2(n525), .B(i_cmd[65]), .ZN(n526) );
  AO21D1BWP30P140LVT U943 ( .A1(i_cmd[65]), .A2(n527), .B(n526), .Z(n545) );
  NR3D0P7BWP30P140LVT U944 ( .A1(i_cmd[113]), .A2(i_cmd[121]), .A3(i_cmd[105]), 
        .ZN(n528) );
  INVD1BWP30P140LVT U945 ( .I(n528), .ZN(n531) );
  MAOI222D1BWP30P140LVT U946 ( .A(i_cmd[113]), .B(i_cmd[121]), .C(i_cmd[105]), 
        .ZN(n529) );
  AOI21D1BWP30P140LVT U947 ( .A1(n531), .A2(n529), .B(i_cmd[97]), .ZN(n530) );
  AO21D1BWP30P140LVT U948 ( .A1(i_cmd[97]), .A2(n531), .B(n530), .Z(n561) );
  MAOI222D1BWP30P140LVT U949 ( .A(i_cmd[49]), .B(i_cmd[57]), .C(i_cmd[41]), 
        .ZN(n532) );
  MAOI222D1BWP30P140LVT U950 ( .A(i_cmd[177]), .B(i_cmd[185]), .C(i_cmd[169]), 
        .ZN(n534) );
  AOI21D1BWP30P140LVT U951 ( .A1(n137), .A2(n534), .B(i_cmd[161]), .ZN(n535)
         );
  AO21D1BWP30P140LVT U952 ( .A1(i_cmd[161]), .A2(n137), .B(n535), .Z(n550) );
  MAOI222D1BWP30P140LVT U953 ( .A(i_cmd[209]), .B(i_cmd[201]), .C(i_cmd[217]), 
        .ZN(n536) );
  AOI21D1BWP30P140LVT U954 ( .A1(n126), .A2(n536), .B(i_cmd[193]), .ZN(n537)
         );
  AO21D1BWP30P140LVT U955 ( .A1(i_cmd[193]), .A2(n126), .B(n537), .Z(n552) );
  NR2D1BWP30P140LVT U956 ( .A1(i_cmd[225]), .A2(i_cmd[241]), .ZN(n538) );
  ND3D1BWP30P140LVT U957 ( .A1(n538), .A2(i_cmd[249]), .A3(n540), .ZN(n581) );
  OR4D1BWP30P140LVT U958 ( .A1(i_cmd[225]), .A2(i_cmd[241]), .A3(i_cmd[249]), 
        .A4(n540), .Z(n585) );
  INVD1BWP30P140LVT U959 ( .I(i_cmd[249]), .ZN(n539) );
  IND4D1BWP30P140LVT U960 ( .A1(i_cmd[241]), .B1(i_cmd[225]), .B2(n540), .B3(
        n539), .ZN(n593) );
  IND4D1BWP30P140LVT U961 ( .A1(i_cmd[225]), .B1(i_cmd[241]), .B2(n540), .B3(
        n539), .ZN(n591) );
  ND4D1BWP30P140LVT U962 ( .A1(n581), .A2(n585), .A3(n593), .A4(n591), .ZN(
        n548) );
  MAOI222D1BWP30P140LVT U963 ( .A(i_cmd[25]), .B(i_cmd[9]), .C(i_cmd[17]), 
        .ZN(n541) );
  AOI21D1BWP30P140LVT U964 ( .A1(n541), .A2(n121), .B(i_cmd[1]), .ZN(n542) );
  AOI211D1BWP30P140LVT U965 ( .A1(i_cmd[1]), .A2(n121), .B(n547), .C(n542), 
        .ZN(n569) );
  INR2D1BWP30P140LVT U966 ( .A1(n567), .B1(n569), .ZN(n556) );
  NR3D0P7BWP30P140LVT U967 ( .A1(i_cmd[137]), .A2(i_cmd[153]), .A3(i_cmd[145]), 
        .ZN(n582) );
  INVD1BWP30P140LVT U968 ( .I(i_cmd[129]), .ZN(n544) );
  MAOI222D1BWP30P140LVT U969 ( .A(i_cmd[137]), .B(i_cmd[153]), .C(i_cmd[145]), 
        .ZN(n543) );
  CKAN2D1BWP30P140LVT U970 ( .A1(n557), .A2(n554), .Z(n560) );
  NR2OPTPAD1BWP30P140LVT U971 ( .A1(n547), .A2(n557), .ZN(n555) );
  INR2D4BWP30P140LVT U972 ( .A1(n568), .B1(n569), .ZN(n564) );
  INR2D1BWP30P140LVT U973 ( .A1(n564), .B1(n548), .ZN(n551) );
  ND3D1BWP30P140LVT U974 ( .A1(n553), .A2(n552), .A3(n551), .ZN(n614) );
  ND4D1BWP30P140LVT U975 ( .A1(n607), .A2(n619), .A3(n614), .A4(n5), .ZN(n563)
         );
  ND4D2BWP30P140LVT U976 ( .A1(n559), .A2(n558), .A3(n557), .A4(n556), .ZN(
        n595) );
  IND3D1BWP30P140LVT U977 ( .A1(n563), .B1(n595), .B2(n620), .ZN(n570) );
  IND3D1BWP30P140LVT U978 ( .A1(n570), .B1(n10), .B2(n590), .ZN(o_valid[1]) );
  ND4D1BWP30P140LVT U979 ( .A1(n574), .A2(n573), .A3(n572), .A4(n571), .ZN(
        n575) );
  NR3D0P7BWP30P140LVT U980 ( .A1(n577), .A2(n576), .A3(n575), .ZN(n580) );
  ND3D1BWP30P140LVT U981 ( .A1(n580), .A2(n579), .A3(n578), .ZN(o_valid[0]) );
  AOI22D1BWP30P140LVT U982 ( .A1(i_data_bus[992]), .A2(n1230), .B1(
        i_data_bus[32]), .B2(n103), .ZN(n589) );
  AOI22D1BWP30P140LVT U983 ( .A1(i_data_bus[544]), .A2(n1233), .B1(
        i_data_bus[96]), .B2(n117), .ZN(n588) );
  INVD1BWP30P140LVT U984 ( .I(n582), .ZN(n583) );
  NR3D0P7BWP30P140LVT U985 ( .A1(n583), .A2(n595), .A3(n5477), .ZN(n584) );
  AOI22D1BWP30P140LVT U986 ( .A1(i_data_bus[0]), .A2(n25), .B1(i_data_bus[576]), .B2(n1234), .ZN(n586) );
  ND4D1BWP30P140LVT U987 ( .A1(n589), .A2(n588), .A3(n587), .A4(n586), .ZN(
        n629) );
  AOI22D1BWP30P140LVT U988 ( .A1(i_data_bus[64]), .A2(n1229), .B1(
        i_data_bus[960]), .B2(n1231), .ZN(n604) );
  AOI22D1BWP30P140LVT U989 ( .A1(i_data_bus[896]), .A2(n594), .B1(
        i_data_bus[608]), .B2(n1240), .ZN(n603) );
  INVD1BWP30P140LVT U990 ( .I(i_cmd[97]), .ZN(n596) );
  NR3D0P7BWP30P140LVT U991 ( .A1(n596), .A2(n5476), .A3(n607), .ZN(n597) );
  BUFFD2BWP30P140LVT U992 ( .I(n597), .Z(n1257) );
  INR3D0BWP30P140LVT U993 ( .A1(i_cmd[121]), .B1(n607), .B2(n4110), .ZN(n598)
         );
  BUFFD2BWP30P140LVT U994 ( .I(n598), .Z(n1247) );
  AOI22D1BWP30P140LVT U995 ( .A1(i_data_bus[384]), .A2(n1257), .B1(
        i_data_bus[480]), .B2(n1247), .ZN(n602) );
  INR3D0BWP30P140LVT U996 ( .A1(i_cmd[105]), .B1(n607), .B2(n4085), .ZN(n599)
         );
  BUFFD2BWP30P140LVT U997 ( .I(n599), .Z(n1245) );
  AOI22D1BWP30P140LVT U998 ( .A1(i_data_bus[416]), .A2(n1245), .B1(
        i_data_bus[832]), .B2(n600), .ZN(n601) );
  ND4D1BWP30P140LVT U999 ( .A1(n604), .A2(n603), .A3(n602), .A4(n601), .ZN(
        n628) );
  NR3D0P7BWP30P140LVT U1000 ( .A1(n137), .A2(n5455), .A3(n614), .ZN(n605) );
  INR3D0BWP30P140LVT U1001 ( .A1(i_cmd[185]), .B1(n614), .B2(n5458), .ZN(n606)
         );
  AOI22D1BWP30P140LVT U1002 ( .A1(i_data_bus[640]), .A2(n1255), .B1(
        i_data_bus[736]), .B2(n1254), .ZN(n613) );
  INR3D2BWP30P140LVT U1003 ( .A1(i_cmd[41]), .B1(n5487), .B2(n5), .ZN(n1265)
         );
  AOI22D1BWP30P140LVT U1004 ( .A1(i_data_bus[768]), .A2(n1253), .B1(
        i_data_bus[160]), .B2(n1265), .ZN(n612) );
  INR3D4BWP30P140LVT U1005 ( .A1(i_cmd[113]), .B1(n607), .B2(n4083), .ZN(n1267) );
  INVD1BWP30P140LVT U1006 ( .I(i_cmd[33]), .ZN(n608) );
  AOI22D1BWP30P140LVT U1007 ( .A1(i_data_bus[448]), .A2(n1267), .B1(
        i_data_bus[128]), .B2(n1263), .ZN(n611) );
  INR3D0BWP30P140LVT U1008 ( .A1(i_cmd[89]), .B1(n4074), .B2(n620), .ZN(n609)
         );
  BUFFD2BWP30P140LVT U1009 ( .I(n609), .Z(n1266) );
  INR3D2BWP30P140LVT U1010 ( .A1(i_cmd[177]), .B1(n614), .B2(n5448), .ZN(n1252) );
  AOI22D1BWP30P140LVT U1011 ( .A1(i_data_bus[352]), .A2(n1266), .B1(
        i_data_bus[704]), .B2(n1252), .ZN(n610) );
  ND4D1BWP30P140LVT U1012 ( .A1(n613), .A2(n612), .A3(n611), .A4(n610), .ZN(
        n627) );
  INR3D2BWP30P140LVT U1013 ( .A1(i_cmd[49]), .B1(n5), .B2(n5494), .ZN(n1258)
         );
  INR3D0BWP30P140LVT U1014 ( .A1(i_cmd[169]), .B1(n614), .B2(n5463), .ZN(n615)
         );
  AOI22D1BWP30P140LVT U1015 ( .A1(i_data_bus[192]), .A2(n1258), .B1(
        i_data_bus[672]), .B2(n1264), .ZN(n625) );
  INR3D2BWP30P140LVT U1016 ( .A1(i_cmd[57]), .B1(n5), .B2(n5471), .ZN(n1269)
         );
  AOI22D1BWP30P140LVT U1017 ( .A1(i_data_bus[224]), .A2(n1269), .B1(
        i_data_bus[864]), .B2(n617), .ZN(n624) );
  INR3D0BWP30P140LVT U1018 ( .A1(i_cmd[73]), .B1(n620), .B2(n4095), .ZN(n618)
         );
  AOI22D1BWP30P140LVT U1019 ( .A1(i_data_bus[288]), .A2(n1244), .B1(
        i_data_bus[800]), .B2(n1256), .ZN(n623) );
  INR3D4BWP30P140LVT U1020 ( .A1(i_cmd[81]), .B1(n620), .B2(n4084), .ZN(n1268)
         );
  INVD1BWP30P140LVT U1021 ( .I(i_cmd[65]), .ZN(n621) );
  AOI22D1BWP30P140LVT U1022 ( .A1(i_data_bus[320]), .A2(n1268), .B1(
        i_data_bus[256]), .B2(n1246), .ZN(n622) );
  ND4D1BWP30P140LVT U1023 ( .A1(n625), .A2(n624), .A3(n623), .A4(n622), .ZN(
        n626) );
  OR4D1BWP30P140LVT U1024 ( .A1(n629), .A2(n628), .A3(n627), .A4(n626), .Z(
        o_data_bus[32]) );
  AOI22D1BWP30P140LVT U1025 ( .A1(n117), .A2(i_data_bus[97]), .B1(n1234), .B2(
        i_data_bus[577]), .ZN(n633) );
  AOI22D1BWP30P140LVT U1026 ( .A1(n1233), .A2(i_data_bus[545]), .B1(n594), 
        .B2(i_data_bus[897]), .ZN(n632) );
  AOI22D1BWP30P140LVT U1027 ( .A1(n1230), .A2(i_data_bus[993]), .B1(n1231), 
        .B2(i_data_bus[961]), .ZN(n631) );
  AOI22D1BWP30P140LVT U1028 ( .A1(n103), .A2(i_data_bus[33]), .B1(n1242), .B2(
        i_data_bus[929]), .ZN(n630) );
  ND4D1BWP30P140LVT U1029 ( .A1(n633), .A2(n632), .A3(n631), .A4(n630), .ZN(
        n649) );
  AOI22D1BWP30P140LVT U1030 ( .A1(n1229), .A2(i_data_bus[65]), .B1(n1240), 
        .B2(i_data_bus[609]), .ZN(n637) );
  AOI22D1BWP30P140LVT U1031 ( .A1(n1241), .A2(i_data_bus[513]), .B1(n25), .B2(
        i_data_bus[1]), .ZN(n636) );
  AOI22D1BWP30P140LVT U1032 ( .A1(n1253), .A2(i_data_bus[769]), .B1(n1252), 
        .B2(i_data_bus[705]), .ZN(n635) );
  AOI22D1BWP30P140LVT U1033 ( .A1(n1257), .A2(i_data_bus[385]), .B1(n1264), 
        .B2(i_data_bus[673]), .ZN(n634) );
  ND4D1BWP30P140LVT U1034 ( .A1(n637), .A2(n636), .A3(n635), .A4(n634), .ZN(
        n648) );
  AOI22D1BWP30P140LVT U1035 ( .A1(n1255), .A2(i_data_bus[641]), .B1(n617), 
        .B2(i_data_bus[865]), .ZN(n641) );
  AOI22D1BWP30P140LVT U1036 ( .A1(n1247), .A2(i_data_bus[481]), .B1(n1256), 
        .B2(i_data_bus[801]), .ZN(n640) );
  AOI22D1BWP30P140LVT U1037 ( .A1(n1265), .A2(i_data_bus[161]), .B1(n1266), 
        .B2(i_data_bus[353]), .ZN(n639) );
  AOI22D1BWP30P140LVT U1038 ( .A1(n1269), .A2(i_data_bus[225]), .B1(n1246), 
        .B2(i_data_bus[257]), .ZN(n638) );
  ND4D1BWP30P140LVT U1039 ( .A1(n641), .A2(n640), .A3(n639), .A4(n638), .ZN(
        n647) );
  AOI22D1BWP30P140LVT U1040 ( .A1(n1267), .A2(i_data_bus[449]), .B1(n1244), 
        .B2(i_data_bus[289]), .ZN(n645) );
  AOI22D1BWP30P140LVT U1041 ( .A1(n1254), .A2(i_data_bus[737]), .B1(n1258), 
        .B2(i_data_bus[193]), .ZN(n644) );
  AOI22D1BWP30P140LVT U1042 ( .A1(n1245), .A2(i_data_bus[417]), .B1(n1263), 
        .B2(i_data_bus[129]), .ZN(n643) );
  AOI22D1BWP30P140LVT U1043 ( .A1(n600), .A2(i_data_bus[833]), .B1(n1268), 
        .B2(i_data_bus[321]), .ZN(n642) );
  ND4D1BWP30P140LVT U1044 ( .A1(n645), .A2(n644), .A3(n643), .A4(n642), .ZN(
        n646) );
  OR4D1BWP30P140LVT U1045 ( .A1(n646), .A2(n648), .A3(n647), .A4(n649), .Z(
        o_data_bus[33]) );
  AOI22D1BWP30P140LVT U1046 ( .A1(n1233), .A2(i_data_bus[546]), .B1(n1234), 
        .B2(i_data_bus[578]), .ZN(n653) );
  AOI22D1BWP30P140LVT U1047 ( .A1(n1232), .A2(i_data_bus[34]), .B1(n594), .B2(
        i_data_bus[898]), .ZN(n651) );
  AOI22D1BWP30P140LVT U1048 ( .A1(n1241), .A2(i_data_bus[514]), .B1(n25), .B2(
        i_data_bus[2]), .ZN(n650) );
  ND4D1BWP30P140LVT U1049 ( .A1(n651), .A2(n652), .A3(n653), .A4(n650), .ZN(
        n669) );
  AOI22D1BWP30P140LVT U1050 ( .A1(n1230), .A2(i_data_bus[994]), .B1(n117), 
        .B2(i_data_bus[98]), .ZN(n657) );
  AOI22D1BWP30P140LVT U1051 ( .A1(n1242), .A2(i_data_bus[930]), .B1(n1240), 
        .B2(i_data_bus[610]), .ZN(n656) );
  AOI22D1BWP30P140LVT U1052 ( .A1(n1265), .A2(i_data_bus[162]), .B1(n617), 
        .B2(i_data_bus[866]), .ZN(n655) );
  AOI22D1BWP30P140LVT U1053 ( .A1(n1258), .A2(i_data_bus[194]), .B1(n1264), 
        .B2(i_data_bus[674]), .ZN(n654) );
  ND4D1BWP30P140LVT U1054 ( .A1(n657), .A2(n656), .A3(n655), .A4(n654), .ZN(
        n668) );
  AOI22D1BWP30P140LVT U1055 ( .A1(n1247), .A2(i_data_bus[482]), .B1(n1244), 
        .B2(i_data_bus[290]), .ZN(n661) );
  AOI22D1BWP30P140LVT U1056 ( .A1(n1257), .A2(i_data_bus[386]), .B1(n1245), 
        .B2(i_data_bus[418]), .ZN(n660) );
  AOI22D1BWP30P140LVT U1057 ( .A1(n1267), .A2(i_data_bus[450]), .B1(n1256), 
        .B2(i_data_bus[802]), .ZN(n659) );
  AOI22D1BWP30P140LVT U1058 ( .A1(n1253), .A2(i_data_bus[770]), .B1(n1269), 
        .B2(i_data_bus[226]), .ZN(n658) );
  ND4D1BWP30P140LVT U1059 ( .A1(n661), .A2(n660), .A3(n659), .A4(n658), .ZN(
        n667) );
  AOI22D1BWP30P140LVT U1060 ( .A1(n600), .A2(i_data_bus[834]), .B1(n1254), 
        .B2(i_data_bus[738]), .ZN(n665) );
  AOI22D1BWP30P140LVT U1061 ( .A1(n1266), .A2(i_data_bus[354]), .B1(n1252), 
        .B2(i_data_bus[706]), .ZN(n664) );
  AOI22D1BWP30P140LVT U1062 ( .A1(n1255), .A2(i_data_bus[642]), .B1(n1263), 
        .B2(i_data_bus[130]), .ZN(n663) );
  AOI22D1BWP30P140LVT U1063 ( .A1(n1268), .A2(i_data_bus[322]), .B1(n1246), 
        .B2(i_data_bus[258]), .ZN(n662) );
  ND4D1BWP30P140LVT U1064 ( .A1(n665), .A2(n664), .A3(n663), .A4(n662), .ZN(
        n666) );
  OR4D1BWP30P140LVT U1065 ( .A1(n669), .A2(n668), .A3(n667), .A4(n666), .Z(
        o_data_bus[34]) );
  AOI22D1BWP30P140LVT U1066 ( .A1(n1234), .A2(i_data_bus[579]), .B1(n594), 
        .B2(i_data_bus[899]), .ZN(n672) );
  AOI22D1BWP30P140LVT U1067 ( .A1(n103), .A2(i_data_bus[35]), .B1(n25), .B2(
        i_data_bus[3]), .ZN(n671) );
  AOI22D1BWP30P140LVT U1068 ( .A1(n117), .A2(i_data_bus[99]), .B1(n1231), .B2(
        i_data_bus[963]), .ZN(n670) );
  AOI22D1BWP30P140LVT U1069 ( .A1(n1233), .A2(i_data_bus[547]), .B1(n1240), 
        .B2(i_data_bus[611]), .ZN(n676) );
  AOI22D1BWP30P140LVT U1070 ( .A1(n1230), .A2(i_data_bus[995]), .B1(n1242), 
        .B2(i_data_bus[931]), .ZN(n675) );
  AOI22D1BWP30P140LVT U1071 ( .A1(n1266), .A2(i_data_bus[355]), .B1(n1246), 
        .B2(i_data_bus[259]), .ZN(n674) );
  AOI22D1BWP30P140LVT U1072 ( .A1(n1257), .A2(i_data_bus[387]), .B1(n600), 
        .B2(i_data_bus[835]), .ZN(n673) );
  ND4D1BWP30P140LVT U1073 ( .A1(n676), .A2(n675), .A3(n674), .A4(n673), .ZN(
        n687) );
  AOI22D1BWP30P140LVT U1074 ( .A1(n1247), .A2(i_data_bus[483]), .B1(n1245), 
        .B2(i_data_bus[419]), .ZN(n680) );
  AOI22D1BWP30P140LVT U1075 ( .A1(n1263), .A2(i_data_bus[131]), .B1(n1268), 
        .B2(i_data_bus[323]), .ZN(n679) );
  AOI22D1BWP30P140LVT U1076 ( .A1(n1254), .A2(i_data_bus[739]), .B1(n1253), 
        .B2(i_data_bus[771]), .ZN(n678) );
  AOI22D1BWP30P140LVT U1077 ( .A1(n1265), .A2(i_data_bus[163]), .B1(n1264), 
        .B2(i_data_bus[675]), .ZN(n677) );
  ND4D1BWP30P140LVT U1078 ( .A1(n680), .A2(n679), .A3(n678), .A4(n677), .ZN(
        n686) );
  AOI22D1BWP30P140LVT U1079 ( .A1(n1255), .A2(i_data_bus[643]), .B1(n1269), 
        .B2(i_data_bus[227]), .ZN(n684) );
  AOI22D1BWP30P140LVT U1080 ( .A1(n617), .A2(i_data_bus[867]), .B1(n1244), 
        .B2(i_data_bus[291]), .ZN(n683) );
  AOI22D1BWP30P140LVT U1081 ( .A1(n1252), .A2(i_data_bus[707]), .B1(n1256), 
        .B2(i_data_bus[803]), .ZN(n682) );
  AOI22D1BWP30P140LVT U1082 ( .A1(n1267), .A2(i_data_bus[451]), .B1(n1258), 
        .B2(i_data_bus[195]), .ZN(n681) );
  ND4D1BWP30P140LVT U1083 ( .A1(n684), .A2(n683), .A3(n682), .A4(n681), .ZN(
        n685) );
  OR4D1BWP30P140LVT U1084 ( .A1(n685), .A2(n687), .A3(n686), .A4(n688), .Z(
        o_data_bus[35]) );
  AOI22D1BWP30P140LVT U1085 ( .A1(n1233), .A2(i_data_bus[548]), .B1(n117), 
        .B2(i_data_bus[100]), .ZN(n692) );
  AOI22D1BWP30P140LVT U1086 ( .A1(n1231), .A2(i_data_bus[964]), .B1(n1240), 
        .B2(i_data_bus[612]), .ZN(n691) );
  AOI22D1BWP30P140LVT U1087 ( .A1(n1242), .A2(i_data_bus[932]), .B1(n594), 
        .B2(i_data_bus[900]), .ZN(n690) );
  AOI22D1BWP30P140LVT U1088 ( .A1(n1241), .A2(i_data_bus[516]), .B1(n1229), 
        .B2(i_data_bus[68]), .ZN(n689) );
  ND4D1BWP30P140LVT U1089 ( .A1(n690), .A2(n691), .A3(n692), .A4(n689), .ZN(
        n708) );
  AOI22D1BWP30P140LVT U1090 ( .A1(n1230), .A2(i_data_bus[996]), .B1(n103), 
        .B2(i_data_bus[36]), .ZN(n696) );
  AOI22D1BWP30P140LVT U1091 ( .A1(n25), .A2(i_data_bus[4]), .B1(n1234), .B2(
        i_data_bus[580]), .ZN(n695) );
  AOI22D1BWP30P140LVT U1092 ( .A1(n1254), .A2(i_data_bus[740]), .B1(n1258), 
        .B2(i_data_bus[196]), .ZN(n694) );
  AOI22D1BWP30P140LVT U1093 ( .A1(n1253), .A2(i_data_bus[772]), .B1(n1252), 
        .B2(i_data_bus[708]), .ZN(n693) );
  ND4D1BWP30P140LVT U1094 ( .A1(n696), .A2(n695), .A3(n694), .A4(n693), .ZN(
        n707) );
  AOI22D1BWP30P140LVT U1095 ( .A1(n1263), .A2(i_data_bus[132]), .B1(n1269), 
        .B2(i_data_bus[228]), .ZN(n700) );
  AOI22D1BWP30P140LVT U1096 ( .A1(n1245), .A2(i_data_bus[420]), .B1(n1267), 
        .B2(i_data_bus[452]), .ZN(n699) );
  AOI22D1BWP30P140LVT U1097 ( .A1(n1247), .A2(i_data_bus[484]), .B1(n617), 
        .B2(i_data_bus[868]), .ZN(n698) );
  AOI22D1BWP30P140LVT U1098 ( .A1(n1265), .A2(i_data_bus[164]), .B1(n1264), 
        .B2(i_data_bus[676]), .ZN(n697) );
  ND4D1BWP30P140LVT U1099 ( .A1(n700), .A2(n699), .A3(n698), .A4(n697), .ZN(
        n706) );
  AOI22D1BWP30P140LVT U1100 ( .A1(n1244), .A2(i_data_bus[292]), .B1(n1268), 
        .B2(i_data_bus[324]), .ZN(n704) );
  AOI22D1BWP30P140LVT U1101 ( .A1(n1255), .A2(i_data_bus[644]), .B1(n1266), 
        .B2(i_data_bus[356]), .ZN(n703) );
  AOI22D1BWP30P140LVT U1102 ( .A1(n600), .A2(i_data_bus[836]), .B1(n1246), 
        .B2(i_data_bus[260]), .ZN(n702) );
  AOI22D1BWP30P140LVT U1103 ( .A1(n1257), .A2(i_data_bus[388]), .B1(n1256), 
        .B2(i_data_bus[804]), .ZN(n701) );
  ND4D1BWP30P140LVT U1104 ( .A1(n704), .A2(n703), .A3(n702), .A4(n701), .ZN(
        n705) );
  OR4D1BWP30P140LVT U1105 ( .A1(n708), .A2(n707), .A3(n706), .A4(n705), .Z(
        o_data_bus[36]) );
  AOI22D1BWP30P140LVT U1106 ( .A1(n1241), .A2(i_data_bus[517]), .B1(n594), 
        .B2(i_data_bus[901]), .ZN(n712) );
  AOI22D1BWP30P140LVT U1107 ( .A1(n1232), .A2(i_data_bus[37]), .B1(n1233), 
        .B2(i_data_bus[549]), .ZN(n711) );
  AOI22D1BWP30P140LVT U1108 ( .A1(n25), .A2(i_data_bus[5]), .B1(n1234), .B2(
        i_data_bus[581]), .ZN(n710) );
  ND4D1BWP30P140LVT U1109 ( .A1(n712), .A2(n711), .A3(n710), .A4(n709), .ZN(
        n728) );
  AOI22D1BWP30P140LVT U1110 ( .A1(n1231), .A2(i_data_bus[965]), .B1(n1240), 
        .B2(i_data_bus[613]), .ZN(n716) );
  AOI22D1BWP30P140LVT U1111 ( .A1(n1230), .A2(i_data_bus[997]), .B1(n1229), 
        .B2(i_data_bus[69]), .ZN(n715) );
  AOI22D1BWP30P140LVT U1112 ( .A1(n1253), .A2(i_data_bus[773]), .B1(n1258), 
        .B2(i_data_bus[197]), .ZN(n714) );
  AOI22D1BWP30P140LVT U1113 ( .A1(n1255), .A2(i_data_bus[645]), .B1(n1264), 
        .B2(i_data_bus[677]), .ZN(n713) );
  ND4D1BWP30P140LVT U1114 ( .A1(n716), .A2(n715), .A3(n714), .A4(n713), .ZN(
        n727) );
  AOI22D1BWP30P140LVT U1115 ( .A1(n600), .A2(i_data_bus[837]), .B1(n1256), 
        .B2(i_data_bus[805]), .ZN(n720) );
  AOI22D1BWP30P140LVT U1116 ( .A1(n1265), .A2(i_data_bus[165]), .B1(n617), 
        .B2(i_data_bus[869]), .ZN(n719) );
  AOI22D1BWP30P140LVT U1117 ( .A1(n1267), .A2(i_data_bus[453]), .B1(n1252), 
        .B2(i_data_bus[709]), .ZN(n718) );
  AOI22D1BWP30P140LVT U1118 ( .A1(n1247), .A2(i_data_bus[485]), .B1(n1266), 
        .B2(i_data_bus[357]), .ZN(n717) );
  ND4D1BWP30P140LVT U1119 ( .A1(n720), .A2(n719), .A3(n718), .A4(n717), .ZN(
        n726) );
  AOI22D1BWP30P140LVT U1120 ( .A1(n1245), .A2(i_data_bus[421]), .B1(n1244), 
        .B2(i_data_bus[293]), .ZN(n724) );
  AOI22D1BWP30P140LVT U1121 ( .A1(n1254), .A2(i_data_bus[741]), .B1(n1263), 
        .B2(i_data_bus[133]), .ZN(n723) );
  AOI22D1BWP30P140LVT U1122 ( .A1(n1268), .A2(i_data_bus[325]), .B1(n1246), 
        .B2(i_data_bus[261]), .ZN(n722) );
  AOI22D1BWP30P140LVT U1123 ( .A1(n1257), .A2(i_data_bus[389]), .B1(n1269), 
        .B2(i_data_bus[229]), .ZN(n721) );
  ND4D1BWP30P140LVT U1124 ( .A1(n724), .A2(n723), .A3(n722), .A4(n721), .ZN(
        n725) );
  OR4D1BWP30P140LVT U1125 ( .A1(n728), .A2(n727), .A3(n726), .A4(n725), .Z(
        o_data_bus[37]) );
  AOI22D1BWP30P140LVT U1126 ( .A1(n1234), .A2(i_data_bus[582]), .B1(n1231), 
        .B2(i_data_bus[966]), .ZN(n732) );
  AOI22D1BWP30P140LVT U1127 ( .A1(n1233), .A2(i_data_bus[550]), .B1(n1240), 
        .B2(i_data_bus[614]), .ZN(n731) );
  AOI22D1BWP30P140LVT U1128 ( .A1(n103), .A2(i_data_bus[38]), .B1(n1242), .B2(
        i_data_bus[934]), .ZN(n730) );
  AOI22D1BWP30P140LVT U1129 ( .A1(n25), .A2(i_data_bus[6]), .B1(n1229), .B2(
        i_data_bus[70]), .ZN(n729) );
  ND4D1BWP30P140LVT U1130 ( .A1(n732), .A2(n730), .A3(n731), .A4(n729), .ZN(
        n748) );
  AOI22D1BWP30P140LVT U1131 ( .A1(n117), .A2(i_data_bus[102]), .B1(n1241), 
        .B2(i_data_bus[518]), .ZN(n736) );
  AOI22D1BWP30P140LVT U1132 ( .A1(n1230), .A2(i_data_bus[998]), .B1(n594), 
        .B2(i_data_bus[902]), .ZN(n735) );
  AOI22D1BWP30P140LVT U1133 ( .A1(n617), .A2(i_data_bus[870]), .B1(n1256), 
        .B2(i_data_bus[806]), .ZN(n734) );
  AOI22D1BWP30P140LVT U1134 ( .A1(n1247), .A2(i_data_bus[486]), .B1(n600), 
        .B2(i_data_bus[838]), .ZN(n733) );
  ND4D1BWP30P140LVT U1135 ( .A1(n736), .A2(n735), .A3(n734), .A4(n733), .ZN(
        n747) );
  AOI22D1BWP30P140LVT U1136 ( .A1(n1254), .A2(i_data_bus[742]), .B1(n1269), 
        .B2(i_data_bus[230]), .ZN(n740) );
  AOI22D1BWP30P140LVT U1137 ( .A1(n1255), .A2(i_data_bus[646]), .B1(n1265), 
        .B2(i_data_bus[166]), .ZN(n739) );
  AOI22D1BWP30P140LVT U1138 ( .A1(n1257), .A2(i_data_bus[390]), .B1(n1267), 
        .B2(i_data_bus[454]), .ZN(n738) );
  AOI22D1BWP30P140LVT U1139 ( .A1(n1266), .A2(i_data_bus[358]), .B1(n1252), 
        .B2(i_data_bus[710]), .ZN(n737) );
  ND4D1BWP30P140LVT U1140 ( .A1(n740), .A2(n739), .A3(n738), .A4(n737), .ZN(
        n746) );
  AOI22D1BWP30P140LVT U1141 ( .A1(n1253), .A2(i_data_bus[774]), .B1(n1258), 
        .B2(i_data_bus[198]), .ZN(n744) );
  AOI22D1BWP30P140LVT U1142 ( .A1(n1245), .A2(i_data_bus[422]), .B1(n1244), 
        .B2(i_data_bus[294]), .ZN(n743) );
  AOI22D1BWP30P140LVT U1143 ( .A1(n1263), .A2(i_data_bus[134]), .B1(n1264), 
        .B2(i_data_bus[678]), .ZN(n742) );
  AOI22D1BWP30P140LVT U1144 ( .A1(n1268), .A2(i_data_bus[326]), .B1(n1246), 
        .B2(i_data_bus[262]), .ZN(n741) );
  ND4D1BWP30P140LVT U1145 ( .A1(n744), .A2(n743), .A3(n742), .A4(n741), .ZN(
        n745) );
  OR4D1BWP30P140LVT U1146 ( .A1(n748), .A2(n747), .A3(n746), .A4(n745), .Z(
        o_data_bus[38]) );
  AOI22D1BWP30P140LVT U1147 ( .A1(n1232), .A2(i_data_bus[39]), .B1(n1240), 
        .B2(i_data_bus[615]), .ZN(n752) );
  AOI22D1BWP30P140LVT U1148 ( .A1(n1233), .A2(i_data_bus[551]), .B1(n1234), 
        .B2(i_data_bus[583]), .ZN(n750) );
  ND4D1BWP30P140LVT U1149 ( .A1(n752), .A2(n751), .A3(n750), .A4(n749), .ZN(
        n768) );
  AOI22D1BWP30P140LVT U1150 ( .A1(n1230), .A2(i_data_bus[999]), .B1(n1242), 
        .B2(i_data_bus[935]), .ZN(n756) );
  AOI22D1BWP30P140LVT U1151 ( .A1(n25), .A2(i_data_bus[7]), .B1(n1229), .B2(
        i_data_bus[71]), .ZN(n755) );
  AOI22D1BWP30P140LVT U1152 ( .A1(n1267), .A2(i_data_bus[455]), .B1(n1266), 
        .B2(i_data_bus[359]), .ZN(n754) );
  AOI22D1BWP30P140LVT U1153 ( .A1(n617), .A2(i_data_bus[871]), .B1(n1246), 
        .B2(i_data_bus[263]), .ZN(n753) );
  ND4D1BWP30P140LVT U1154 ( .A1(n756), .A2(n755), .A3(n754), .A4(n753), .ZN(
        n767) );
  AOI22D1BWP30P140LVT U1155 ( .A1(n1257), .A2(i_data_bus[391]), .B1(n1264), 
        .B2(i_data_bus[679]), .ZN(n760) );
  AOI22D1BWP30P140LVT U1156 ( .A1(n1247), .A2(i_data_bus[487]), .B1(n1256), 
        .B2(i_data_bus[807]), .ZN(n759) );
  AOI22D1BWP30P140LVT U1157 ( .A1(n600), .A2(i_data_bus[839]), .B1(n1254), 
        .B2(i_data_bus[743]), .ZN(n758) );
  AOI22D1BWP30P140LVT U1158 ( .A1(n1253), .A2(i_data_bus[775]), .B1(n1252), 
        .B2(i_data_bus[711]), .ZN(n757) );
  ND4D1BWP30P140LVT U1159 ( .A1(n760), .A2(n759), .A3(n758), .A4(n757), .ZN(
        n766) );
  AOI22D1BWP30P140LVT U1160 ( .A1(n1265), .A2(i_data_bus[167]), .B1(n1263), 
        .B2(i_data_bus[135]), .ZN(n764) );
  AOI22D1BWP30P140LVT U1161 ( .A1(n1255), .A2(i_data_bus[647]), .B1(n1244), 
        .B2(i_data_bus[295]), .ZN(n763) );
  AOI22D1BWP30P140LVT U1162 ( .A1(n1245), .A2(i_data_bus[423]), .B1(n1268), 
        .B2(i_data_bus[327]), .ZN(n762) );
  AOI22D1BWP30P140LVT U1163 ( .A1(n1258), .A2(i_data_bus[199]), .B1(n1269), 
        .B2(i_data_bus[231]), .ZN(n761) );
  ND4D1BWP30P140LVT U1164 ( .A1(n764), .A2(n763), .A3(n762), .A4(n761), .ZN(
        n765) );
  OR4D1BWP30P140LVT U1165 ( .A1(n768), .A2(n767), .A3(n766), .A4(n765), .Z(
        o_data_bus[39]) );
  AOI22D1BWP30P140LVT U1166 ( .A1(n1242), .A2(i_data_bus[936]), .B1(n1240), 
        .B2(i_data_bus[616]), .ZN(n771) );
  AOI22D1BWP30P140LVT U1167 ( .A1(n1233), .A2(i_data_bus[552]), .B1(n117), 
        .B2(i_data_bus[104]), .ZN(n770) );
  AOI22D1BWP30P140LVT U1168 ( .A1(n1230), .A2(i_data_bus[1000]), .B1(n594), 
        .B2(i_data_bus[904]), .ZN(n769) );
  ND4D1BWP30P140LVT U1169 ( .A1(n769), .A2(n772), .A3(n770), .A4(n771), .ZN(
        n788) );
  AOI22D1BWP30P140LVT U1170 ( .A1(n1241), .A2(i_data_bus[520]), .B1(n1234), 
        .B2(i_data_bus[584]), .ZN(n776) );
  AOI22D1BWP30P140LVT U1171 ( .A1(n1232), .A2(i_data_bus[40]), .B1(n1229), 
        .B2(i_data_bus[72]), .ZN(n775) );
  AOI22D1BWP30P140LVT U1172 ( .A1(n1267), .A2(i_data_bus[456]), .B1(n1246), 
        .B2(i_data_bus[264]), .ZN(n774) );
  AOI22D1BWP30P140LVT U1173 ( .A1(n1245), .A2(i_data_bus[424]), .B1(n1265), 
        .B2(i_data_bus[168]), .ZN(n773) );
  ND4D1BWP30P140LVT U1174 ( .A1(n776), .A2(n775), .A3(n774), .A4(n773), .ZN(
        n787) );
  AOI22D1BWP30P140LVT U1175 ( .A1(n600), .A2(i_data_bus[840]), .B1(n1254), 
        .B2(i_data_bus[744]), .ZN(n780) );
  AOI22D1BWP30P140LVT U1176 ( .A1(n1264), .A2(i_data_bus[680]), .B1(n1268), 
        .B2(i_data_bus[328]), .ZN(n779) );
  AOI22D1BWP30P140LVT U1177 ( .A1(n1258), .A2(i_data_bus[200]), .B1(n1256), 
        .B2(i_data_bus[808]), .ZN(n778) );
  AOI22D1BWP30P140LVT U1178 ( .A1(n1247), .A2(i_data_bus[488]), .B1(n1244), 
        .B2(i_data_bus[296]), .ZN(n777) );
  ND4D1BWP30P140LVT U1179 ( .A1(n780), .A2(n779), .A3(n778), .A4(n777), .ZN(
        n786) );
  AOI22D1BWP30P140LVT U1180 ( .A1(n1252), .A2(i_data_bus[712]), .B1(n617), 
        .B2(i_data_bus[872]), .ZN(n784) );
  AOI22D1BWP30P140LVT U1181 ( .A1(n1257), .A2(i_data_bus[392]), .B1(n1266), 
        .B2(i_data_bus[360]), .ZN(n783) );
  AOI22D1BWP30P140LVT U1182 ( .A1(n1263), .A2(i_data_bus[136]), .B1(n1269), 
        .B2(i_data_bus[232]), .ZN(n782) );
  AOI22D1BWP30P140LVT U1183 ( .A1(n1255), .A2(i_data_bus[648]), .B1(n1253), 
        .B2(i_data_bus[776]), .ZN(n781) );
  ND4D1BWP30P140LVT U1184 ( .A1(n784), .A2(n783), .A3(n782), .A4(n781), .ZN(
        n785) );
  OR4D1BWP30P140LVT U1185 ( .A1(n788), .A2(n787), .A3(n786), .A4(n785), .Z(
        o_data_bus[40]) );
  AOI22D1BWP30P140LVT U1186 ( .A1(n1241), .A2(i_data_bus[521]), .B1(n25), .B2(
        i_data_bus[9]), .ZN(n792) );
  AOI22D1BWP30P140LVT U1187 ( .A1(n1234), .A2(i_data_bus[585]), .B1(n1240), 
        .B2(i_data_bus[617]), .ZN(n790) );
  AOI22D1BWP30P140LVT U1188 ( .A1(n1233), .A2(i_data_bus[553]), .B1(n117), 
        .B2(i_data_bus[105]), .ZN(n789) );
  ND4D1BWP30P140LVT U1189 ( .A1(n792), .A2(n791), .A3(n790), .A4(n789), .ZN(
        n808) );
  AOI22D1BWP30P140LVT U1190 ( .A1(n1230), .A2(i_data_bus[1001]), .B1(n1231), 
        .B2(i_data_bus[969]), .ZN(n796) );
  AOI22D1BWP30P140LVT U1191 ( .A1(n1232), .A2(i_data_bus[41]), .B1(n1242), 
        .B2(i_data_bus[937]), .ZN(n795) );
  AOI22D1BWP30P140LVT U1192 ( .A1(n1247), .A2(i_data_bus[489]), .B1(n1258), 
        .B2(i_data_bus[201]), .ZN(n794) );
  AOI22D1BWP30P140LVT U1193 ( .A1(n1254), .A2(i_data_bus[745]), .B1(n1269), 
        .B2(i_data_bus[233]), .ZN(n793) );
  ND4D1BWP30P140LVT U1194 ( .A1(n796), .A2(n795), .A3(n794), .A4(n793), .ZN(
        n807) );
  AOI22D1BWP30P140LVT U1195 ( .A1(n1264), .A2(i_data_bus[681]), .B1(n1244), 
        .B2(i_data_bus[297]), .ZN(n800) );
  AOI22D1BWP30P140LVT U1196 ( .A1(n1265), .A2(i_data_bus[169]), .B1(n617), 
        .B2(i_data_bus[873]), .ZN(n799) );
  AOI22D1BWP30P140LVT U1197 ( .A1(n1263), .A2(i_data_bus[137]), .B1(n1268), 
        .B2(i_data_bus[329]), .ZN(n798) );
  AOI22D1BWP30P140LVT U1198 ( .A1(n1245), .A2(i_data_bus[425]), .B1(n1252), 
        .B2(i_data_bus[713]), .ZN(n797) );
  ND4D1BWP30P140LVT U1199 ( .A1(n800), .A2(n799), .A3(n798), .A4(n797), .ZN(
        n806) );
  AOI22D1BWP30P140LVT U1200 ( .A1(n1256), .A2(i_data_bus[809]), .B1(n1246), 
        .B2(i_data_bus[265]), .ZN(n804) );
  AOI22D1BWP30P140LVT U1201 ( .A1(n1253), .A2(i_data_bus[777]), .B1(n1266), 
        .B2(i_data_bus[361]), .ZN(n803) );
  AOI22D1BWP30P140LVT U1202 ( .A1(n1257), .A2(i_data_bus[393]), .B1(n1267), 
        .B2(i_data_bus[457]), .ZN(n802) );
  AOI22D1BWP30P140LVT U1203 ( .A1(n600), .A2(i_data_bus[841]), .B1(n1255), 
        .B2(i_data_bus[649]), .ZN(n801) );
  ND4D1BWP30P140LVT U1204 ( .A1(n804), .A2(n803), .A3(n802), .A4(n801), .ZN(
        n805) );
  OR4D1BWP30P140LVT U1205 ( .A1(n808), .A2(n807), .A3(n806), .A4(n805), .Z(
        o_data_bus[41]) );
  AOI22D1BWP30P140LVT U1206 ( .A1(n1230), .A2(i_data_bus[1002]), .B1(n1233), 
        .B2(i_data_bus[554]), .ZN(n812) );
  AOI22D1BWP30P140LVT U1207 ( .A1(n1232), .A2(i_data_bus[42]), .B1(n25), .B2(
        i_data_bus[10]), .ZN(n811) );
  AOI22D1BWP30P140LVT U1208 ( .A1(n1231), .A2(i_data_bus[970]), .B1(n1240), 
        .B2(i_data_bus[618]), .ZN(n810) );
  AOI22D1BWP30P140LVT U1209 ( .A1(n117), .A2(i_data_bus[106]), .B1(n1229), 
        .B2(i_data_bus[74]), .ZN(n809) );
  ND4D1BWP30P140LVT U1210 ( .A1(n812), .A2(n811), .A3(n810), .A4(n809), .ZN(
        n828) );
  AOI22D1BWP30P140LVT U1211 ( .A1(n1234), .A2(i_data_bus[586]), .B1(n594), 
        .B2(i_data_bus[906]), .ZN(n816) );
  AOI22D1BWP30P140LVT U1212 ( .A1(n1241), .A2(i_data_bus[522]), .B1(n1242), 
        .B2(i_data_bus[938]), .ZN(n815) );
  AOI22D1BWP30P140LVT U1213 ( .A1(n1258), .A2(i_data_bus[202]), .B1(n1268), 
        .B2(i_data_bus[330]), .ZN(n814) );
  AOI22D1BWP30P140LVT U1214 ( .A1(n1247), .A2(i_data_bus[490]), .B1(n1269), 
        .B2(i_data_bus[234]), .ZN(n813) );
  ND4D1BWP30P140LVT U1215 ( .A1(n816), .A2(n815), .A3(n814), .A4(n813), .ZN(
        n827) );
  AOI22D1BWP30P140LVT U1216 ( .A1(n1255), .A2(i_data_bus[650]), .B1(n1253), 
        .B2(i_data_bus[778]), .ZN(n820) );
  AOI22D1BWP30P140LVT U1217 ( .A1(n600), .A2(i_data_bus[842]), .B1(n1265), 
        .B2(i_data_bus[170]), .ZN(n819) );
  AOI22D1BWP30P140LVT U1218 ( .A1(n1266), .A2(i_data_bus[362]), .B1(n1244), 
        .B2(i_data_bus[298]), .ZN(n818) );
  AOI22D1BWP30P140LVT U1219 ( .A1(n1257), .A2(i_data_bus[394]), .B1(n617), 
        .B2(i_data_bus[874]), .ZN(n817) );
  ND4D1BWP30P140LVT U1220 ( .A1(n820), .A2(n819), .A3(n818), .A4(n817), .ZN(
        n826) );
  AOI22D1BWP30P140LVT U1221 ( .A1(n1245), .A2(i_data_bus[426]), .B1(n1267), 
        .B2(i_data_bus[458]), .ZN(n824) );
  AOI22D1BWP30P140LVT U1222 ( .A1(n1252), .A2(i_data_bus[714]), .B1(n1256), 
        .B2(i_data_bus[810]), .ZN(n823) );
  AOI22D1BWP30P140LVT U1223 ( .A1(n1254), .A2(i_data_bus[746]), .B1(n1264), 
        .B2(i_data_bus[682]), .ZN(n822) );
  AOI22D1BWP30P140LVT U1224 ( .A1(n1263), .A2(i_data_bus[138]), .B1(n1246), 
        .B2(i_data_bus[266]), .ZN(n821) );
  ND4D1BWP30P140LVT U1225 ( .A1(n824), .A2(n823), .A3(n822), .A4(n821), .ZN(
        n825) );
  OR4D1BWP30P140LVT U1226 ( .A1(n828), .A2(n827), .A3(n826), .A4(n825), .Z(
        o_data_bus[42]) );
  AOI22D1BWP30P140LVT U1227 ( .A1(n1241), .A2(i_data_bus[523]), .B1(n1242), 
        .B2(i_data_bus[939]), .ZN(n832) );
  AOI22D1BWP30P140LVT U1228 ( .A1(n594), .A2(i_data_bus[907]), .B1(n1240), 
        .B2(i_data_bus[619]), .ZN(n831) );
  AOI22D1BWP30P140LVT U1229 ( .A1(n1230), .A2(i_data_bus[1003]), .B1(n25), 
        .B2(i_data_bus[11]), .ZN(n830) );
  ND4D1BWP30P140LVT U1230 ( .A1(n832), .A2(n831), .A3(n830), .A4(n829), .ZN(
        n848) );
  AOI22D1BWP30P140LVT U1231 ( .A1(n103), .A2(i_data_bus[43]), .B1(n1229), .B2(
        i_data_bus[75]), .ZN(n836) );
  AOI22D1BWP30P140LVT U1232 ( .A1(n1233), .A2(i_data_bus[555]), .B1(n1234), 
        .B2(i_data_bus[587]), .ZN(n835) );
  AOI22D1BWP30P140LVT U1233 ( .A1(n1266), .A2(i_data_bus[363]), .B1(n1258), 
        .B2(i_data_bus[203]), .ZN(n834) );
  AOI22D1BWP30P140LVT U1234 ( .A1(n1247), .A2(i_data_bus[491]), .B1(n1245), 
        .B2(i_data_bus[427]), .ZN(n833) );
  ND4D1BWP30P140LVT U1235 ( .A1(n836), .A2(n835), .A3(n834), .A4(n833), .ZN(
        n847) );
  AOI22D1BWP30P140LVT U1236 ( .A1(n1257), .A2(i_data_bus[395]), .B1(n1265), 
        .B2(i_data_bus[171]), .ZN(n840) );
  AOI22D1BWP30P140LVT U1237 ( .A1(n1267), .A2(i_data_bus[459]), .B1(n617), 
        .B2(i_data_bus[875]), .ZN(n839) );
  AOI22D1BWP30P140LVT U1238 ( .A1(n1254), .A2(i_data_bus[747]), .B1(n1263), 
        .B2(i_data_bus[139]), .ZN(n838) );
  AOI22D1BWP30P140LVT U1239 ( .A1(n600), .A2(i_data_bus[843]), .B1(n1256), 
        .B2(i_data_bus[811]), .ZN(n837) );
  ND4D1BWP30P140LVT U1240 ( .A1(n840), .A2(n839), .A3(n838), .A4(n837), .ZN(
        n846) );
  AOI22D1BWP30P140LVT U1241 ( .A1(n1253), .A2(i_data_bus[779]), .B1(n1269), 
        .B2(i_data_bus[235]), .ZN(n844) );
  AOI22D1BWP30P140LVT U1242 ( .A1(n1244), .A2(i_data_bus[299]), .B1(n1268), 
        .B2(i_data_bus[331]), .ZN(n843) );
  AOI22D1BWP30P140LVT U1243 ( .A1(n1255), .A2(i_data_bus[651]), .B1(n1264), 
        .B2(i_data_bus[683]), .ZN(n842) );
  AOI22D1BWP30P140LVT U1244 ( .A1(n1252), .A2(i_data_bus[715]), .B1(n1246), 
        .B2(i_data_bus[267]), .ZN(n841) );
  ND4D1BWP30P140LVT U1245 ( .A1(n844), .A2(n843), .A3(n842), .A4(n841), .ZN(
        n845) );
  OR4D1BWP30P140LVT U1246 ( .A1(n848), .A2(n847), .A3(n846), .A4(n845), .Z(
        o_data_bus[43]) );
  AOI22D1BWP30P140LVT U1247 ( .A1(n1242), .A2(i_data_bus[940]), .B1(n25), .B2(
        i_data_bus[12]), .ZN(n852) );
  AOI22D1BWP30P140LVT U1248 ( .A1(n1233), .A2(i_data_bus[556]), .B1(n1240), 
        .B2(i_data_bus[620]), .ZN(n851) );
  AOI22D1BWP30P140LVT U1249 ( .A1(n1232), .A2(i_data_bus[44]), .B1(n1229), 
        .B2(i_data_bus[76]), .ZN(n850) );
  ND4D1BWP30P140LVT U1250 ( .A1(n852), .A2(n851), .A3(n850), .A4(n849), .ZN(
        n868) );
  AOI22D1BWP30P140LVT U1251 ( .A1(n1230), .A2(i_data_bus[1004]), .B1(n1234), 
        .B2(i_data_bus[588]), .ZN(n856) );
  AOI22D1BWP30P140LVT U1252 ( .A1(n1253), .A2(i_data_bus[780]), .B1(n1267), 
        .B2(i_data_bus[460]), .ZN(n854) );
  AOI22D1BWP30P140LVT U1253 ( .A1(n1252), .A2(i_data_bus[716]), .B1(n1244), 
        .B2(i_data_bus[300]), .ZN(n853) );
  ND4D1BWP30P140LVT U1254 ( .A1(n856), .A2(n855), .A3(n854), .A4(n853), .ZN(
        n867) );
  AOI22D1BWP30P140LVT U1255 ( .A1(n1266), .A2(i_data_bus[364]), .B1(n1264), 
        .B2(i_data_bus[684]), .ZN(n860) );
  AOI22D1BWP30P140LVT U1256 ( .A1(n1245), .A2(i_data_bus[428]), .B1(n1246), 
        .B2(i_data_bus[268]), .ZN(n859) );
  AOI22D1BWP30P140LVT U1257 ( .A1(n1254), .A2(i_data_bus[748]), .B1(n1263), 
        .B2(i_data_bus[140]), .ZN(n858) );
  AOI22D1BWP30P140LVT U1258 ( .A1(n1258), .A2(i_data_bus[204]), .B1(n1256), 
        .B2(i_data_bus[812]), .ZN(n857) );
  ND4D1BWP30P140LVT U1259 ( .A1(n860), .A2(n859), .A3(n858), .A4(n857), .ZN(
        n866) );
  AOI22D1BWP30P140LVT U1260 ( .A1(n1257), .A2(i_data_bus[396]), .B1(n1269), 
        .B2(i_data_bus[236]), .ZN(n864) );
  AOI22D1BWP30P140LVT U1261 ( .A1(n1247), .A2(i_data_bus[492]), .B1(n600), 
        .B2(i_data_bus[844]), .ZN(n863) );
  AOI22D1BWP30P140LVT U1262 ( .A1(n1255), .A2(i_data_bus[652]), .B1(n617), 
        .B2(i_data_bus[876]), .ZN(n862) );
  AOI22D1BWP30P140LVT U1263 ( .A1(n1265), .A2(i_data_bus[172]), .B1(n1268), 
        .B2(i_data_bus[332]), .ZN(n861) );
  ND4D1BWP30P140LVT U1264 ( .A1(n864), .A2(n863), .A3(n862), .A4(n861), .ZN(
        n865) );
  OR4D1BWP30P140LVT U1265 ( .A1(n868), .A2(n867), .A3(n866), .A4(n865), .Z(
        o_data_bus[44]) );
  AOI22D1BWP30P140LVT U1266 ( .A1(n103), .A2(i_data_bus[45]), .B1(n1241), .B2(
        i_data_bus[525]), .ZN(n872) );
  AOI22D1BWP30P140LVT U1267 ( .A1(n594), .A2(i_data_bus[909]), .B1(n1240), 
        .B2(i_data_bus[621]), .ZN(n871) );
  AOI22D1BWP30P140LVT U1268 ( .A1(n1230), .A2(i_data_bus[1005]), .B1(n1234), 
        .B2(i_data_bus[589]), .ZN(n869) );
  ND4D1BWP30P140LVT U1269 ( .A1(n872), .A2(n871), .A3(n870), .A4(n869), .ZN(
        n888) );
  AOI22D1BWP30P140LVT U1270 ( .A1(n117), .A2(i_data_bus[109]), .B1(n1229), 
        .B2(i_data_bus[77]), .ZN(n876) );
  AOI22D1BWP30P140LVT U1271 ( .A1(n1242), .A2(i_data_bus[941]), .B1(n25), .B2(
        i_data_bus[13]), .ZN(n875) );
  AOI22D1BWP30P140LVT U1272 ( .A1(n1257), .A2(i_data_bus[397]), .B1(n1269), 
        .B2(i_data_bus[237]), .ZN(n874) );
  AOI22D1BWP30P140LVT U1273 ( .A1(n1266), .A2(i_data_bus[365]), .B1(n1246), 
        .B2(i_data_bus[269]), .ZN(n873) );
  ND4D1BWP30P140LVT U1274 ( .A1(n876), .A2(n875), .A3(n874), .A4(n873), .ZN(
        n887) );
  AOI22D1BWP30P140LVT U1275 ( .A1(n1247), .A2(i_data_bus[493]), .B1(n1245), 
        .B2(i_data_bus[429]), .ZN(n880) );
  AOI22D1BWP30P140LVT U1276 ( .A1(n1263), .A2(i_data_bus[141]), .B1(n617), 
        .B2(i_data_bus[877]), .ZN(n879) );
  AOI22D1BWP30P140LVT U1277 ( .A1(n1254), .A2(i_data_bus[749]), .B1(n1253), 
        .B2(i_data_bus[781]), .ZN(n878) );
  AOI22D1BWP30P140LVT U1278 ( .A1(n1258), .A2(i_data_bus[205]), .B1(n1244), 
        .B2(i_data_bus[301]), .ZN(n877) );
  ND4D1BWP30P140LVT U1279 ( .A1(n880), .A2(n879), .A3(n878), .A4(n877), .ZN(
        n886) );
  AOI22D1BWP30P140LVT U1280 ( .A1(n600), .A2(i_data_bus[845]), .B1(n1264), 
        .B2(i_data_bus[685]), .ZN(n884) );
  AOI22D1BWP30P140LVT U1281 ( .A1(n1255), .A2(i_data_bus[653]), .B1(n1268), 
        .B2(i_data_bus[333]), .ZN(n883) );
  AOI22D1BWP30P140LVT U1282 ( .A1(n1265), .A2(i_data_bus[173]), .B1(n1256), 
        .B2(i_data_bus[813]), .ZN(n882) );
  AOI22D1BWP30P140LVT U1283 ( .A1(n1267), .A2(i_data_bus[461]), .B1(n1252), 
        .B2(i_data_bus[717]), .ZN(n881) );
  ND4D1BWP30P140LVT U1284 ( .A1(n884), .A2(n883), .A3(n882), .A4(n881), .ZN(
        n885) );
  OR4D1BWP30P140LVT U1285 ( .A1(n888), .A2(n887), .A3(n886), .A4(n885), .Z(
        o_data_bus[45]) );
  AOI22D1BWP30P140LVT U1286 ( .A1(n117), .A2(i_data_bus[110]), .B1(n594), .B2(
        i_data_bus[910]), .ZN(n892) );
  AOI22D1BWP30P140LVT U1287 ( .A1(n1230), .A2(i_data_bus[1006]), .B1(n1229), 
        .B2(i_data_bus[78]), .ZN(n891) );
  AOI22D1BWP30P140LVT U1288 ( .A1(n25), .A2(i_data_bus[14]), .B1(n1234), .B2(
        i_data_bus[590]), .ZN(n890) );
  AOI22D1BWP30P140LVT U1289 ( .A1(n103), .A2(i_data_bus[46]), .B1(n1233), .B2(
        i_data_bus[558]), .ZN(n889) );
  ND4D1BWP30P140LVT U1290 ( .A1(n892), .A2(n891), .A3(n890), .A4(n889), .ZN(
        n908) );
  AOI22D1BWP30P140LVT U1291 ( .A1(n1242), .A2(i_data_bus[942]), .B1(n1231), 
        .B2(i_data_bus[974]), .ZN(n896) );
  AOI22D1BWP30P140LVT U1292 ( .A1(n1241), .A2(i_data_bus[526]), .B1(n1240), 
        .B2(i_data_bus[622]), .ZN(n895) );
  AOI22D1BWP30P140LVT U1293 ( .A1(n1265), .A2(i_data_bus[174]), .B1(n1246), 
        .B2(i_data_bus[270]), .ZN(n894) );
  AOI22D1BWP30P140LVT U1294 ( .A1(n1266), .A2(i_data_bus[366]), .B1(n1258), 
        .B2(i_data_bus[206]), .ZN(n893) );
  ND4D1BWP30P140LVT U1295 ( .A1(n896), .A2(n895), .A3(n894), .A4(n893), .ZN(
        n907) );
  AOI22D1BWP30P140LVT U1296 ( .A1(n1267), .A2(i_data_bus[462]), .B1(n1269), 
        .B2(i_data_bus[238]), .ZN(n900) );
  AOI22D1BWP30P140LVT U1297 ( .A1(n1263), .A2(i_data_bus[142]), .B1(n1256), 
        .B2(i_data_bus[814]), .ZN(n899) );
  AOI22D1BWP30P140LVT U1298 ( .A1(n600), .A2(i_data_bus[846]), .B1(n1244), 
        .B2(i_data_bus[302]), .ZN(n898) );
  AOI22D1BWP30P140LVT U1299 ( .A1(n1253), .A2(i_data_bus[782]), .B1(n1268), 
        .B2(i_data_bus[334]), .ZN(n897) );
  ND4D1BWP30P140LVT U1300 ( .A1(n900), .A2(n899), .A3(n898), .A4(n897), .ZN(
        n906) );
  AOI22D1BWP30P140LVT U1301 ( .A1(n1264), .A2(i_data_bus[686]), .B1(n617), 
        .B2(i_data_bus[878]), .ZN(n904) );
  AOI22D1BWP30P140LVT U1302 ( .A1(n1257), .A2(i_data_bus[398]), .B1(n1245), 
        .B2(i_data_bus[430]), .ZN(n903) );
  AOI22D1BWP30P140LVT U1303 ( .A1(n1247), .A2(i_data_bus[494]), .B1(n1254), 
        .B2(i_data_bus[750]), .ZN(n902) );
  AOI22D1BWP30P140LVT U1304 ( .A1(n1255), .A2(i_data_bus[654]), .B1(n1252), 
        .B2(i_data_bus[718]), .ZN(n901) );
  ND4D1BWP30P140LVT U1305 ( .A1(n904), .A2(n903), .A3(n902), .A4(n901), .ZN(
        n905) );
  OR4D1BWP30P140LVT U1306 ( .A1(n908), .A2(n907), .A3(n906), .A4(n905), .Z(
        o_data_bus[46]) );
  AOI22D1BWP30P140LVT U1307 ( .A1(n1229), .A2(i_data_bus[79]), .B1(n1231), 
        .B2(i_data_bus[975]), .ZN(n912) );
  AOI22D1BWP30P140LVT U1308 ( .A1(n1233), .A2(i_data_bus[559]), .B1(n117), 
        .B2(i_data_bus[111]), .ZN(n910) );
  AOI22D1BWP30P140LVT U1309 ( .A1(n1232), .A2(i_data_bus[47]), .B1(n1241), 
        .B2(i_data_bus[527]), .ZN(n909) );
  ND4D1BWP30P140LVT U1310 ( .A1(n912), .A2(n911), .A3(n910), .A4(n909), .ZN(
        n928) );
  AOI22D1BWP30P140LVT U1311 ( .A1(n25), .A2(i_data_bus[15]), .B1(n1240), .B2(
        i_data_bus[623]), .ZN(n916) );
  AOI22D1BWP30P140LVT U1312 ( .A1(n1230), .A2(i_data_bus[1007]), .B1(n1242), 
        .B2(i_data_bus[943]), .ZN(n915) );
  AOI22D1BWP30P140LVT U1313 ( .A1(n1254), .A2(i_data_bus[751]), .B1(n1252), 
        .B2(i_data_bus[719]), .ZN(n914) );
  AOI22D1BWP30P140LVT U1314 ( .A1(n600), .A2(i_data_bus[847]), .B1(n1246), 
        .B2(i_data_bus[271]), .ZN(n913) );
  ND4D1BWP30P140LVT U1315 ( .A1(n916), .A2(n915), .A3(n914), .A4(n913), .ZN(
        n927) );
  AOI22D1BWP30P140LVT U1316 ( .A1(n1245), .A2(i_data_bus[431]), .B1(n1258), 
        .B2(i_data_bus[207]), .ZN(n920) );
  AOI22D1BWP30P140LVT U1317 ( .A1(n1265), .A2(i_data_bus[175]), .B1(n1269), 
        .B2(i_data_bus[239]), .ZN(n919) );
  AOI22D1BWP30P140LVT U1318 ( .A1(n1247), .A2(i_data_bus[495]), .B1(n1263), 
        .B2(i_data_bus[143]), .ZN(n918) );
  AOI22D1BWP30P140LVT U1319 ( .A1(n1255), .A2(i_data_bus[655]), .B1(n1267), 
        .B2(i_data_bus[463]), .ZN(n917) );
  ND4D1BWP30P140LVT U1320 ( .A1(n920), .A2(n919), .A3(n918), .A4(n917), .ZN(
        n926) );
  AOI22D1BWP30P140LVT U1321 ( .A1(n1253), .A2(i_data_bus[783]), .B1(n617), 
        .B2(i_data_bus[879]), .ZN(n924) );
  AOI22D1BWP30P140LVT U1322 ( .A1(n1257), .A2(i_data_bus[399]), .B1(n1256), 
        .B2(i_data_bus[815]), .ZN(n923) );
  AOI22D1BWP30P140LVT U1323 ( .A1(n1264), .A2(i_data_bus[687]), .B1(n1268), 
        .B2(i_data_bus[335]), .ZN(n922) );
  AOI22D1BWP30P140LVT U1324 ( .A1(n1266), .A2(i_data_bus[367]), .B1(n1244), 
        .B2(i_data_bus[303]), .ZN(n921) );
  ND4D1BWP30P140LVT U1325 ( .A1(n924), .A2(n923), .A3(n922), .A4(n921), .ZN(
        n925) );
  OR4D1BWP30P140LVT U1326 ( .A1(n928), .A2(n927), .A3(n926), .A4(n925), .Z(
        o_data_bus[47]) );
  AOI22D1BWP30P140LVT U1327 ( .A1(n1233), .A2(i_data_bus[560]), .B1(n1242), 
        .B2(i_data_bus[944]), .ZN(n932) );
  AOI22D1BWP30P140LVT U1328 ( .A1(n1232), .A2(i_data_bus[48]), .B1(n1229), 
        .B2(i_data_bus[80]), .ZN(n931) );
  AOI22D1BWP30P140LVT U1329 ( .A1(n1241), .A2(i_data_bus[528]), .B1(n1240), 
        .B2(i_data_bus[624]), .ZN(n930) );
  AOI22D1BWP30P140LVT U1330 ( .A1(n1231), .A2(i_data_bus[976]), .B1(n594), 
        .B2(i_data_bus[912]), .ZN(n929) );
  ND4D1BWP30P140LVT U1331 ( .A1(n932), .A2(n931), .A3(n930), .A4(n929), .ZN(
        n948) );
  AOI22D1BWP30P140LVT U1332 ( .A1(n117), .A2(i_data_bus[112]), .B1(n1234), 
        .B2(i_data_bus[592]), .ZN(n936) );
  AOI22D1BWP30P140LVT U1333 ( .A1(n1230), .A2(i_data_bus[1008]), .B1(n25), 
        .B2(i_data_bus[16]), .ZN(n935) );
  AOI22D1BWP30P140LVT U1334 ( .A1(n1245), .A2(i_data_bus[432]), .B1(n1244), 
        .B2(i_data_bus[304]), .ZN(n934) );
  AOI22D1BWP30P140LVT U1335 ( .A1(n1247), .A2(i_data_bus[496]), .B1(n1268), 
        .B2(i_data_bus[336]), .ZN(n933) );
  ND4D1BWP30P140LVT U1336 ( .A1(n936), .A2(n935), .A3(n934), .A4(n933), .ZN(
        n947) );
  AOI22D1BWP30P140LVT U1337 ( .A1(n1263), .A2(i_data_bus[144]), .B1(n617), 
        .B2(i_data_bus[880]), .ZN(n940) );
  AOI22D1BWP30P140LVT U1338 ( .A1(n1255), .A2(i_data_bus[656]), .B1(n1253), 
        .B2(i_data_bus[784]), .ZN(n939) );
  AOI22D1BWP30P140LVT U1339 ( .A1(n1254), .A2(i_data_bus[752]), .B1(n1252), 
        .B2(i_data_bus[720]), .ZN(n938) );
  AOI22D1BWP30P140LVT U1340 ( .A1(n1258), .A2(i_data_bus[208]), .B1(n1256), 
        .B2(i_data_bus[816]), .ZN(n937) );
  ND4D1BWP30P140LVT U1341 ( .A1(n940), .A2(n939), .A3(n938), .A4(n937), .ZN(
        n946) );
  AOI22D1BWP30P140LVT U1342 ( .A1(n1267), .A2(i_data_bus[464]), .B1(n1246), 
        .B2(i_data_bus[272]), .ZN(n944) );
  AOI22D1BWP30P140LVT U1343 ( .A1(n1265), .A2(i_data_bus[176]), .B1(n1266), 
        .B2(i_data_bus[368]), .ZN(n943) );
  AOI22D1BWP30P140LVT U1344 ( .A1(n1257), .A2(i_data_bus[400]), .B1(n1269), 
        .B2(i_data_bus[240]), .ZN(n942) );
  AOI22D1BWP30P140LVT U1345 ( .A1(n600), .A2(i_data_bus[848]), .B1(n1264), 
        .B2(i_data_bus[688]), .ZN(n941) );
  ND4D1BWP30P140LVT U1346 ( .A1(n944), .A2(n943), .A3(n942), .A4(n941), .ZN(
        n945) );
  OR4D1BWP30P140LVT U1347 ( .A1(n945), .A2(n947), .A3(n946), .A4(n948), .Z(
        o_data_bus[48]) );
  AOI22D1BWP30P140LVT U1348 ( .A1(n25), .A2(i_data_bus[17]), .B1(n1240), .B2(
        i_data_bus[625]), .ZN(n952) );
  AOI22D1BWP30P140LVT U1349 ( .A1(n1230), .A2(i_data_bus[1009]), .B1(n103), 
        .B2(i_data_bus[49]), .ZN(n951) );
  AOI22D1BWP30P140LVT U1350 ( .A1(n1242), .A2(i_data_bus[945]), .B1(n1234), 
        .B2(i_data_bus[593]), .ZN(n949) );
  ND4D1BWP30P140LVT U1351 ( .A1(n952), .A2(n951), .A3(n950), .A4(n949), .ZN(
        n968) );
  AOI22D1BWP30P140LVT U1352 ( .A1(n117), .A2(i_data_bus[113]), .B1(n1231), 
        .B2(i_data_bus[977]), .ZN(n956) );
  AOI22D1BWP30P140LVT U1353 ( .A1(n1233), .A2(i_data_bus[561]), .B1(n1241), 
        .B2(i_data_bus[529]), .ZN(n955) );
  AOI22D1BWP30P140LVT U1354 ( .A1(n1264), .A2(i_data_bus[689]), .B1(n617), 
        .B2(i_data_bus[881]), .ZN(n954) );
  AOI22D1BWP30P140LVT U1355 ( .A1(n1245), .A2(i_data_bus[433]), .B1(n600), 
        .B2(i_data_bus[849]), .ZN(n953) );
  ND4D1BWP30P140LVT U1356 ( .A1(n956), .A2(n955), .A3(n954), .A4(n953), .ZN(
        n967) );
  AOI22D1BWP30P140LVT U1357 ( .A1(n1263), .A2(i_data_bus[145]), .B1(n1268), 
        .B2(i_data_bus[337]), .ZN(n960) );
  AOI22D1BWP30P140LVT U1358 ( .A1(n1257), .A2(i_data_bus[401]), .B1(n1269), 
        .B2(i_data_bus[241]), .ZN(n959) );
  AOI22D1BWP30P140LVT U1359 ( .A1(n1253), .A2(i_data_bus[785]), .B1(n1258), 
        .B2(i_data_bus[209]), .ZN(n958) );
  AOI22D1BWP30P140LVT U1360 ( .A1(n1252), .A2(i_data_bus[721]), .B1(n1246), 
        .B2(i_data_bus[273]), .ZN(n957) );
  ND4D1BWP30P140LVT U1361 ( .A1(n960), .A2(n959), .A3(n958), .A4(n957), .ZN(
        n966) );
  AOI22D1BWP30P140LVT U1362 ( .A1(n1265), .A2(i_data_bus[177]), .B1(n1244), 
        .B2(i_data_bus[305]), .ZN(n964) );
  AOI22D1BWP30P140LVT U1363 ( .A1(n1255), .A2(i_data_bus[657]), .B1(n1254), 
        .B2(i_data_bus[753]), .ZN(n963) );
  AOI22D1BWP30P140LVT U1364 ( .A1(n1247), .A2(i_data_bus[497]), .B1(n1267), 
        .B2(i_data_bus[465]), .ZN(n962) );
  AOI22D1BWP30P140LVT U1365 ( .A1(n1266), .A2(i_data_bus[369]), .B1(n1256), 
        .B2(i_data_bus[817]), .ZN(n961) );
  ND4D1BWP30P140LVT U1366 ( .A1(n964), .A2(n963), .A3(n962), .A4(n961), .ZN(
        n965) );
  OR4D1BWP30P140LVT U1367 ( .A1(n968), .A2(n967), .A3(n966), .A4(n965), .Z(
        o_data_bus[49]) );
  AOI22D1BWP30P140LVT U1368 ( .A1(n1234), .A2(i_data_bus[594]), .B1(n1240), 
        .B2(i_data_bus[626]), .ZN(n972) );
  AOI22D1BWP30P140LVT U1369 ( .A1(n103), .A2(i_data_bus[50]), .B1(n1231), .B2(
        i_data_bus[978]), .ZN(n971) );
  AOI22D1BWP30P140LVT U1370 ( .A1(n117), .A2(i_data_bus[114]), .B1(n1241), 
        .B2(i_data_bus[530]), .ZN(n970) );
  AOI22D1BWP30P140LVT U1371 ( .A1(n1230), .A2(i_data_bus[1010]), .B1(n1233), 
        .B2(i_data_bus[562]), .ZN(n969) );
  ND4D1BWP30P140LVT U1372 ( .A1(n971), .A2(n972), .A3(n970), .A4(n969), .ZN(
        n988) );
  AOI22D1BWP30P140LVT U1373 ( .A1(n1229), .A2(i_data_bus[82]), .B1(n594), .B2(
        i_data_bus[914]), .ZN(n976) );
  AOI22D1BWP30P140LVT U1374 ( .A1(n1242), .A2(i_data_bus[946]), .B1(n25), .B2(
        i_data_bus[18]), .ZN(n975) );
  AOI22D1BWP30P140LVT U1375 ( .A1(n1252), .A2(i_data_bus[722]), .B1(n617), 
        .B2(i_data_bus[882]), .ZN(n974) );
  AOI22D1BWP30P140LVT U1376 ( .A1(n1257), .A2(i_data_bus[402]), .B1(n1269), 
        .B2(i_data_bus[242]), .ZN(n973) );
  ND4D1BWP30P140LVT U1377 ( .A1(n976), .A2(n975), .A3(n974), .A4(n973), .ZN(
        n987) );
  AOI22D1BWP30P140LVT U1378 ( .A1(n1258), .A2(i_data_bus[210]), .B1(n1256), 
        .B2(i_data_bus[818]), .ZN(n980) );
  AOI22D1BWP30P140LVT U1379 ( .A1(n1266), .A2(i_data_bus[370]), .B1(n1264), 
        .B2(i_data_bus[690]), .ZN(n979) );
  AOI22D1BWP30P140LVT U1380 ( .A1(n1247), .A2(i_data_bus[498]), .B1(n1265), 
        .B2(i_data_bus[178]), .ZN(n978) );
  AOI22D1BWP30P140LVT U1381 ( .A1(n600), .A2(i_data_bus[850]), .B1(n1244), 
        .B2(i_data_bus[306]), .ZN(n977) );
  ND4D1BWP30P140LVT U1382 ( .A1(n980), .A2(n979), .A3(n978), .A4(n977), .ZN(
        n986) );
  AOI22D1BWP30P140LVT U1383 ( .A1(n1255), .A2(i_data_bus[658]), .B1(n1267), 
        .B2(i_data_bus[466]), .ZN(n984) );
  AOI22D1BWP30P140LVT U1384 ( .A1(n1263), .A2(i_data_bus[146]), .B1(n1246), 
        .B2(i_data_bus[274]), .ZN(n983) );
  AOI22D1BWP30P140LVT U1385 ( .A1(n1254), .A2(i_data_bus[754]), .B1(n1253), 
        .B2(i_data_bus[786]), .ZN(n982) );
  AOI22D1BWP30P140LVT U1386 ( .A1(n1245), .A2(i_data_bus[434]), .B1(n1268), 
        .B2(i_data_bus[338]), .ZN(n981) );
  ND4D1BWP30P140LVT U1387 ( .A1(n984), .A2(n983), .A3(n982), .A4(n981), .ZN(
        n985) );
  OR4D1BWP30P140LVT U1388 ( .A1(n988), .A2(n986), .A3(n987), .A4(n985), .Z(
        o_data_bus[50]) );
  AOI22D1BWP30P140LVT U1389 ( .A1(n1233), .A2(i_data_bus[563]), .B1(n1231), 
        .B2(i_data_bus[979]), .ZN(n992) );
  AOI22D1BWP30P140LVT U1390 ( .A1(n103), .A2(i_data_bus[51]), .B1(n1241), .B2(
        i_data_bus[531]), .ZN(n991) );
  AOI22D1BWP30P140LVT U1391 ( .A1(n1230), .A2(i_data_bus[1011]), .B1(n117), 
        .B2(i_data_bus[115]), .ZN(n990) );
  AOI22D1BWP30P140LVT U1392 ( .A1(n1242), .A2(i_data_bus[947]), .B1(n1229), 
        .B2(i_data_bus[83]), .ZN(n989) );
  ND4D1BWP30P140LVT U1393 ( .A1(n992), .A2(n991), .A3(n990), .A4(n989), .ZN(
        n1008) );
  AOI22D1BWP30P140LVT U1394 ( .A1(n25), .A2(i_data_bus[19]), .B1(n594), .B2(
        i_data_bus[915]), .ZN(n996) );
  AOI22D1BWP30P140LVT U1395 ( .A1(n1234), .A2(i_data_bus[595]), .B1(n1240), 
        .B2(i_data_bus[627]), .ZN(n995) );
  AOI22D1BWP30P140LVT U1396 ( .A1(n1254), .A2(i_data_bus[755]), .B1(n1266), 
        .B2(i_data_bus[371]), .ZN(n994) );
  AOI22D1BWP30P140LVT U1397 ( .A1(n1265), .A2(i_data_bus[179]), .B1(n1258), 
        .B2(i_data_bus[211]), .ZN(n993) );
  ND4D1BWP30P140LVT U1398 ( .A1(n996), .A2(n995), .A3(n994), .A4(n993), .ZN(
        n1007) );
  AOI22D1BWP30P140LVT U1399 ( .A1(n1257), .A2(i_data_bus[403]), .B1(n1244), 
        .B2(i_data_bus[307]), .ZN(n1000) );
  AOI22D1BWP30P140LVT U1400 ( .A1(n1263), .A2(i_data_bus[147]), .B1(n1268), 
        .B2(i_data_bus[339]), .ZN(n999) );
  AOI22D1BWP30P140LVT U1401 ( .A1(n1269), .A2(i_data_bus[243]), .B1(n1256), 
        .B2(i_data_bus[819]), .ZN(n998) );
  AOI22D1BWP30P140LVT U1402 ( .A1(n1255), .A2(i_data_bus[659]), .B1(n1253), 
        .B2(i_data_bus[787]), .ZN(n997) );
  ND4D1BWP30P140LVT U1403 ( .A1(n1000), .A2(n999), .A3(n998), .A4(n997), .ZN(
        n1006) );
  AOI22D1BWP30P140LVT U1404 ( .A1(n600), .A2(i_data_bus[851]), .B1(n617), .B2(
        i_data_bus[883]), .ZN(n1004) );
  AOI22D1BWP30P140LVT U1405 ( .A1(n1247), .A2(i_data_bus[499]), .B1(n1264), 
        .B2(i_data_bus[691]), .ZN(n1003) );
  AOI22D1BWP30P140LVT U1406 ( .A1(n1245), .A2(i_data_bus[435]), .B1(n1252), 
        .B2(i_data_bus[723]), .ZN(n1002) );
  AOI22D1BWP30P140LVT U1407 ( .A1(n1267), .A2(i_data_bus[467]), .B1(n1246), 
        .B2(i_data_bus[275]), .ZN(n1001) );
  ND4D1BWP30P140LVT U1408 ( .A1(n1004), .A2(n1003), .A3(n1002), .A4(n1001), 
        .ZN(n1005) );
  OR4D1BWP30P140LVT U1409 ( .A1(n1008), .A2(n1007), .A3(n1006), .A4(n1005), 
        .Z(o_data_bus[51]) );
  AOI22D1BWP30P140LVT U1410 ( .A1(n1241), .A2(i_data_bus[532]), .B1(n1234), 
        .B2(i_data_bus[596]), .ZN(n1012) );
  AOI22D1BWP30P140LVT U1411 ( .A1(n1232), .A2(i_data_bus[52]), .B1(n1231), 
        .B2(i_data_bus[980]), .ZN(n1011) );
  AOI22D1BWP30P140LVT U1412 ( .A1(n1230), .A2(i_data_bus[1012]), .B1(n1233), 
        .B2(i_data_bus[564]), .ZN(n1010) );
  AOI22D1BWP30P140LVT U1413 ( .A1(n25), .A2(i_data_bus[20]), .B1(n1240), .B2(
        i_data_bus[628]), .ZN(n1009) );
  ND4D1BWP30P140LVT U1414 ( .A1(n1011), .A2(n1012), .A3(n1010), .A4(n1009), 
        .ZN(n1028) );
  AOI22D1BWP30P140LVT U1415 ( .A1(n1242), .A2(i_data_bus[948]), .B1(n1229), 
        .B2(i_data_bus[84]), .ZN(n1016) );
  AOI22D1BWP30P140LVT U1416 ( .A1(n117), .A2(i_data_bus[116]), .B1(n594), .B2(
        i_data_bus[916]), .ZN(n1015) );
  AOI22D1BWP30P140LVT U1417 ( .A1(n1252), .A2(i_data_bus[724]), .B1(n1258), 
        .B2(i_data_bus[212]), .ZN(n1014) );
  AOI22D1BWP30P140LVT U1418 ( .A1(n1269), .A2(i_data_bus[244]), .B1(n1268), 
        .B2(i_data_bus[340]), .ZN(n1013) );
  ND4D1BWP30P140LVT U1419 ( .A1(n1016), .A2(n1015), .A3(n1014), .A4(n1013), 
        .ZN(n1027) );
  AOI22D1BWP30P140LVT U1420 ( .A1(n1265), .A2(i_data_bus[180]), .B1(n1256), 
        .B2(i_data_bus[820]), .ZN(n1020) );
  AOI22D1BWP30P140LVT U1421 ( .A1(n600), .A2(i_data_bus[852]), .B1(n1253), 
        .B2(i_data_bus[788]), .ZN(n1019) );
  AOI22D1BWP30P140LVT U1422 ( .A1(n1254), .A2(i_data_bus[756]), .B1(n1246), 
        .B2(i_data_bus[276]), .ZN(n1018) );
  AOI22D1BWP30P140LVT U1423 ( .A1(n1255), .A2(i_data_bus[660]), .B1(n617), 
        .B2(i_data_bus[884]), .ZN(n1017) );
  ND4D1BWP30P140LVT U1424 ( .A1(n1020), .A2(n1019), .A3(n1018), .A4(n1017), 
        .ZN(n1026) );
  AOI22D1BWP30P140LVT U1425 ( .A1(n1257), .A2(i_data_bus[404]), .B1(n1245), 
        .B2(i_data_bus[436]), .ZN(n1024) );
  AOI22D1BWP30P140LVT U1426 ( .A1(n1267), .A2(i_data_bus[468]), .B1(n1264), 
        .B2(i_data_bus[692]), .ZN(n1023) );
  AOI22D1BWP30P140LVT U1427 ( .A1(n1263), .A2(i_data_bus[148]), .B1(n1244), 
        .B2(i_data_bus[308]), .ZN(n1022) );
  AOI22D1BWP30P140LVT U1428 ( .A1(n1247), .A2(i_data_bus[500]), .B1(n1266), 
        .B2(i_data_bus[372]), .ZN(n1021) );
  ND4D1BWP30P140LVT U1429 ( .A1(n1024), .A2(n1023), .A3(n1022), .A4(n1021), 
        .ZN(n1025) );
  OR4D1BWP30P140LVT U1430 ( .A1(n1028), .A2(n1027), .A3(n1026), .A4(n1025), 
        .Z(o_data_bus[52]) );
  AOI22D1BWP30P140LVT U1431 ( .A1(n103), .A2(i_data_bus[53]), .B1(n1242), .B2(
        i_data_bus[949]), .ZN(n1032) );
  AOI22D1BWP30P140LVT U1432 ( .A1(n117), .A2(i_data_bus[117]), .B1(n1240), 
        .B2(i_data_bus[629]), .ZN(n1031) );
  AOI22D1BWP30P140LVT U1433 ( .A1(n1231), .A2(i_data_bus[981]), .B1(n594), 
        .B2(i_data_bus[917]), .ZN(n1030) );
  AOI22D1BWP30P140LVT U1434 ( .A1(n25), .A2(i_data_bus[21]), .B1(n1234), .B2(
        i_data_bus[597]), .ZN(n1029) );
  ND4D1BWP30P140LVT U1435 ( .A1(n1030), .A2(n1032), .A3(n1031), .A4(n1029), 
        .ZN(n1048) );
  AOI22D1BWP30P140LVT U1436 ( .A1(n1233), .A2(i_data_bus[565]), .B1(n1241), 
        .B2(i_data_bus[533]), .ZN(n1036) );
  AOI22D1BWP30P140LVT U1437 ( .A1(n1230), .A2(i_data_bus[1013]), .B1(n1229), 
        .B2(i_data_bus[85]), .ZN(n1035) );
  AOI22D1BWP30P140LVT U1438 ( .A1(n1255), .A2(i_data_bus[661]), .B1(n1254), 
        .B2(i_data_bus[757]), .ZN(n1034) );
  AOI22D1BWP30P140LVT U1439 ( .A1(n600), .A2(i_data_bus[853]), .B1(n1268), 
        .B2(i_data_bus[341]), .ZN(n1033) );
  ND4D1BWP30P140LVT U1440 ( .A1(n1036), .A2(n1035), .A3(n1034), .A4(n1033), 
        .ZN(n1047) );
  AOI22D1BWP30P140LVT U1441 ( .A1(n1253), .A2(i_data_bus[789]), .B1(n1263), 
        .B2(i_data_bus[149]), .ZN(n1040) );
  AOI22D1BWP30P140LVT U1442 ( .A1(n1265), .A2(i_data_bus[181]), .B1(n1256), 
        .B2(i_data_bus[821]), .ZN(n1039) );
  AOI22D1BWP30P140LVT U1443 ( .A1(n1247), .A2(i_data_bus[501]), .B1(n1245), 
        .B2(i_data_bus[437]), .ZN(n1038) );
  AOI22D1BWP30P140LVT U1444 ( .A1(n1252), .A2(i_data_bus[725]), .B1(n1258), 
        .B2(i_data_bus[213]), .ZN(n1037) );
  ND4D1BWP30P140LVT U1445 ( .A1(n1040), .A2(n1039), .A3(n1038), .A4(n1037), 
        .ZN(n1046) );
  AOI22D1BWP30P140LVT U1446 ( .A1(n1264), .A2(i_data_bus[693]), .B1(n1244), 
        .B2(i_data_bus[309]), .ZN(n1044) );
  AOI22D1BWP30P140LVT U1447 ( .A1(n1267), .A2(i_data_bus[469]), .B1(n1269), 
        .B2(i_data_bus[245]), .ZN(n1043) );
  AOI22D1BWP30P140LVT U1448 ( .A1(n1257), .A2(i_data_bus[405]), .B1(n1246), 
        .B2(i_data_bus[277]), .ZN(n1042) );
  AOI22D1BWP30P140LVT U1449 ( .A1(n1266), .A2(i_data_bus[373]), .B1(n617), 
        .B2(i_data_bus[885]), .ZN(n1041) );
  ND4D1BWP30P140LVT U1450 ( .A1(n1044), .A2(n1043), .A3(n1042), .A4(n1041), 
        .ZN(n1045) );
  OR4D1BWP30P140LVT U1451 ( .A1(n1048), .A2(n1047), .A3(n1046), .A4(n1045), 
        .Z(o_data_bus[53]) );
  AOI22D1BWP30P140LVT U1452 ( .A1(n1230), .A2(i_data_bus[1014]), .B1(n1232), 
        .B2(i_data_bus[54]), .ZN(n1052) );
  AOI22D1BWP30P140LVT U1453 ( .A1(n1233), .A2(i_data_bus[566]), .B1(n1241), 
        .B2(i_data_bus[534]), .ZN(n1051) );
  AOI22D1BWP30P140LVT U1454 ( .A1(n117), .A2(i_data_bus[118]), .B1(n1234), 
        .B2(i_data_bus[598]), .ZN(n1050) );
  AOI22D1BWP30P140LVT U1455 ( .A1(n1242), .A2(i_data_bus[950]), .B1(n594), 
        .B2(i_data_bus[918]), .ZN(n1049) );
  ND4D1BWP30P140LVT U1456 ( .A1(n1049), .A2(n1051), .A3(n1050), .A4(n1052), 
        .ZN(n1068) );
  AOI22D1BWP30P140LVT U1457 ( .A1(n25), .A2(i_data_bus[22]), .B1(n1229), .B2(
        i_data_bus[86]), .ZN(n1056) );
  AOI22D1BWP30P140LVT U1458 ( .A1(n1231), .A2(i_data_bus[982]), .B1(n1240), 
        .B2(i_data_bus[630]), .ZN(n1055) );
  AOI22D1BWP30P140LVT U1459 ( .A1(n1264), .A2(i_data_bus[694]), .B1(n1256), 
        .B2(i_data_bus[822]), .ZN(n1054) );
  AOI22D1BWP30P140LVT U1460 ( .A1(n1245), .A2(i_data_bus[438]), .B1(n1254), 
        .B2(i_data_bus[758]), .ZN(n1053) );
  ND4D1BWP30P140LVT U1461 ( .A1(n1056), .A2(n1055), .A3(n1054), .A4(n1053), 
        .ZN(n1067) );
  AOI22D1BWP30P140LVT U1462 ( .A1(n1253), .A2(i_data_bus[790]), .B1(n1269), 
        .B2(i_data_bus[246]), .ZN(n1060) );
  AOI22D1BWP30P140LVT U1463 ( .A1(n1257), .A2(i_data_bus[406]), .B1(n1266), 
        .B2(i_data_bus[374]), .ZN(n1059) );
  AOI22D1BWP30P140LVT U1464 ( .A1(n1247), .A2(i_data_bus[502]), .B1(n1265), 
        .B2(i_data_bus[182]), .ZN(n1058) );
  AOI22D1BWP30P140LVT U1465 ( .A1(n1263), .A2(i_data_bus[150]), .B1(n1252), 
        .B2(i_data_bus[726]), .ZN(n1057) );
  ND4D1BWP30P140LVT U1466 ( .A1(n1060), .A2(n1059), .A3(n1058), .A4(n1057), 
        .ZN(n1066) );
  AOI22D1BWP30P140LVT U1467 ( .A1(n617), .A2(i_data_bus[886]), .B1(n1244), 
        .B2(i_data_bus[310]), .ZN(n1064) );
  AOI22D1BWP30P140LVT U1468 ( .A1(n1267), .A2(i_data_bus[470]), .B1(n1268), 
        .B2(i_data_bus[342]), .ZN(n1063) );
  AOI22D1BWP30P140LVT U1469 ( .A1(n600), .A2(i_data_bus[854]), .B1(n1246), 
        .B2(i_data_bus[278]), .ZN(n1062) );
  AOI22D1BWP30P140LVT U1470 ( .A1(n1255), .A2(i_data_bus[662]), .B1(n1258), 
        .B2(i_data_bus[214]), .ZN(n1061) );
  ND4D1BWP30P140LVT U1471 ( .A1(n1064), .A2(n1063), .A3(n1062), .A4(n1061), 
        .ZN(n1065) );
  OR4D1BWP30P140LVT U1472 ( .A1(n1068), .A2(n1067), .A3(n1066), .A4(n1065), 
        .Z(o_data_bus[54]) );
  AOI22D1BWP30P140LVT U1473 ( .A1(n25), .A2(i_data_bus[23]), .B1(n1240), .B2(
        i_data_bus[631]), .ZN(n1072) );
  AOI22D1BWP30P140LVT U1474 ( .A1(n1230), .A2(i_data_bus[1015]), .B1(n1232), 
        .B2(i_data_bus[55]), .ZN(n1071) );
  AOI22D1BWP30P140LVT U1475 ( .A1(n1234), .A2(i_data_bus[599]), .B1(n1229), 
        .B2(i_data_bus[87]), .ZN(n1070) );
  ND4D1BWP30P140LVT U1476 ( .A1(n1072), .A2(n1071), .A3(n1070), .A4(n1069), 
        .ZN(n1088) );
  AOI22D1BWP30P140LVT U1477 ( .A1(n1241), .A2(i_data_bus[535]), .B1(n1231), 
        .B2(i_data_bus[983]), .ZN(n1076) );
  AOI22D1BWP30P140LVT U1478 ( .A1(n1233), .A2(i_data_bus[567]), .B1(n594), 
        .B2(i_data_bus[919]), .ZN(n1075) );
  AOI22D1BWP30P140LVT U1479 ( .A1(n1264), .A2(i_data_bus[695]), .B1(n1269), 
        .B2(i_data_bus[247]), .ZN(n1074) );
  AOI22D1BWP30P140LVT U1480 ( .A1(n1267), .A2(i_data_bus[471]), .B1(n617), 
        .B2(i_data_bus[887]), .ZN(n1073) );
  ND4D1BWP30P140LVT U1481 ( .A1(n1076), .A2(n1075), .A3(n1074), .A4(n1073), 
        .ZN(n1087) );
  AOI22D1BWP30P140LVT U1482 ( .A1(n1265), .A2(i_data_bus[183]), .B1(n1244), 
        .B2(i_data_bus[311]), .ZN(n1080) );
  AOI22D1BWP30P140LVT U1483 ( .A1(n1254), .A2(i_data_bus[759]), .B1(n1246), 
        .B2(i_data_bus[279]), .ZN(n1079) );
  AOI22D1BWP30P140LVT U1484 ( .A1(n1247), .A2(i_data_bus[503]), .B1(n1258), 
        .B2(i_data_bus[215]), .ZN(n1078) );
  AOI22D1BWP30P140LVT U1485 ( .A1(n1245), .A2(i_data_bus[439]), .B1(n1252), 
        .B2(i_data_bus[727]), .ZN(n1077) );
  ND4D1BWP30P140LVT U1486 ( .A1(n1080), .A2(n1079), .A3(n1078), .A4(n1077), 
        .ZN(n1086) );
  AOI22D1BWP30P140LVT U1487 ( .A1(n1257), .A2(i_data_bus[407]), .B1(n1263), 
        .B2(i_data_bus[151]), .ZN(n1084) );
  AOI22D1BWP30P140LVT U1488 ( .A1(n1255), .A2(i_data_bus[663]), .B1(n1256), 
        .B2(i_data_bus[823]), .ZN(n1083) );
  AOI22D1BWP30P140LVT U1489 ( .A1(n1253), .A2(i_data_bus[791]), .B1(n1266), 
        .B2(i_data_bus[375]), .ZN(n1082) );
  AOI22D1BWP30P140LVT U1490 ( .A1(n600), .A2(i_data_bus[855]), .B1(n1268), 
        .B2(i_data_bus[343]), .ZN(n1081) );
  ND4D1BWP30P140LVT U1491 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n1081), 
        .ZN(n1085) );
  OR4D1BWP30P140LVT U1492 ( .A1(n1088), .A2(n1087), .A3(n1086), .A4(n1085), 
        .Z(o_data_bus[55]) );
  AOI22D1BWP30P140LVT U1493 ( .A1(n1231), .A2(i_data_bus[984]), .B1(n1240), 
        .B2(i_data_bus[632]), .ZN(n1092) );
  AOI22D1BWP30P140LVT U1494 ( .A1(n117), .A2(i_data_bus[120]), .B1(n1229), 
        .B2(i_data_bus[88]), .ZN(n1091) );
  AOI22D1BWP30P140LVT U1495 ( .A1(n1230), .A2(i_data_bus[1016]), .B1(n1234), 
        .B2(i_data_bus[600]), .ZN(n1090) );
  AOI22D1BWP30P140LVT U1496 ( .A1(n1241), .A2(i_data_bus[536]), .B1(n25), .B2(
        i_data_bus[24]), .ZN(n1089) );
  ND4D1BWP30P140LVT U1497 ( .A1(n1092), .A2(n1091), .A3(n1090), .A4(n1089), 
        .ZN(n1108) );
  AOI22D1BWP30P140LVT U1498 ( .A1(n1232), .A2(i_data_bus[56]), .B1(n1242), 
        .B2(i_data_bus[952]), .ZN(n1096) );
  AOI22D1BWP30P140LVT U1499 ( .A1(n1233), .A2(i_data_bus[568]), .B1(n594), 
        .B2(i_data_bus[920]), .ZN(n1095) );
  AOI22D1BWP30P140LVT U1500 ( .A1(n1253), .A2(i_data_bus[792]), .B1(n1246), 
        .B2(i_data_bus[280]), .ZN(n1094) );
  AOI22D1BWP30P140LVT U1501 ( .A1(n1264), .A2(i_data_bus[696]), .B1(n1269), 
        .B2(i_data_bus[248]), .ZN(n1093) );
  ND4D1BWP30P140LVT U1502 ( .A1(n1096), .A2(n1095), .A3(n1094), .A4(n1093), 
        .ZN(n1107) );
  AOI22D1BWP30P140LVT U1503 ( .A1(n1257), .A2(i_data_bus[408]), .B1(n1268), 
        .B2(i_data_bus[344]), .ZN(n1100) );
  AOI22D1BWP30P140LVT U1504 ( .A1(n1245), .A2(i_data_bus[440]), .B1(n600), 
        .B2(i_data_bus[856]), .ZN(n1099) );
  AOI22D1BWP30P140LVT U1505 ( .A1(n1255), .A2(i_data_bus[664]), .B1(n1256), 
        .B2(i_data_bus[824]), .ZN(n1098) );
  AOI22D1BWP30P140LVT U1506 ( .A1(n1266), .A2(i_data_bus[376]), .B1(n1252), 
        .B2(i_data_bus[728]), .ZN(n1097) );
  ND4D1BWP30P140LVT U1507 ( .A1(n1100), .A2(n1099), .A3(n1098), .A4(n1097), 
        .ZN(n1106) );
  AOI22D1BWP30P140LVT U1508 ( .A1(n1263), .A2(i_data_bus[152]), .B1(n617), 
        .B2(i_data_bus[888]), .ZN(n1104) );
  AOI22D1BWP30P140LVT U1509 ( .A1(n1265), .A2(i_data_bus[184]), .B1(n1267), 
        .B2(i_data_bus[472]), .ZN(n1103) );
  AOI22D1BWP30P140LVT U1510 ( .A1(n1247), .A2(i_data_bus[504]), .B1(n1258), 
        .B2(i_data_bus[216]), .ZN(n1102) );
  AOI22D1BWP30P140LVT U1511 ( .A1(n1254), .A2(i_data_bus[760]), .B1(n1244), 
        .B2(i_data_bus[312]), .ZN(n1101) );
  ND4D1BWP30P140LVT U1512 ( .A1(n1104), .A2(n1103), .A3(n1102), .A4(n1101), 
        .ZN(n1105) );
  OR4D1BWP30P140LVT U1513 ( .A1(n1108), .A2(n1107), .A3(n1106), .A4(n1105), 
        .Z(o_data_bus[56]) );
  AOI22D1BWP30P140LVT U1514 ( .A1(n1230), .A2(i_data_bus[1017]), .B1(n1232), 
        .B2(i_data_bus[57]), .ZN(n1112) );
  AOI22D1BWP30P140LVT U1515 ( .A1(n1234), .A2(i_data_bus[601]), .B1(n1240), 
        .B2(i_data_bus[633]), .ZN(n1110) );
  AOI22D1BWP30P140LVT U1516 ( .A1(n117), .A2(i_data_bus[121]), .B1(n1241), 
        .B2(i_data_bus[537]), .ZN(n1109) );
  ND4D1BWP30P140LVT U1517 ( .A1(n1112), .A2(n1111), .A3(n1110), .A4(n1109), 
        .ZN(n1128) );
  AOI22D1BWP30P140LVT U1518 ( .A1(n25), .A2(i_data_bus[25]), .B1(n1231), .B2(
        i_data_bus[985]), .ZN(n1116) );
  AOI22D1BWP30P140LVT U1519 ( .A1(n1242), .A2(i_data_bus[953]), .B1(n1229), 
        .B2(i_data_bus[89]), .ZN(n1115) );
  AOI22D1BWP30P140LVT U1520 ( .A1(n1252), .A2(i_data_bus[729]), .B1(n1256), 
        .B2(i_data_bus[825]), .ZN(n1114) );
  AOI22D1BWP30P140LVT U1521 ( .A1(n1255), .A2(i_data_bus[665]), .B1(n1264), 
        .B2(i_data_bus[697]), .ZN(n1113) );
  ND4D1BWP30P140LVT U1522 ( .A1(n1116), .A2(n1115), .A3(n1114), .A4(n1113), 
        .ZN(n1127) );
  AOI22D1BWP30P140LVT U1523 ( .A1(n1265), .A2(i_data_bus[185]), .B1(n1268), 
        .B2(i_data_bus[345]), .ZN(n1120) );
  AOI22D1BWP30P140LVT U1524 ( .A1(n1253), .A2(i_data_bus[793]), .B1(n1266), 
        .B2(i_data_bus[377]), .ZN(n1119) );
  AOI22D1BWP30P140LVT U1525 ( .A1(n1254), .A2(i_data_bus[761]), .B1(n1267), 
        .B2(i_data_bus[473]), .ZN(n1118) );
  AOI22D1BWP30P140LVT U1526 ( .A1(n1263), .A2(i_data_bus[153]), .B1(n1246), 
        .B2(i_data_bus[281]), .ZN(n1117) );
  ND4D1BWP30P140LVT U1527 ( .A1(n1120), .A2(n1119), .A3(n1118), .A4(n1117), 
        .ZN(n1126) );
  AOI22D1BWP30P140LVT U1528 ( .A1(n1257), .A2(i_data_bus[409]), .B1(n1258), 
        .B2(i_data_bus[217]), .ZN(n1124) );
  AOI22D1BWP30P140LVT U1529 ( .A1(n617), .A2(i_data_bus[889]), .B1(n1244), 
        .B2(i_data_bus[313]), .ZN(n1123) );
  AOI22D1BWP30P140LVT U1530 ( .A1(n1247), .A2(i_data_bus[505]), .B1(n600), 
        .B2(i_data_bus[857]), .ZN(n1122) );
  AOI22D1BWP30P140LVT U1531 ( .A1(n1245), .A2(i_data_bus[441]), .B1(n1269), 
        .B2(i_data_bus[249]), .ZN(n1121) );
  ND4D1BWP30P140LVT U1532 ( .A1(n1124), .A2(n1123), .A3(n1122), .A4(n1121), 
        .ZN(n1125) );
  OR4D1BWP30P140LVT U1533 ( .A1(n1128), .A2(n1127), .A3(n1126), .A4(n1125), 
        .Z(o_data_bus[57]) );
  AOI22D1BWP30P140LVT U1534 ( .A1(n117), .A2(i_data_bus[122]), .B1(n1234), 
        .B2(i_data_bus[602]), .ZN(n1132) );
  AOI22D1BWP30P140LVT U1535 ( .A1(n1230), .A2(i_data_bus[1018]), .B1(n1229), 
        .B2(i_data_bus[90]), .ZN(n1131) );
  AOI22D1BWP30P140LVT U1536 ( .A1(n1242), .A2(i_data_bus[954]), .B1(n1231), 
        .B2(i_data_bus[986]), .ZN(n1130) );
  ND4D1BWP30P140LVT U1537 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1129), 
        .ZN(n1148) );
  AOI22D1BWP30P140LVT U1538 ( .A1(n1233), .A2(i_data_bus[570]), .B1(n1240), 
        .B2(i_data_bus[634]), .ZN(n1136) );
  AOI22D1BWP30P140LVT U1539 ( .A1(n103), .A2(i_data_bus[58]), .B1(n25), .B2(
        i_data_bus[26]), .ZN(n1135) );
  AOI22D1BWP30P140LVT U1540 ( .A1(n1245), .A2(i_data_bus[442]), .B1(n1258), 
        .B2(i_data_bus[218]), .ZN(n1134) );
  AOI22D1BWP30P140LVT U1541 ( .A1(n617), .A2(i_data_bus[890]), .B1(n1256), 
        .B2(i_data_bus[826]), .ZN(n1133) );
  ND4D1BWP30P140LVT U1542 ( .A1(n1136), .A2(n1135), .A3(n1134), .A4(n1133), 
        .ZN(n1147) );
  AOI22D1BWP30P140LVT U1543 ( .A1(n600), .A2(i_data_bus[858]), .B1(n1244), 
        .B2(i_data_bus[314]), .ZN(n1140) );
  AOI22D1BWP30P140LVT U1544 ( .A1(n1264), .A2(i_data_bus[698]), .B1(n1268), 
        .B2(i_data_bus[346]), .ZN(n1139) );
  AOI22D1BWP30P140LVT U1545 ( .A1(n1265), .A2(i_data_bus[186]), .B1(n1246), 
        .B2(i_data_bus[282]), .ZN(n1138) );
  AOI22D1BWP30P140LVT U1546 ( .A1(n1254), .A2(i_data_bus[762]), .B1(n1253), 
        .B2(i_data_bus[794]), .ZN(n1137) );
  ND4D1BWP30P140LVT U1547 ( .A1(n1140), .A2(n1139), .A3(n1138), .A4(n1137), 
        .ZN(n1146) );
  AOI22D1BWP30P140LVT U1548 ( .A1(n1247), .A2(i_data_bus[506]), .B1(n1269), 
        .B2(i_data_bus[250]), .ZN(n1144) );
  AOI22D1BWP30P140LVT U1549 ( .A1(n1257), .A2(i_data_bus[410]), .B1(n1255), 
        .B2(i_data_bus[666]), .ZN(n1143) );
  AOI22D1BWP30P140LVT U1550 ( .A1(n1263), .A2(i_data_bus[154]), .B1(n1252), 
        .B2(i_data_bus[730]), .ZN(n1142) );
  AOI22D1BWP30P140LVT U1551 ( .A1(n1267), .A2(i_data_bus[474]), .B1(n1266), 
        .B2(i_data_bus[378]), .ZN(n1141) );
  ND4D1BWP30P140LVT U1552 ( .A1(n1144), .A2(n1143), .A3(n1142), .A4(n1141), 
        .ZN(n1145) );
  OR4D1BWP30P140LVT U1553 ( .A1(n1148), .A2(n1147), .A3(n1146), .A4(n1145), 
        .Z(o_data_bus[58]) );
  AOI22D1BWP30P140LVT U1554 ( .A1(n117), .A2(i_data_bus[123]), .B1(n1231), 
        .B2(i_data_bus[987]), .ZN(n1152) );
  AOI22D1BWP30P140LVT U1555 ( .A1(n1230), .A2(i_data_bus[1019]), .B1(n1233), 
        .B2(i_data_bus[571]), .ZN(n1151) );
  AOI22D1BWP30P140LVT U1556 ( .A1(n1241), .A2(i_data_bus[539]), .B1(n1234), 
        .B2(i_data_bus[603]), .ZN(n1150) );
  AOI22D1BWP30P140LVT U1557 ( .A1(n1229), .A2(i_data_bus[91]), .B1(n1240), 
        .B2(i_data_bus[635]), .ZN(n1149) );
  ND4D1BWP30P140LVT U1558 ( .A1(n1152), .A2(n1151), .A3(n1150), .A4(n1149), 
        .ZN(n1168) );
  AOI22D1BWP30P140LVT U1559 ( .A1(n25), .A2(i_data_bus[27]), .B1(n594), .B2(
        i_data_bus[923]), .ZN(n1156) );
  AOI22D1BWP30P140LVT U1560 ( .A1(n103), .A2(i_data_bus[59]), .B1(n1242), .B2(
        i_data_bus[955]), .ZN(n1155) );
  AOI22D1BWP30P140LVT U1561 ( .A1(n1257), .A2(i_data_bus[411]), .B1(n1247), 
        .B2(i_data_bus[507]), .ZN(n1154) );
  AOI22D1BWP30P140LVT U1562 ( .A1(n1252), .A2(i_data_bus[731]), .B1(n1256), 
        .B2(i_data_bus[827]), .ZN(n1153) );
  ND4D1BWP30P140LVT U1563 ( .A1(n1156), .A2(n1155), .A3(n1154), .A4(n1153), 
        .ZN(n1167) );
  AOI22D1BWP30P140LVT U1564 ( .A1(n1245), .A2(i_data_bus[443]), .B1(n1263), 
        .B2(i_data_bus[155]), .ZN(n1160) );
  AOI22D1BWP30P140LVT U1565 ( .A1(n617), .A2(i_data_bus[891]), .B1(n1244), 
        .B2(i_data_bus[315]), .ZN(n1159) );
  AOI22D1BWP30P140LVT U1566 ( .A1(n1266), .A2(i_data_bus[379]), .B1(n1258), 
        .B2(i_data_bus[219]), .ZN(n1158) );
  AOI22D1BWP30P140LVT U1567 ( .A1(n1269), .A2(i_data_bus[251]), .B1(n1246), 
        .B2(i_data_bus[283]), .ZN(n1157) );
  ND4D1BWP30P140LVT U1568 ( .A1(n1160), .A2(n1159), .A3(n1158), .A4(n1157), 
        .ZN(n1166) );
  AOI22D1BWP30P140LVT U1569 ( .A1(n1254), .A2(i_data_bus[763]), .B1(n1253), 
        .B2(i_data_bus[795]), .ZN(n1164) );
  AOI22D1BWP30P140LVT U1570 ( .A1(n1255), .A2(i_data_bus[667]), .B1(n1267), 
        .B2(i_data_bus[475]), .ZN(n1163) );
  AOI22D1BWP30P140LVT U1571 ( .A1(n600), .A2(i_data_bus[859]), .B1(n1268), 
        .B2(i_data_bus[347]), .ZN(n1162) );
  AOI22D1BWP30P140LVT U1572 ( .A1(n1265), .A2(i_data_bus[187]), .B1(n1264), 
        .B2(i_data_bus[699]), .ZN(n1161) );
  ND4D1BWP30P140LVT U1573 ( .A1(n1164), .A2(n1163), .A3(n1162), .A4(n1161), 
        .ZN(n1165) );
  OR4D1BWP30P140LVT U1574 ( .A1(n1168), .A2(n1167), .A3(n1166), .A4(n1165), 
        .Z(o_data_bus[59]) );
  AOI22D1BWP30P140LVT U1575 ( .A1(n1242), .A2(i_data_bus[956]), .B1(n594), 
        .B2(i_data_bus[924]), .ZN(n1171) );
  AOI22D1BWP30P140LVT U1576 ( .A1(n1234), .A2(i_data_bus[604]), .B1(n1240), 
        .B2(i_data_bus[636]), .ZN(n1170) );
  AOI22D1BWP30P140LVT U1577 ( .A1(n117), .A2(i_data_bus[124]), .B1(n1229), 
        .B2(i_data_bus[92]), .ZN(n1169) );
  ND4D1BWP30P140LVT U1578 ( .A1(n1171), .A2(n1172), .A3(n1170), .A4(n1169), 
        .ZN(n1188) );
  AOI22D1BWP30P140LVT U1579 ( .A1(n1233), .A2(i_data_bus[572]), .B1(n25), .B2(
        i_data_bus[28]), .ZN(n1176) );
  AOI22D1BWP30P140LVT U1580 ( .A1(n1230), .A2(i_data_bus[1020]), .B1(n103), 
        .B2(i_data_bus[60]), .ZN(n1175) );
  AOI22D1BWP30P140LVT U1581 ( .A1(n1266), .A2(i_data_bus[380]), .B1(n1268), 
        .B2(i_data_bus[348]), .ZN(n1174) );
  AOI22D1BWP30P140LVT U1582 ( .A1(n1245), .A2(i_data_bus[444]), .B1(n1253), 
        .B2(i_data_bus[796]), .ZN(n1173) );
  ND4D1BWP30P140LVT U1583 ( .A1(n1176), .A2(n1175), .A3(n1174), .A4(n1173), 
        .ZN(n1187) );
  AOI22D1BWP30P140LVT U1584 ( .A1(n1252), .A2(i_data_bus[732]), .B1(n1269), 
        .B2(i_data_bus[252]), .ZN(n1180) );
  AOI22D1BWP30P140LVT U1585 ( .A1(n1247), .A2(i_data_bus[508]), .B1(n617), 
        .B2(i_data_bus[892]), .ZN(n1179) );
  AOI22D1BWP30P140LVT U1586 ( .A1(n1263), .A2(i_data_bus[156]), .B1(n1256), 
        .B2(i_data_bus[828]), .ZN(n1178) );
  AOI22D1BWP30P140LVT U1587 ( .A1(n1257), .A2(i_data_bus[412]), .B1(n1258), 
        .B2(i_data_bus[220]), .ZN(n1177) );
  ND4D1BWP30P140LVT U1588 ( .A1(n1180), .A2(n1179), .A3(n1178), .A4(n1177), 
        .ZN(n1186) );
  AOI22D1BWP30P140LVT U1589 ( .A1(n1255), .A2(i_data_bus[668]), .B1(n1254), 
        .B2(i_data_bus[764]), .ZN(n1184) );
  AOI22D1BWP30P140LVT U1590 ( .A1(n600), .A2(i_data_bus[860]), .B1(n1265), 
        .B2(i_data_bus[188]), .ZN(n1183) );
  AOI22D1BWP30P140LVT U1591 ( .A1(n1267), .A2(i_data_bus[476]), .B1(n1264), 
        .B2(i_data_bus[700]), .ZN(n1182) );
  AOI22D1BWP30P140LVT U1592 ( .A1(n1244), .A2(i_data_bus[316]), .B1(n1246), 
        .B2(i_data_bus[284]), .ZN(n1181) );
  ND4D1BWP30P140LVT U1593 ( .A1(n1184), .A2(n1183), .A3(n1182), .A4(n1181), 
        .ZN(n1185) );
  OR4D1BWP30P140LVT U1594 ( .A1(n1188), .A2(n1187), .A3(n1186), .A4(n1185), 
        .Z(o_data_bus[60]) );
  AOI22D1BWP30P140LVT U1595 ( .A1(n1242), .A2(i_data_bus[957]), .B1(n594), 
        .B2(i_data_bus[925]), .ZN(n1192) );
  AOI22D1BWP30P140LVT U1596 ( .A1(n1233), .A2(i_data_bus[573]), .B1(n25), .B2(
        i_data_bus[29]), .ZN(n1191) );
  AOI22D1BWP30P140LVT U1597 ( .A1(n1231), .A2(i_data_bus[989]), .B1(n1240), 
        .B2(i_data_bus[637]), .ZN(n1190) );
  AOI22D1BWP30P140LVT U1598 ( .A1(n1230), .A2(i_data_bus[1021]), .B1(n117), 
        .B2(i_data_bus[125]), .ZN(n1189) );
  ND4D1BWP30P140LVT U1599 ( .A1(n1192), .A2(n1191), .A3(n1190), .A4(n1189), 
        .ZN(n1208) );
  AOI22D1BWP30P140LVT U1600 ( .A1(n1241), .A2(i_data_bus[541]), .B1(n1234), 
        .B2(i_data_bus[605]), .ZN(n1196) );
  AOI22D1BWP30P140LVT U1601 ( .A1(n1232), .A2(i_data_bus[61]), .B1(n1229), 
        .B2(i_data_bus[93]), .ZN(n1195) );
  AOI22D1BWP30P140LVT U1602 ( .A1(n1263), .A2(i_data_bus[157]), .B1(n1264), 
        .B2(i_data_bus[701]), .ZN(n1194) );
  AOI22D1BWP30P140LVT U1603 ( .A1(n1245), .A2(i_data_bus[445]), .B1(n1255), 
        .B2(i_data_bus[669]), .ZN(n1193) );
  ND4D1BWP30P140LVT U1604 ( .A1(n1196), .A2(n1195), .A3(n1194), .A4(n1193), 
        .ZN(n1207) );
  AOI22D1BWP30P140LVT U1605 ( .A1(n1254), .A2(i_data_bus[765]), .B1(n1244), 
        .B2(i_data_bus[317]), .ZN(n1200) );
  AOI22D1BWP30P140LVT U1606 ( .A1(n1247), .A2(i_data_bus[509]), .B1(n1265), 
        .B2(i_data_bus[189]), .ZN(n1199) );
  AOI22D1BWP30P140LVT U1607 ( .A1(n1253), .A2(i_data_bus[797]), .B1(n1268), 
        .B2(i_data_bus[349]), .ZN(n1198) );
  AOI22D1BWP30P140LVT U1608 ( .A1(n1267), .A2(i_data_bus[477]), .B1(n1252), 
        .B2(i_data_bus[733]), .ZN(n1197) );
  ND4D1BWP30P140LVT U1609 ( .A1(n1200), .A2(n1199), .A3(n1198), .A4(n1197), 
        .ZN(n1206) );
  AOI22D1BWP30P140LVT U1610 ( .A1(n1257), .A2(i_data_bus[413]), .B1(n1266), 
        .B2(i_data_bus[381]), .ZN(n1204) );
  AOI22D1BWP30P140LVT U1611 ( .A1(n1269), .A2(i_data_bus[253]), .B1(n1246), 
        .B2(i_data_bus[285]), .ZN(n1203) );
  AOI22D1BWP30P140LVT U1612 ( .A1(n600), .A2(i_data_bus[861]), .B1(n1256), 
        .B2(i_data_bus[829]), .ZN(n1202) );
  AOI22D1BWP30P140LVT U1613 ( .A1(n1258), .A2(i_data_bus[221]), .B1(n617), 
        .B2(i_data_bus[893]), .ZN(n1201) );
  ND4D1BWP30P140LVT U1614 ( .A1(n1204), .A2(n1203), .A3(n1202), .A4(n1201), 
        .ZN(n1205) );
  OR4D1BWP30P140LVT U1615 ( .A1(n1208), .A2(n1207), .A3(n1206), .A4(n1205), 
        .Z(o_data_bus[61]) );
  AOI22D1BWP30P140LVT U1616 ( .A1(n1232), .A2(i_data_bus[62]), .B1(n594), .B2(
        i_data_bus[926]), .ZN(n1212) );
  AOI22D1BWP30P140LVT U1617 ( .A1(n1233), .A2(i_data_bus[574]), .B1(n117), 
        .B2(i_data_bus[126]), .ZN(n1210) );
  AOI22D1BWP30P140LVT U1618 ( .A1(n1230), .A2(i_data_bus[1022]), .B1(n1231), 
        .B2(i_data_bus[990]), .ZN(n1209) );
  ND4D1BWP30P140LVT U1619 ( .A1(n1212), .A2(n1209), .A3(n1211), .A4(n1210), 
        .ZN(n1228) );
  AOI22D1BWP30P140LVT U1620 ( .A1(n25), .A2(i_data_bus[30]), .B1(n1229), .B2(
        i_data_bus[94]), .ZN(n1216) );
  AOI22D1BWP30P140LVT U1621 ( .A1(n1234), .A2(i_data_bus[606]), .B1(n1240), 
        .B2(i_data_bus[638]), .ZN(n1215) );
  AOI22D1BWP30P140LVT U1622 ( .A1(n1255), .A2(i_data_bus[670]), .B1(n1258), 
        .B2(i_data_bus[222]), .ZN(n1214) );
  AOI22D1BWP30P140LVT U1623 ( .A1(n1245), .A2(i_data_bus[446]), .B1(n1268), 
        .B2(i_data_bus[350]), .ZN(n1213) );
  ND4D1BWP30P140LVT U1624 ( .A1(n1216), .A2(n1215), .A3(n1214), .A4(n1213), 
        .ZN(n1227) );
  AOI22D1BWP30P140LVT U1625 ( .A1(n600), .A2(i_data_bus[862]), .B1(n1244), 
        .B2(i_data_bus[318]), .ZN(n1220) );
  AOI22D1BWP30P140LVT U1626 ( .A1(n1253), .A2(i_data_bus[798]), .B1(n1246), 
        .B2(i_data_bus[286]), .ZN(n1219) );
  AOI22D1BWP30P140LVT U1627 ( .A1(n1254), .A2(i_data_bus[766]), .B1(n1265), 
        .B2(i_data_bus[190]), .ZN(n1218) );
  AOI22D1BWP30P140LVT U1628 ( .A1(n1269), .A2(i_data_bus[254]), .B1(n1256), 
        .B2(i_data_bus[830]), .ZN(n1217) );
  ND4D1BWP30P140LVT U1629 ( .A1(n1220), .A2(n1219), .A3(n1218), .A4(n1217), 
        .ZN(n1226) );
  AOI22D1BWP30P140LVT U1630 ( .A1(n1257), .A2(i_data_bus[414]), .B1(n1267), 
        .B2(i_data_bus[478]), .ZN(n1224) );
  AOI22D1BWP30P140LVT U1631 ( .A1(n1247), .A2(i_data_bus[510]), .B1(n1264), 
        .B2(i_data_bus[702]), .ZN(n1223) );
  AOI22D1BWP30P140LVT U1632 ( .A1(n1266), .A2(i_data_bus[382]), .B1(n1252), 
        .B2(i_data_bus[734]), .ZN(n1222) );
  AOI22D1BWP30P140LVT U1633 ( .A1(n1263), .A2(i_data_bus[158]), .B1(n617), 
        .B2(i_data_bus[894]), .ZN(n1221) );
  ND4D1BWP30P140LVT U1634 ( .A1(n1224), .A2(n1223), .A3(n1222), .A4(n1221), 
        .ZN(n1225) );
  OR4D1BWP30P140LVT U1635 ( .A1(n1225), .A2(n1227), .A3(n1226), .A4(n1228), 
        .Z(o_data_bus[62]) );
  AOI22D1BWP30P140LVT U1636 ( .A1(n1230), .A2(i_data_bus[1023]), .B1(n1229), 
        .B2(i_data_bus[95]), .ZN(n1239) );
  AOI22D1BWP30P140LVT U1637 ( .A1(n103), .A2(i_data_bus[63]), .B1(n1231), .B2(
        i_data_bus[991]), .ZN(n1238) );
  AOI22D1BWP30P140LVT U1638 ( .A1(n25), .A2(i_data_bus[31]), .B1(n1234), .B2(
        i_data_bus[607]), .ZN(n1236) );
  ND4D1BWP30P140LVT U1639 ( .A1(n1238), .A2(n1239), .A3(n1237), .A4(n1236), 
        .ZN(n1277) );
  AOI22D1BWP30P140LVT U1640 ( .A1(n1241), .A2(i_data_bus[543]), .B1(n1240), 
        .B2(i_data_bus[639]), .ZN(n1251) );
  AOI22D1BWP30P140LVT U1641 ( .A1(n117), .A2(i_data_bus[127]), .B1(n1242), 
        .B2(i_data_bus[959]), .ZN(n1250) );
  AOI22D1BWP30P140LVT U1642 ( .A1(n1245), .A2(i_data_bus[447]), .B1(n1244), 
        .B2(i_data_bus[319]), .ZN(n1249) );
  AOI22D1BWP30P140LVT U1643 ( .A1(n1247), .A2(i_data_bus[511]), .B1(n1246), 
        .B2(i_data_bus[287]), .ZN(n1248) );
  ND4D1BWP30P140LVT U1644 ( .A1(n1251), .A2(n1250), .A3(n1249), .A4(n1248), 
        .ZN(n1276) );
  AOI22D1BWP30P140LVT U1645 ( .A1(n1253), .A2(i_data_bus[799]), .B1(n1252), 
        .B2(i_data_bus[735]), .ZN(n1262) );
  AOI22D1BWP30P140LVT U1646 ( .A1(n1255), .A2(i_data_bus[671]), .B1(n1254), 
        .B2(i_data_bus[767]), .ZN(n1261) );
  AOI22D1BWP30P140LVT U1647 ( .A1(n1257), .A2(i_data_bus[415]), .B1(n1256), 
        .B2(i_data_bus[831]), .ZN(n1260) );
  AOI22D1BWP30P140LVT U1648 ( .A1(n600), .A2(i_data_bus[863]), .B1(n1258), 
        .B2(i_data_bus[223]), .ZN(n1259) );
  ND4D1BWP30P140LVT U1649 ( .A1(n1262), .A2(n1261), .A3(n1260), .A4(n1259), 
        .ZN(n1275) );
  AOI22D1BWP30P140LVT U1650 ( .A1(n1263), .A2(i_data_bus[159]), .B1(n617), 
        .B2(i_data_bus[895]), .ZN(n1273) );
  AOI22D1BWP30P140LVT U1651 ( .A1(n1265), .A2(i_data_bus[191]), .B1(n1264), 
        .B2(i_data_bus[703]), .ZN(n1272) );
  AOI22D1BWP30P140LVT U1652 ( .A1(n1267), .A2(i_data_bus[479]), .B1(n1266), 
        .B2(i_data_bus[383]), .ZN(n1271) );
  AOI22D1BWP30P140LVT U1653 ( .A1(n1269), .A2(i_data_bus[255]), .B1(n1268), 
        .B2(i_data_bus[351]), .ZN(n1270) );
  ND4D1BWP30P140LVT U1654 ( .A1(n1273), .A2(n1272), .A3(n1271), .A4(n1270), 
        .ZN(n1274) );
  OR4D1BWP30P140LVT U1655 ( .A1(n1277), .A2(n1276), .A3(n1275), .A4(n1274), 
        .Z(o_data_bus[63]) );
  INR3D2BWP30P140LVT U1656 ( .A1(i_cmd[107]), .B1(n4085), .B2(n1287), .ZN(
        n1921) );
  AOI22D1BWP30P140LVT U1657 ( .A1(i_data_bus[608]), .A2(n1910), .B1(
        i_data_bus[416]), .B2(n1921), .ZN(n1283) );
  INR3D2BWP30P140LVT U1658 ( .A1(i_cmd[83]), .B1(n4084), .B2(n1295), .ZN(n1913) );
  AOI22D1BWP30P140LVT U1659 ( .A1(i_data_bus[64]), .A2(n1925), .B1(
        i_data_bus[320]), .B2(n1913), .ZN(n1282) );
  AOI22D1BWP30P140LVT U1660 ( .A1(i_data_bus[544]), .A2(n1924), .B1(
        i_data_bus[0]), .B2(n2), .ZN(n1281) );
  INR3D2BWP30P140LVT U1661 ( .A1(i_cmd[115]), .B1(n4083), .B2(n1287), .ZN(
        n1933) );
  AOI22D1BWP30P140LVT U1662 ( .A1(i_data_bus[384]), .A2(n1279), .B1(
        i_data_bus[448]), .B2(n1933), .ZN(n1280) );
  ND4D1BWP30P140LVT U1663 ( .A1(n1283), .A2(n1282), .A3(n1281), .A4(n1280), 
        .ZN(n1316) );
  INR3D2BWP30P140LVT U1664 ( .A1(i_cmd[75]), .B1(n4095), .B2(n1295), .ZN(n1922) );
  AOI22D1BWP30P140LVT U1665 ( .A1(i_data_bus[224]), .A2(n1911), .B1(
        i_data_bus[288]), .B2(n1922), .ZN(n1291) );
  INVD1BWP30P140LVT U1666 ( .I(i_cmd[131]), .ZN(n1284) );
  AOI22D1BWP30P140LVT U1667 ( .A1(i_data_bus[512]), .A2(n1927), .B1(
        i_data_bus[960]), .B2(n1923), .ZN(n1290) );
  INR3D2BWP30P140LVT U1668 ( .A1(i_cmd[123]), .B1(n4110), .B2(n1287), .ZN(
        n1932) );
  AOI22D1BWP30P140LVT U1669 ( .A1(i_data_bus[992]), .A2(n1934), .B1(
        i_data_bus[480]), .B2(n1932), .ZN(n1289) );
  INR3D2BWP30P140LVT U1670 ( .A1(n1294), .B1(n5493), .B2(n133), .ZN(n1935) );
  AOI22D1BWP30P140LVT U1671 ( .A1(i_data_bus[128]), .A2(n1935), .B1(
        i_data_bus[192]), .B2(n1916), .ZN(n1288) );
  ND4D1BWP30P140LVT U1672 ( .A1(n1291), .A2(n1290), .A3(n1289), .A4(n1288), 
        .ZN(n1315) );
  INVD1BWP30P140LVT U1673 ( .I(i_cmd[67]), .ZN(n1292) );
  AOI22D1BWP30P140LVT U1674 ( .A1(i_data_bus[96]), .A2(n1936), .B1(
        i_data_bus[256]), .B2(n1293), .ZN(n1304) );
  INR3D2BWP30P140LVT U1675 ( .A1(i_cmd[91]), .B1(n4074), .B2(n1295), .ZN(n1926) );
  AOI22D1BWP30P140LVT U1676 ( .A1(i_data_bus[160]), .A2(n1915), .B1(
        i_data_bus[352]), .B2(n1926), .ZN(n1303) );
  AOI22D1BWP30P140LVT U1677 ( .A1(i_data_bus[576]), .A2(n1912), .B1(
        i_data_bus[896]), .B2(n128), .ZN(n1302) );
  AOI22D1BWP30P140LVT U1678 ( .A1(i_data_bus[32]), .A2(n1914), .B1(
        i_data_bus[928]), .B2(n127), .ZN(n1301) );
  ND4D1BWP30P140LVT U1679 ( .A1(n1304), .A2(n1303), .A3(n1302), .A4(n1301), 
        .ZN(n1314) );
  INR3D2BWP30P140LVT U1680 ( .A1(i_cmd[211]), .B1(n5461), .B2(n1306), .ZN(
        n1948) );
  INVD1BWP30P140LVT U1681 ( .I(i_cmd[163]), .ZN(n1305) );
  AOI22D1BWP30P140LVT U1682 ( .A1(i_data_bus[832]), .A2(n1948), .B1(
        i_data_bus[640]), .B2(n1944), .ZN(n1312) );
  INR3D2BWP30P140LVT U1683 ( .A1(i_cmd[179]), .B1(n5448), .B2(n1308), .ZN(
        n1942) );
  INR3D2BWP30P140LVT U1684 ( .A1(i_cmd[219]), .B1(n5457), .B2(n1306), .ZN(
        n1941) );
  AOI22D1BWP30P140LVT U1685 ( .A1(i_data_bus[704]), .A2(n1942), .B1(
        i_data_bus[864]), .B2(n1941), .ZN(n1311) );
  INR3D2BWP30P140LVT U1686 ( .A1(i_cmd[187]), .B1(n5458), .B2(n1308), .ZN(
        n1945) );
  INR3D2BWP30P140LVT U1687 ( .A1(i_cmd[203]), .B1(n5459), .B2(n1306), .ZN(
        n1943) );
  AOI22D1BWP30P140LVT U1688 ( .A1(i_data_bus[736]), .A2(n1945), .B1(
        i_data_bus[800]), .B2(n1943), .ZN(n1310) );
  INVD1BWP30P140LVT U1689 ( .I(i_cmd[195]), .ZN(n1307) );
  NR3D1P5BWP30P140LVT U1690 ( .A1(n5444), .A2(n1307), .A3(n1306), .ZN(n1946)
         );
  INR3D2BWP30P140LVT U1691 ( .A1(i_cmd[171]), .B1(n5463), .B2(n1308), .ZN(
        n1947) );
  AOI22D1BWP30P140LVT U1692 ( .A1(i_data_bus[768]), .A2(n1946), .B1(
        i_data_bus[672]), .B2(n1947), .ZN(n1309) );
  ND4D1BWP30P140LVT U1693 ( .A1(n1312), .A2(n1311), .A3(n1310), .A4(n1309), 
        .ZN(n1313) );
  OR4D1BWP30P140LVT U1694 ( .A1(n1316), .A2(n1315), .A3(n1314), .A4(n1313), 
        .Z(o_data_bus[96]) );
  AOI22D1BWP30P140LVT U1695 ( .A1(i_data_bus[385]), .A2(n1279), .B1(
        i_data_bus[225]), .B2(n1911), .ZN(n1320) );
  AOI22D1BWP30P140LVT U1696 ( .A1(i_data_bus[65]), .A2(n1925), .B1(
        i_data_bus[513]), .B2(n1927), .ZN(n1319) );
  AOI22D1BWP30P140LVT U1697 ( .A1(i_data_bus[929]), .A2(n127), .B1(
        i_data_bus[129]), .B2(n1935), .ZN(n1318) );
  AOI22D1BWP30P140LVT U1698 ( .A1(i_data_bus[33]), .A2(n1914), .B1(
        i_data_bus[161]), .B2(n1915), .ZN(n1317) );
  ND4D1BWP30P140LVT U1699 ( .A1(n1320), .A2(n1319), .A3(n1318), .A4(n1317), 
        .ZN(n1336) );
  AOI22D1BWP30P140LVT U1700 ( .A1(i_data_bus[97]), .A2(n1936), .B1(
        i_data_bus[1]), .B2(n2), .ZN(n1324) );
  AOI22D1BWP30P140LVT U1701 ( .A1(i_data_bus[257]), .A2(n1293), .B1(
        i_data_bus[449]), .B2(n1933), .ZN(n1323) );
  AOI22D1BWP30P140LVT U1702 ( .A1(i_data_bus[897]), .A2(n128), .B1(
        i_data_bus[481]), .B2(n1932), .ZN(n1322) );
  AOI22D1BWP30P140LVT U1703 ( .A1(i_data_bus[289]), .A2(n1922), .B1(
        i_data_bus[321]), .B2(n1913), .ZN(n1321) );
  ND4D1BWP30P140LVT U1704 ( .A1(n1324), .A2(n1323), .A3(n1322), .A4(n1321), 
        .ZN(n1335) );
  AOI22D1BWP30P140LVT U1705 ( .A1(i_data_bus[993]), .A2(n1934), .B1(
        i_data_bus[609]), .B2(n1910), .ZN(n1328) );
  AOI22D1BWP30P140LVT U1706 ( .A1(i_data_bus[961]), .A2(n1923), .B1(
        i_data_bus[193]), .B2(n1916), .ZN(n1327) );
  AOI22D1BWP30P140LVT U1707 ( .A1(i_data_bus[577]), .A2(n1912), .B1(
        i_data_bus[417]), .B2(n1921), .ZN(n1326) );
  AOI22D1BWP30P140LVT U1708 ( .A1(i_data_bus[545]), .A2(n1924), .B1(
        i_data_bus[353]), .B2(n1926), .ZN(n1325) );
  ND4D1BWP30P140LVT U1709 ( .A1(n1328), .A2(n1327), .A3(n1326), .A4(n1325), 
        .ZN(n1334) );
  AOI22D1BWP30P140LVT U1710 ( .A1(i_data_bus[769]), .A2(n1946), .B1(
        i_data_bus[737]), .B2(n1945), .ZN(n1332) );
  AOI22D1BWP30P140LVT U1711 ( .A1(i_data_bus[705]), .A2(n1942), .B1(
        i_data_bus[641]), .B2(n1944), .ZN(n1331) );
  AOI22D1BWP30P140LVT U1712 ( .A1(i_data_bus[673]), .A2(n1947), .B1(
        i_data_bus[865]), .B2(n1941), .ZN(n1330) );
  AOI22D1BWP30P140LVT U1713 ( .A1(i_data_bus[801]), .A2(n1943), .B1(
        i_data_bus[833]), .B2(n1948), .ZN(n1329) );
  ND4D1BWP30P140LVT U1714 ( .A1(n1332), .A2(n1331), .A3(n1330), .A4(n1329), 
        .ZN(n1333) );
  OR4D1BWP30P140LVT U1715 ( .A1(n1336), .A2(n1335), .A3(n1334), .A4(n1333), 
        .Z(o_data_bus[97]) );
  AOI22D1BWP30P140LVT U1716 ( .A1(i_data_bus[546]), .A2(n1924), .B1(
        i_data_bus[226]), .B2(n1911), .ZN(n1340) );
  AOI22D1BWP30P140LVT U1717 ( .A1(i_data_bus[578]), .A2(n1912), .B1(
        i_data_bus[130]), .B2(n1935), .ZN(n1339) );
  AOI22D1BWP30P140LVT U1718 ( .A1(i_data_bus[2]), .A2(n2), .B1(i_data_bus[194]), .B2(n1916), .ZN(n1338) );
  AOI22D1BWP30P140LVT U1719 ( .A1(i_data_bus[162]), .A2(n1915), .B1(
        i_data_bus[450]), .B2(n1933), .ZN(n1337) );
  ND4D1BWP30P140LVT U1720 ( .A1(n1340), .A2(n1339), .A3(n1338), .A4(n1337), 
        .ZN(n1356) );
  AOI22D1BWP30P140LVT U1721 ( .A1(i_data_bus[482]), .A2(n1932), .B1(
        i_data_bus[258]), .B2(n1293), .ZN(n1344) );
  AOI22D1BWP30P140LVT U1722 ( .A1(i_data_bus[994]), .A2(n1934), .B1(
        i_data_bus[354]), .B2(n1926), .ZN(n1343) );
  AOI22D1BWP30P140LVT U1723 ( .A1(i_data_bus[98]), .A2(n1936), .B1(
        i_data_bus[418]), .B2(n1921), .ZN(n1342) );
  AOI22D1BWP30P140LVT U1724 ( .A1(i_data_bus[930]), .A2(n127), .B1(
        i_data_bus[290]), .B2(n1922), .ZN(n1341) );
  ND4D1BWP30P140LVT U1725 ( .A1(n1344), .A2(n1343), .A3(n1342), .A4(n1341), 
        .ZN(n1355) );
  AOI22D1BWP30P140LVT U1726 ( .A1(i_data_bus[898]), .A2(n128), .B1(
        i_data_bus[514]), .B2(n1927), .ZN(n1348) );
  AOI22D1BWP30P140LVT U1727 ( .A1(i_data_bus[386]), .A2(n1279), .B1(
        i_data_bus[322]), .B2(n1913), .ZN(n1347) );
  AOI22D1BWP30P140LVT U1728 ( .A1(i_data_bus[66]), .A2(n1925), .B1(
        i_data_bus[610]), .B2(n1910), .ZN(n1346) );
  ND4D1BWP30P140LVT U1729 ( .A1(n1348), .A2(n1347), .A3(n1346), .A4(n1345), 
        .ZN(n1354) );
  AOI22D1BWP30P140LVT U1730 ( .A1(i_data_bus[834]), .A2(n1948), .B1(
        i_data_bus[642]), .B2(n1944), .ZN(n1352) );
  AOI22D1BWP30P140LVT U1731 ( .A1(i_data_bus[866]), .A2(n1941), .B1(
        i_data_bus[738]), .B2(n1945), .ZN(n1351) );
  AOI22D1BWP30P140LVT U1732 ( .A1(i_data_bus[674]), .A2(n1947), .B1(
        i_data_bus[706]), .B2(n1942), .ZN(n1350) );
  AOI22D1BWP30P140LVT U1733 ( .A1(i_data_bus[802]), .A2(n1943), .B1(
        i_data_bus[770]), .B2(n1946), .ZN(n1349) );
  ND4D1BWP30P140LVT U1734 ( .A1(n1352), .A2(n1351), .A3(n1350), .A4(n1349), 
        .ZN(n1353) );
  OR4D1BWP30P140LVT U1735 ( .A1(n1356), .A2(n1355), .A3(n1354), .A4(n1353), 
        .Z(o_data_bus[98]) );
  AOI22D1BWP30P140LVT U1736 ( .A1(i_data_bus[67]), .A2(n1925), .B1(
        i_data_bus[899]), .B2(n128), .ZN(n1360) );
  AOI22D1BWP30P140LVT U1737 ( .A1(i_data_bus[35]), .A2(n1914), .B1(
        i_data_bus[451]), .B2(n1933), .ZN(n1359) );
  AOI22D1BWP30P140LVT U1738 ( .A1(i_data_bus[963]), .A2(n1923), .B1(
        i_data_bus[163]), .B2(n1915), .ZN(n1358) );
  AOI22D1BWP30P140LVT U1739 ( .A1(i_data_bus[259]), .A2(n1293), .B1(
        i_data_bus[227]), .B2(n1911), .ZN(n1357) );
  ND4D1BWP30P140LVT U1740 ( .A1(n1360), .A2(n1359), .A3(n1358), .A4(n1357), 
        .ZN(n1376) );
  AOI22D1BWP30P140LVT U1741 ( .A1(i_data_bus[579]), .A2(n1912), .B1(
        i_data_bus[3]), .B2(n2), .ZN(n1364) );
  AOI22D1BWP30P140LVT U1742 ( .A1(i_data_bus[515]), .A2(n1927), .B1(
        i_data_bus[547]), .B2(n1924), .ZN(n1363) );
  AOI22D1BWP30P140LVT U1743 ( .A1(i_data_bus[995]), .A2(n1934), .B1(
        i_data_bus[483]), .B2(n1932), .ZN(n1362) );
  AOI22D1BWP30P140LVT U1744 ( .A1(i_data_bus[419]), .A2(n1921), .B1(
        i_data_bus[323]), .B2(n1913), .ZN(n1361) );
  ND4D1BWP30P140LVT U1745 ( .A1(n1364), .A2(n1363), .A3(n1362), .A4(n1361), 
        .ZN(n1375) );
  AOI22D1BWP30P140LVT U1746 ( .A1(i_data_bus[931]), .A2(n127), .B1(
        i_data_bus[355]), .B2(n1926), .ZN(n1368) );
  AOI22D1BWP30P140LVT U1747 ( .A1(i_data_bus[611]), .A2(n1910), .B1(
        i_data_bus[291]), .B2(n1922), .ZN(n1367) );
  AOI22D1BWP30P140LVT U1748 ( .A1(i_data_bus[387]), .A2(n1279), .B1(
        i_data_bus[195]), .B2(n1916), .ZN(n1366) );
  AOI22D1BWP30P140LVT U1749 ( .A1(i_data_bus[99]), .A2(n1936), .B1(
        i_data_bus[131]), .B2(n1935), .ZN(n1365) );
  ND4D1BWP30P140LVT U1750 ( .A1(n1368), .A2(n1367), .A3(n1366), .A4(n1365), 
        .ZN(n1374) );
  AOI22D1BWP30P140LVT U1751 ( .A1(i_data_bus[835]), .A2(n1948), .B1(
        i_data_bus[739]), .B2(n1945), .ZN(n1372) );
  AOI22D1BWP30P140LVT U1752 ( .A1(i_data_bus[771]), .A2(n1946), .B1(
        i_data_bus[803]), .B2(n1943), .ZN(n1371) );
  AOI22D1BWP30P140LVT U1753 ( .A1(i_data_bus[643]), .A2(n1944), .B1(
        i_data_bus[707]), .B2(n1942), .ZN(n1370) );
  AOI22D1BWP30P140LVT U1754 ( .A1(i_data_bus[675]), .A2(n1947), .B1(
        i_data_bus[867]), .B2(n1941), .ZN(n1369) );
  ND4D1BWP30P140LVT U1755 ( .A1(n1372), .A2(n1371), .A3(n1370), .A4(n1369), 
        .ZN(n1373) );
  OR4D1BWP30P140LVT U1756 ( .A1(n1376), .A2(n1375), .A3(n1374), .A4(n1373), 
        .Z(o_data_bus[99]) );
  AOI22D1BWP30P140LVT U1757 ( .A1(i_data_bus[900]), .A2(n128), .B1(
        i_data_bus[356]), .B2(n1926), .ZN(n1379) );
  AOI22D1BWP30P140LVT U1758 ( .A1(i_data_bus[996]), .A2(n1934), .B1(
        i_data_bus[484]), .B2(n1932), .ZN(n1377) );
  ND4D1BWP30P140LVT U1759 ( .A1(n1380), .A2(n1379), .A3(n1378), .A4(n1377), 
        .ZN(n1396) );
  AOI22D1BWP30P140LVT U1760 ( .A1(i_data_bus[516]), .A2(n1927), .B1(
        i_data_bus[420]), .B2(n1921), .ZN(n1384) );
  AOI22D1BWP30P140LVT U1761 ( .A1(i_data_bus[324]), .A2(n1913), .B1(
        i_data_bus[260]), .B2(n1293), .ZN(n1383) );
  AOI22D1BWP30P140LVT U1762 ( .A1(i_data_bus[932]), .A2(n127), .B1(
        i_data_bus[164]), .B2(n1915), .ZN(n1382) );
  AOI22D1BWP30P140LVT U1763 ( .A1(i_data_bus[100]), .A2(n1936), .B1(
        i_data_bus[196]), .B2(n1916), .ZN(n1381) );
  ND4D1BWP30P140LVT U1764 ( .A1(n1384), .A2(n1383), .A3(n1382), .A4(n1381), 
        .ZN(n1395) );
  AOI22D1BWP30P140LVT U1765 ( .A1(i_data_bus[228]), .A2(n1911), .B1(
        i_data_bus[452]), .B2(n1933), .ZN(n1388) );
  AOI22D1BWP30P140LVT U1766 ( .A1(i_data_bus[612]), .A2(n1910), .B1(
        i_data_bus[292]), .B2(n1922), .ZN(n1387) );
  AOI22D1BWP30P140LVT U1767 ( .A1(i_data_bus[4]), .A2(n2), .B1(i_data_bus[580]), .B2(n1912), .ZN(n1386) );
  AOI22D1BWP30P140LVT U1768 ( .A1(i_data_bus[132]), .A2(n1935), .B1(
        i_data_bus[388]), .B2(n1279), .ZN(n1385) );
  ND4D1BWP30P140LVT U1769 ( .A1(n1388), .A2(n1387), .A3(n1386), .A4(n1385), 
        .ZN(n1394) );
  AOI22D1BWP30P140LVT U1770 ( .A1(i_data_bus[740]), .A2(n1945), .B1(
        i_data_bus[772]), .B2(n1946), .ZN(n1392) );
  AOI22D1BWP30P140LVT U1771 ( .A1(i_data_bus[836]), .A2(n1948), .B1(
        i_data_bus[804]), .B2(n1943), .ZN(n1391) );
  AOI22D1BWP30P140LVT U1772 ( .A1(i_data_bus[708]), .A2(n1942), .B1(
        i_data_bus[644]), .B2(n1944), .ZN(n1390) );
  AOI22D1BWP30P140LVT U1773 ( .A1(i_data_bus[868]), .A2(n1941), .B1(
        i_data_bus[676]), .B2(n1947), .ZN(n1389) );
  ND4D1BWP30P140LVT U1774 ( .A1(n1392), .A2(n1391), .A3(n1390), .A4(n1389), 
        .ZN(n1393) );
  OR4D1BWP30P140LVT U1775 ( .A1(n1396), .A2(n1395), .A3(n1394), .A4(n1393), 
        .Z(o_data_bus[100]) );
  AOI22D1BWP30P140LVT U1776 ( .A1(i_data_bus[133]), .A2(n1935), .B1(
        i_data_bus[229]), .B2(n1911), .ZN(n1400) );
  AOI22D1BWP30P140LVT U1777 ( .A1(i_data_bus[933]), .A2(n127), .B1(
        i_data_bus[613]), .B2(n1910), .ZN(n1399) );
  AOI22D1BWP30P140LVT U1778 ( .A1(i_data_bus[997]), .A2(n1934), .B1(
        i_data_bus[261]), .B2(n1293), .ZN(n1398) );
  AOI22D1BWP30P140LVT U1779 ( .A1(i_data_bus[101]), .A2(n1936), .B1(
        i_data_bus[965]), .B2(n1923), .ZN(n1397) );
  ND4D1BWP30P140LVT U1780 ( .A1(n1400), .A2(n1399), .A3(n1398), .A4(n1397), 
        .ZN(n1416) );
  AOI22D1BWP30P140LVT U1781 ( .A1(i_data_bus[581]), .A2(n1912), .B1(
        i_data_bus[421]), .B2(n1921), .ZN(n1404) );
  AOI22D1BWP30P140LVT U1782 ( .A1(i_data_bus[197]), .A2(n1916), .B1(
        i_data_bus[453]), .B2(n1933), .ZN(n1403) );
  AOI22D1BWP30P140LVT U1783 ( .A1(i_data_bus[517]), .A2(n1927), .B1(
        i_data_bus[549]), .B2(n1924), .ZN(n1402) );
  AOI22D1BWP30P140LVT U1784 ( .A1(i_data_bus[485]), .A2(n1932), .B1(
        i_data_bus[293]), .B2(n1922), .ZN(n1401) );
  ND4D1BWP30P140LVT U1785 ( .A1(n1404), .A2(n1403), .A3(n1402), .A4(n1401), 
        .ZN(n1415) );
  AOI22D1BWP30P140LVT U1786 ( .A1(i_data_bus[69]), .A2(n1925), .B1(
        i_data_bus[357]), .B2(n1926), .ZN(n1408) );
  AOI22D1BWP30P140LVT U1787 ( .A1(i_data_bus[5]), .A2(n2), .B1(i_data_bus[325]), .B2(n1913), .ZN(n1407) );
  AOI22D1BWP30P140LVT U1788 ( .A1(i_data_bus[37]), .A2(n1914), .B1(
        i_data_bus[389]), .B2(n1279), .ZN(n1406) );
  AOI22D1BWP30P140LVT U1789 ( .A1(i_data_bus[901]), .A2(n128), .B1(
        i_data_bus[165]), .B2(n1915), .ZN(n1405) );
  ND4D1BWP30P140LVT U1790 ( .A1(n1408), .A2(n1407), .A3(n1406), .A4(n1405), 
        .ZN(n1414) );
  AOI22D1BWP30P140LVT U1791 ( .A1(i_data_bus[773]), .A2(n1946), .B1(
        i_data_bus[837]), .B2(n1948), .ZN(n1412) );
  AOI22D1BWP30P140LVT U1792 ( .A1(i_data_bus[869]), .A2(n1941), .B1(
        i_data_bus[741]), .B2(n1945), .ZN(n1411) );
  AOI22D1BWP30P140LVT U1793 ( .A1(i_data_bus[677]), .A2(n1947), .B1(
        i_data_bus[805]), .B2(n1943), .ZN(n1410) );
  AOI22D1BWP30P140LVT U1794 ( .A1(i_data_bus[645]), .A2(n1944), .B1(
        i_data_bus[709]), .B2(n1942), .ZN(n1409) );
  ND4D1BWP30P140LVT U1795 ( .A1(n1412), .A2(n1411), .A3(n1410), .A4(n1409), 
        .ZN(n1413) );
  OR4D1BWP30P140LVT U1796 ( .A1(n1416), .A2(n1415), .A3(n1414), .A4(n1413), 
        .Z(o_data_bus[101]) );
  AOI22D1BWP30P140LVT U1797 ( .A1(i_data_bus[966]), .A2(n1923), .B1(
        i_data_bus[518]), .B2(n1927), .ZN(n1420) );
  AOI22D1BWP30P140LVT U1798 ( .A1(i_data_bus[6]), .A2(n2), .B1(i_data_bus[102]), .B2(n1936), .ZN(n1419) );
  AOI22D1BWP30P140LVT U1799 ( .A1(i_data_bus[902]), .A2(n128), .B1(
        i_data_bus[326]), .B2(n1913), .ZN(n1418) );
  AOI22D1BWP30P140LVT U1800 ( .A1(i_data_bus[582]), .A2(n1912), .B1(
        i_data_bus[38]), .B2(n1914), .ZN(n1417) );
  AOI22D1BWP30P140LVT U1801 ( .A1(i_data_bus[358]), .A2(n1926), .B1(
        i_data_bus[294]), .B2(n1922), .ZN(n1424) );
  AOI22D1BWP30P140LVT U1802 ( .A1(i_data_bus[166]), .A2(n1915), .B1(
        i_data_bus[422]), .B2(n1921), .ZN(n1423) );
  AOI22D1BWP30P140LVT U1803 ( .A1(i_data_bus[486]), .A2(n1932), .B1(
        i_data_bus[390]), .B2(n1279), .ZN(n1422) );
  AOI22D1BWP30P140LVT U1804 ( .A1(i_data_bus[550]), .A2(n1924), .B1(
        i_data_bus[230]), .B2(n1911), .ZN(n1421) );
  AOI22D1BWP30P140LVT U1805 ( .A1(i_data_bus[998]), .A2(n1934), .B1(
        i_data_bus[262]), .B2(n1293), .ZN(n1428) );
  AOI22D1BWP30P140LVT U1806 ( .A1(i_data_bus[614]), .A2(n1910), .B1(
        i_data_bus[934]), .B2(n127), .ZN(n1427) );
  AOI22D1BWP30P140LVT U1807 ( .A1(i_data_bus[198]), .A2(n1916), .B1(
        i_data_bus[134]), .B2(n1935), .ZN(n1426) );
  AOI22D1BWP30P140LVT U1808 ( .A1(i_data_bus[70]), .A2(n1925), .B1(
        i_data_bus[454]), .B2(n1933), .ZN(n1425) );
  AOI22D1BWP30P140LVT U1809 ( .A1(i_data_bus[838]), .A2(n1948), .B1(
        i_data_bus[646]), .B2(n1944), .ZN(n1432) );
  AOI22D1BWP30P140LVT U1810 ( .A1(i_data_bus[870]), .A2(n1941), .B1(
        i_data_bus[678]), .B2(n1947), .ZN(n1431) );
  AOI22D1BWP30P140LVT U1811 ( .A1(i_data_bus[742]), .A2(n1945), .B1(
        i_data_bus[774]), .B2(n1946), .ZN(n1430) );
  AOI22D1BWP30P140LVT U1812 ( .A1(i_data_bus[806]), .A2(n1943), .B1(
        i_data_bus[710]), .B2(n1942), .ZN(n1429) );
  ND4D1BWP30P140LVT U1813 ( .A1(n1432), .A2(n1431), .A3(n1430), .A4(n1429), 
        .ZN(n1433) );
  AOI22D1BWP30P140LVT U1814 ( .A1(i_data_bus[551]), .A2(n1924), .B1(
        i_data_bus[135]), .B2(n1935), .ZN(n1437) );
  AOI22D1BWP30P140LVT U1815 ( .A1(i_data_bus[39]), .A2(n1914), .B1(
        i_data_bus[999]), .B2(n1934), .ZN(n1436) );
  AOI22D1BWP30P140LVT U1816 ( .A1(i_data_bus[295]), .A2(n1922), .B1(
        i_data_bus[199]), .B2(n1916), .ZN(n1435) );
  AOI22D1BWP30P140LVT U1817 ( .A1(i_data_bus[903]), .A2(n128), .B1(
        i_data_bus[167]), .B2(n1915), .ZN(n1434) );
  ND4D1BWP30P140LVT U1818 ( .A1(n1437), .A2(n1436), .A3(n1435), .A4(n1434), 
        .ZN(n1453) );
  AOI22D1BWP30P140LVT U1819 ( .A1(i_data_bus[519]), .A2(n1927), .B1(
        i_data_bus[487]), .B2(n1932), .ZN(n1441) );
  AOI22D1BWP30P140LVT U1820 ( .A1(i_data_bus[103]), .A2(n1936), .B1(
        i_data_bus[935]), .B2(n127), .ZN(n1440) );
  AOI22D1BWP30P140LVT U1821 ( .A1(i_data_bus[583]), .A2(n1912), .B1(
        i_data_bus[263]), .B2(n1293), .ZN(n1439) );
  AOI22D1BWP30P140LVT U1822 ( .A1(i_data_bus[455]), .A2(n1933), .B1(
        i_data_bus[231]), .B2(n1911), .ZN(n1438) );
  ND4D1BWP30P140LVT U1823 ( .A1(n1441), .A2(n1440), .A3(n1439), .A4(n1438), 
        .ZN(n1452) );
  AOI22D1BWP30P140LVT U1824 ( .A1(i_data_bus[391]), .A2(n1279), .B1(
        i_data_bus[423]), .B2(n1921), .ZN(n1445) );
  AOI22D1BWP30P140LVT U1825 ( .A1(i_data_bus[615]), .A2(n1910), .B1(
        i_data_bus[7]), .B2(n2), .ZN(n1444) );
  AOI22D1BWP30P140LVT U1826 ( .A1(i_data_bus[359]), .A2(n1926), .B1(
        i_data_bus[327]), .B2(n1913), .ZN(n1442) );
  ND4D1BWP30P140LVT U1827 ( .A1(n1445), .A2(n1444), .A3(n1443), .A4(n1442), 
        .ZN(n1451) );
  AOI22D1BWP30P140LVT U1828 ( .A1(i_data_bus[743]), .A2(n1945), .B1(
        i_data_bus[775]), .B2(n1946), .ZN(n1449) );
  AOI22D1BWP30P140LVT U1829 ( .A1(i_data_bus[807]), .A2(n1943), .B1(
        i_data_bus[647]), .B2(n1944), .ZN(n1448) );
  AOI22D1BWP30P140LVT U1830 ( .A1(i_data_bus[679]), .A2(n1947), .B1(
        i_data_bus[711]), .B2(n1942), .ZN(n1447) );
  AOI22D1BWP30P140LVT U1831 ( .A1(i_data_bus[871]), .A2(n1941), .B1(
        i_data_bus[839]), .B2(n1948), .ZN(n1446) );
  ND4D1BWP30P140LVT U1832 ( .A1(n1449), .A2(n1448), .A3(n1447), .A4(n1446), 
        .ZN(n1450) );
  OR4D1BWP30P140LVT U1833 ( .A1(n1453), .A2(n1452), .A3(n1451), .A4(n1450), 
        .Z(o_data_bus[103]) );
  AOI22D1BWP30P140LVT U1834 ( .A1(i_data_bus[584]), .A2(n1912), .B1(
        i_data_bus[200]), .B2(n1916), .ZN(n1457) );
  AOI22D1BWP30P140LVT U1835 ( .A1(i_data_bus[104]), .A2(n1936), .B1(
        i_data_bus[168]), .B2(n1915), .ZN(n1456) );
  AOI22D1BWP30P140LVT U1836 ( .A1(i_data_bus[520]), .A2(n1927), .B1(
        i_data_bus[456]), .B2(n1933), .ZN(n1455) );
  AOI22D1BWP30P140LVT U1837 ( .A1(i_data_bus[968]), .A2(n1923), .B1(
        i_data_bus[424]), .B2(n1921), .ZN(n1454) );
  ND4D1BWP30P140LVT U1838 ( .A1(n1457), .A2(n1456), .A3(n1455), .A4(n1454), 
        .ZN(n1473) );
  AOI22D1BWP30P140LVT U1839 ( .A1(i_data_bus[360]), .A2(n1926), .B1(
        i_data_bus[232]), .B2(n1911), .ZN(n1461) );
  AOI22D1BWP30P140LVT U1840 ( .A1(i_data_bus[1000]), .A2(n1934), .B1(
        i_data_bus[136]), .B2(n1935), .ZN(n1460) );
  AOI22D1BWP30P140LVT U1841 ( .A1(i_data_bus[8]), .A2(n2), .B1(i_data_bus[488]), .B2(n1932), .ZN(n1459) );
  AOI22D1BWP30P140LVT U1842 ( .A1(i_data_bus[936]), .A2(n127), .B1(
        i_data_bus[392]), .B2(n1279), .ZN(n1458) );
  ND4D1BWP30P140LVT U1843 ( .A1(n1461), .A2(n1460), .A3(n1459), .A4(n1458), 
        .ZN(n1472) );
  AOI22D1BWP30P140LVT U1844 ( .A1(i_data_bus[616]), .A2(n1910), .B1(
        i_data_bus[328]), .B2(n1913), .ZN(n1465) );
  AOI22D1BWP30P140LVT U1845 ( .A1(i_data_bus[264]), .A2(n1293), .B1(
        i_data_bus[296]), .B2(n1922), .ZN(n1464) );
  ND4D1BWP30P140LVT U1846 ( .A1(n1465), .A2(n1464), .A3(n1463), .A4(n1462), 
        .ZN(n1471) );
  AOI22D1BWP30P140LVT U1847 ( .A1(i_data_bus[680]), .A2(n1947), .B1(
        i_data_bus[808]), .B2(n1943), .ZN(n1469) );
  AOI22D1BWP30P140LVT U1848 ( .A1(i_data_bus[712]), .A2(n1942), .B1(
        i_data_bus[776]), .B2(n1946), .ZN(n1468) );
  AOI22D1BWP30P140LVT U1849 ( .A1(i_data_bus[744]), .A2(n1945), .B1(
        i_data_bus[648]), .B2(n1944), .ZN(n1467) );
  AOI22D1BWP30P140LVT U1850 ( .A1(i_data_bus[840]), .A2(n1948), .B1(
        i_data_bus[872]), .B2(n1941), .ZN(n1466) );
  ND4D1BWP30P140LVT U1851 ( .A1(n1469), .A2(n1468), .A3(n1467), .A4(n1466), 
        .ZN(n1470) );
  OR4D1BWP30P140LVT U1852 ( .A1(n1473), .A2(n1472), .A3(n1471), .A4(n1470), 
        .Z(o_data_bus[104]) );
  AOI22D1BWP30P140LVT U1853 ( .A1(i_data_bus[1001]), .A2(n1934), .B1(
        i_data_bus[169]), .B2(n1915), .ZN(n1476) );
  AOI22D1BWP30P140LVT U1854 ( .A1(i_data_bus[489]), .A2(n1932), .B1(
        i_data_bus[137]), .B2(n1935), .ZN(n1474) );
  ND4D1BWP30P140LVT U1855 ( .A1(n1477), .A2(n1476), .A3(n1475), .A4(n1474), 
        .ZN(n1493) );
  AOI22D1BWP30P140LVT U1856 ( .A1(i_data_bus[617]), .A2(n1910), .B1(
        i_data_bus[297]), .B2(n1922), .ZN(n1481) );
  AOI22D1BWP30P140LVT U1857 ( .A1(i_data_bus[105]), .A2(n1936), .B1(
        i_data_bus[457]), .B2(n1933), .ZN(n1480) );
  AOI22D1BWP30P140LVT U1858 ( .A1(i_data_bus[969]), .A2(n1923), .B1(
        i_data_bus[329]), .B2(n1913), .ZN(n1479) );
  AOI22D1BWP30P140LVT U1859 ( .A1(i_data_bus[585]), .A2(n1912), .B1(
        i_data_bus[361]), .B2(n1926), .ZN(n1478) );
  ND4D1BWP30P140LVT U1860 ( .A1(n1481), .A2(n1480), .A3(n1479), .A4(n1478), 
        .ZN(n1492) );
  AOI22D1BWP30P140LVT U1861 ( .A1(i_data_bus[937]), .A2(n127), .B1(
        i_data_bus[425]), .B2(n1921), .ZN(n1485) );
  AOI22D1BWP30P140LVT U1862 ( .A1(i_data_bus[201]), .A2(n1916), .B1(
        i_data_bus[265]), .B2(n1293), .ZN(n1484) );
  AOI22D1BWP30P140LVT U1863 ( .A1(i_data_bus[9]), .A2(n2), .B1(i_data_bus[553]), .B2(n1924), .ZN(n1483) );
  AOI22D1BWP30P140LVT U1864 ( .A1(i_data_bus[233]), .A2(n1911), .B1(
        i_data_bus[393]), .B2(n1279), .ZN(n1482) );
  ND4D1BWP30P140LVT U1865 ( .A1(n1485), .A2(n1484), .A3(n1483), .A4(n1482), 
        .ZN(n1491) );
  AOI22D1BWP30P140LVT U1866 ( .A1(i_data_bus[873]), .A2(n1941), .B1(
        i_data_bus[841]), .B2(n1948), .ZN(n1489) );
  AOI22D1BWP30P140LVT U1867 ( .A1(i_data_bus[809]), .A2(n1943), .B1(
        i_data_bus[777]), .B2(n1946), .ZN(n1488) );
  AOI22D1BWP30P140LVT U1868 ( .A1(i_data_bus[681]), .A2(n1947), .B1(
        i_data_bus[713]), .B2(n1942), .ZN(n1487) );
  AOI22D1BWP30P140LVT U1869 ( .A1(i_data_bus[745]), .A2(n1945), .B1(
        i_data_bus[649]), .B2(n1944), .ZN(n1486) );
  ND4D1BWP30P140LVT U1870 ( .A1(n1489), .A2(n1488), .A3(n1487), .A4(n1486), 
        .ZN(n1490) );
  OR4D1BWP30P140LVT U1871 ( .A1(n1493), .A2(n1492), .A3(n1491), .A4(n1490), 
        .Z(o_data_bus[105]) );
  AOI22D1BWP30P140LVT U1872 ( .A1(i_data_bus[906]), .A2(n128), .B1(
        i_data_bus[394]), .B2(n1279), .ZN(n1497) );
  AOI22D1BWP30P140LVT U1873 ( .A1(i_data_bus[106]), .A2(n1936), .B1(
        i_data_bus[938]), .B2(n127), .ZN(n1496) );
  AOI22D1BWP30P140LVT U1874 ( .A1(i_data_bus[202]), .A2(n1916), .B1(
        i_data_bus[298]), .B2(n1922), .ZN(n1495) );
  AOI22D1BWP30P140LVT U1875 ( .A1(i_data_bus[490]), .A2(n1932), .B1(
        i_data_bus[266]), .B2(n1293), .ZN(n1494) );
  ND4D1BWP30P140LVT U1876 ( .A1(n1497), .A2(n1496), .A3(n1495), .A4(n1494), 
        .ZN(n1513) );
  AOI22D1BWP30P140LVT U1877 ( .A1(i_data_bus[554]), .A2(n1924), .B1(
        i_data_bus[458]), .B2(n1933), .ZN(n1501) );
  AOI22D1BWP30P140LVT U1878 ( .A1(i_data_bus[234]), .A2(n1911), .B1(
        i_data_bus[426]), .B2(n1921), .ZN(n1500) );
  AOI22D1BWP30P140LVT U1879 ( .A1(i_data_bus[1002]), .A2(n1934), .B1(
        i_data_bus[138]), .B2(n1935), .ZN(n1499) );
  AOI22D1BWP30P140LVT U1880 ( .A1(i_data_bus[970]), .A2(n1923), .B1(
        i_data_bus[362]), .B2(n1926), .ZN(n1498) );
  ND4D1BWP30P140LVT U1881 ( .A1(n1501), .A2(n1500), .A3(n1499), .A4(n1498), 
        .ZN(n1512) );
  AOI22D1BWP30P140LVT U1882 ( .A1(i_data_bus[74]), .A2(n1925), .B1(
        i_data_bus[522]), .B2(n1927), .ZN(n1505) );
  AOI22D1BWP30P140LVT U1883 ( .A1(i_data_bus[586]), .A2(n1912), .B1(
        i_data_bus[330]), .B2(n1913), .ZN(n1504) );
  AOI22D1BWP30P140LVT U1884 ( .A1(i_data_bus[10]), .A2(n2), .B1(
        i_data_bus[618]), .B2(n1910), .ZN(n1503) );
  AOI22D1BWP30P140LVT U1885 ( .A1(i_data_bus[42]), .A2(n1914), .B1(
        i_data_bus[170]), .B2(n1915), .ZN(n1502) );
  ND4D1BWP30P140LVT U1886 ( .A1(n1505), .A2(n1504), .A3(n1503), .A4(n1502), 
        .ZN(n1511) );
  AOI22D1BWP30P140LVT U1887 ( .A1(i_data_bus[874]), .A2(n1941), .B1(
        i_data_bus[714]), .B2(n1942), .ZN(n1509) );
  AOI22D1BWP30P140LVT U1888 ( .A1(i_data_bus[842]), .A2(n1948), .B1(
        i_data_bus[682]), .B2(n1947), .ZN(n1508) );
  AOI22D1BWP30P140LVT U1889 ( .A1(i_data_bus[778]), .A2(n1946), .B1(
        i_data_bus[810]), .B2(n1943), .ZN(n1507) );
  AOI22D1BWP30P140LVT U1890 ( .A1(i_data_bus[650]), .A2(n1944), .B1(
        i_data_bus[746]), .B2(n1945), .ZN(n1506) );
  ND4D1BWP30P140LVT U1891 ( .A1(n1509), .A2(n1508), .A3(n1507), .A4(n1506), 
        .ZN(n1510) );
  OR4D1BWP30P140LVT U1892 ( .A1(n1513), .A2(n1512), .A3(n1511), .A4(n1510), 
        .Z(o_data_bus[106]) );
  AOI22D1BWP30P140LVT U1893 ( .A1(i_data_bus[523]), .A2(n1927), .B1(
        i_data_bus[203]), .B2(n1916), .ZN(n1517) );
  AOI22D1BWP30P140LVT U1894 ( .A1(i_data_bus[555]), .A2(n1924), .B1(
        i_data_bus[139]), .B2(n1935), .ZN(n1516) );
  AOI22D1BWP30P140LVT U1895 ( .A1(i_data_bus[43]), .A2(n1914), .B1(
        i_data_bus[171]), .B2(n1915), .ZN(n1515) );
  AOI22D1BWP30P140LVT U1896 ( .A1(i_data_bus[427]), .A2(n1921), .B1(
        i_data_bus[299]), .B2(n1922), .ZN(n1514) );
  ND4D1BWP30P140LVT U1897 ( .A1(n1517), .A2(n1516), .A3(n1515), .A4(n1514), 
        .ZN(n1533) );
  AOI22D1BWP30P140LVT U1898 ( .A1(i_data_bus[235]), .A2(n1911), .B1(
        i_data_bus[267]), .B2(n1293), .ZN(n1521) );
  AOI22D1BWP30P140LVT U1899 ( .A1(i_data_bus[907]), .A2(n128), .B1(
        i_data_bus[363]), .B2(n1926), .ZN(n1520) );
  AOI22D1BWP30P140LVT U1900 ( .A1(i_data_bus[1003]), .A2(n1934), .B1(
        i_data_bus[491]), .B2(n1932), .ZN(n1519) );
  AOI22D1BWP30P140LVT U1901 ( .A1(i_data_bus[587]), .A2(n1912), .B1(
        i_data_bus[395]), .B2(n1279), .ZN(n1518) );
  ND4D1BWP30P140LVT U1902 ( .A1(n1521), .A2(n1520), .A3(n1519), .A4(n1518), 
        .ZN(n1532) );
  AOI22D1BWP30P140LVT U1903 ( .A1(i_data_bus[11]), .A2(n2), .B1(
        i_data_bus[459]), .B2(n1933), .ZN(n1525) );
  AOI22D1BWP30P140LVT U1904 ( .A1(i_data_bus[619]), .A2(n1910), .B1(
        i_data_bus[331]), .B2(n1913), .ZN(n1524) );
  AOI22D1BWP30P140LVT U1905 ( .A1(i_data_bus[939]), .A2(n127), .B1(
        i_data_bus[107]), .B2(n1936), .ZN(n1523) );
  ND4D1BWP30P140LVT U1906 ( .A1(n1523), .A2(n1524), .A3(n1525), .A4(n1522), 
        .ZN(n1531) );
  AOI22D1BWP30P140LVT U1907 ( .A1(i_data_bus[843]), .A2(n1948), .B1(
        i_data_bus[779]), .B2(n1946), .ZN(n1529) );
  AOI22D1BWP30P140LVT U1908 ( .A1(i_data_bus[875]), .A2(n1941), .B1(
        i_data_bus[715]), .B2(n1942), .ZN(n1528) );
  AOI22D1BWP30P140LVT U1909 ( .A1(i_data_bus[811]), .A2(n1943), .B1(
        i_data_bus[683]), .B2(n1947), .ZN(n1527) );
  AOI22D1BWP30P140LVT U1910 ( .A1(i_data_bus[747]), .A2(n1945), .B1(
        i_data_bus[651]), .B2(n1944), .ZN(n1526) );
  ND4D1BWP30P140LVT U1911 ( .A1(n1529), .A2(n1528), .A3(n1527), .A4(n1526), 
        .ZN(n1530) );
  OR4D1BWP30P140LVT U1912 ( .A1(n1533), .A2(n1532), .A3(n1530), .A4(n1531), 
        .Z(o_data_bus[107]) );
  AOI22D1BWP30P140LVT U1913 ( .A1(i_data_bus[556]), .A2(n1924), .B1(
        i_data_bus[588]), .B2(n1912), .ZN(n1537) );
  AOI22D1BWP30P140LVT U1914 ( .A1(i_data_bus[1004]), .A2(n1934), .B1(
        i_data_bus[364]), .B2(n1926), .ZN(n1536) );
  AOI22D1BWP30P140LVT U1915 ( .A1(i_data_bus[428]), .A2(n1921), .B1(
        i_data_bus[204]), .B2(n1916), .ZN(n1535) );
  AOI22D1BWP30P140LVT U1916 ( .A1(i_data_bus[12]), .A2(n2), .B1(
        i_data_bus[908]), .B2(n128), .ZN(n1534) );
  ND4D1BWP30P140LVT U1917 ( .A1(n1537), .A2(n1536), .A3(n1535), .A4(n1534), 
        .ZN(n1553) );
  AOI22D1BWP30P140LVT U1918 ( .A1(i_data_bus[140]), .A2(n1935), .B1(
        i_data_bus[396]), .B2(n1279), .ZN(n1540) );
  AOI22D1BWP30P140LVT U1919 ( .A1(i_data_bus[236]), .A2(n1911), .B1(
        i_data_bus[172]), .B2(n1915), .ZN(n1539) );
  AOI22D1BWP30P140LVT U1920 ( .A1(i_data_bus[460]), .A2(n1933), .B1(
        i_data_bus[268]), .B2(n1293), .ZN(n1538) );
  ND4D1BWP30P140LVT U1921 ( .A1(n1541), .A2(n1540), .A3(n1539), .A4(n1538), 
        .ZN(n1552) );
  AOI22D1BWP30P140LVT U1922 ( .A1(i_data_bus[300]), .A2(n1922), .B1(
        i_data_bus[332]), .B2(n1913), .ZN(n1545) );
  AOI22D1BWP30P140LVT U1923 ( .A1(i_data_bus[76]), .A2(n1925), .B1(
        i_data_bus[492]), .B2(n1932), .ZN(n1544) );
  AOI22D1BWP30P140LVT U1924 ( .A1(i_data_bus[940]), .A2(n127), .B1(
        i_data_bus[524]), .B2(n1927), .ZN(n1542) );
  ND4D1BWP30P140LVT U1925 ( .A1(n1545), .A2(n1544), .A3(n1543), .A4(n1542), 
        .ZN(n1551) );
  AOI22D1BWP30P140LVT U1926 ( .A1(i_data_bus[780]), .A2(n1946), .B1(
        i_data_bus[652]), .B2(n1944), .ZN(n1549) );
  AOI22D1BWP30P140LVT U1927 ( .A1(i_data_bus[812]), .A2(n1943), .B1(
        i_data_bus[876]), .B2(n1941), .ZN(n1548) );
  AOI22D1BWP30P140LVT U1928 ( .A1(i_data_bus[684]), .A2(n1947), .B1(
        i_data_bus[844]), .B2(n1948), .ZN(n1547) );
  AOI22D1BWP30P140LVT U1929 ( .A1(i_data_bus[716]), .A2(n1942), .B1(
        i_data_bus[748]), .B2(n1945), .ZN(n1546) );
  ND4D1BWP30P140LVT U1930 ( .A1(n1549), .A2(n1548), .A3(n1547), .A4(n1546), 
        .ZN(n1550) );
  OR4D1BWP30P140LVT U1931 ( .A1(n1553), .A2(n1552), .A3(n1551), .A4(n1550), 
        .Z(o_data_bus[108]) );
  AOI22D1BWP30P140LVT U1932 ( .A1(i_data_bus[973]), .A2(n1923), .B1(
        i_data_bus[493]), .B2(n1932), .ZN(n1557) );
  AOI22D1BWP30P140LVT U1933 ( .A1(i_data_bus[397]), .A2(n1279), .B1(
        i_data_bus[365]), .B2(n1926), .ZN(n1556) );
  AOI22D1BWP30P140LVT U1934 ( .A1(i_data_bus[621]), .A2(n1910), .B1(
        i_data_bus[141]), .B2(n1935), .ZN(n1555) );
  AOI22D1BWP30P140LVT U1935 ( .A1(i_data_bus[589]), .A2(n1912), .B1(
        i_data_bus[13]), .B2(n2), .ZN(n1554) );
  ND4D1BWP30P140LVT U1936 ( .A1(n1557), .A2(n1556), .A3(n1555), .A4(n1554), 
        .ZN(n1573) );
  AOI22D1BWP30P140LVT U1937 ( .A1(i_data_bus[45]), .A2(n1914), .B1(
        i_data_bus[525]), .B2(n1927), .ZN(n1561) );
  AOI22D1BWP30P140LVT U1938 ( .A1(i_data_bus[941]), .A2(n127), .B1(
        i_data_bus[461]), .B2(n1933), .ZN(n1560) );
  AOI22D1BWP30P140LVT U1939 ( .A1(i_data_bus[77]), .A2(n1925), .B1(
        i_data_bus[205]), .B2(n1916), .ZN(n1558) );
  ND4D1BWP30P140LVT U1940 ( .A1(n1561), .A2(n1560), .A3(n1559), .A4(n1558), 
        .ZN(n1572) );
  AOI22D1BWP30P140LVT U1941 ( .A1(i_data_bus[429]), .A2(n1921), .B1(
        i_data_bus[301]), .B2(n1922), .ZN(n1565) );
  AOI22D1BWP30P140LVT U1942 ( .A1(i_data_bus[237]), .A2(n1911), .B1(
        i_data_bus[269]), .B2(n1293), .ZN(n1564) );
  AOI22D1BWP30P140LVT U1943 ( .A1(i_data_bus[1005]), .A2(n1934), .B1(
        i_data_bus[173]), .B2(n1915), .ZN(n1563) );
  AOI22D1BWP30P140LVT U1944 ( .A1(i_data_bus[557]), .A2(n1924), .B1(
        i_data_bus[333]), .B2(n1913), .ZN(n1562) );
  ND4D1BWP30P140LVT U1945 ( .A1(n1565), .A2(n1564), .A3(n1563), .A4(n1562), 
        .ZN(n1571) );
  AOI22D1BWP30P140LVT U1946 ( .A1(i_data_bus[877]), .A2(n1941), .B1(
        i_data_bus[717]), .B2(n1942), .ZN(n1569) );
  AOI22D1BWP30P140LVT U1947 ( .A1(i_data_bus[781]), .A2(n1946), .B1(
        i_data_bus[813]), .B2(n1943), .ZN(n1568) );
  AOI22D1BWP30P140LVT U1948 ( .A1(i_data_bus[749]), .A2(n1945), .B1(
        i_data_bus[685]), .B2(n1947), .ZN(n1567) );
  AOI22D1BWP30P140LVT U1949 ( .A1(i_data_bus[845]), .A2(n1948), .B1(
        i_data_bus[653]), .B2(n1944), .ZN(n1566) );
  ND4D1BWP30P140LVT U1950 ( .A1(n1569), .A2(n1568), .A3(n1567), .A4(n1566), 
        .ZN(n1570) );
  OR4D1BWP30P140LVT U1951 ( .A1(n1573), .A2(n1572), .A3(n1571), .A4(n1570), 
        .Z(o_data_bus[109]) );
  AOI22D1BWP30P140LVT U1952 ( .A1(i_data_bus[14]), .A2(n2), .B1(
        i_data_bus[398]), .B2(n1279), .ZN(n1577) );
  AOI22D1BWP30P140LVT U1953 ( .A1(i_data_bus[910]), .A2(n128), .B1(
        i_data_bus[974]), .B2(n1923), .ZN(n1576) );
  AOI22D1BWP30P140LVT U1954 ( .A1(i_data_bus[558]), .A2(n1924), .B1(
        i_data_bus[302]), .B2(n1922), .ZN(n1575) );
  AOI22D1BWP30P140LVT U1955 ( .A1(i_data_bus[174]), .A2(n1915), .B1(
        i_data_bus[334]), .B2(n1913), .ZN(n1574) );
  ND4D1BWP30P140LVT U1956 ( .A1(n1577), .A2(n1576), .A3(n1575), .A4(n1574), 
        .ZN(n1593) );
  AOI22D1BWP30P140LVT U1957 ( .A1(i_data_bus[622]), .A2(n1910), .B1(
        i_data_bus[270]), .B2(n1293), .ZN(n1581) );
  AOI22D1BWP30P140LVT U1958 ( .A1(i_data_bus[78]), .A2(n1925), .B1(
        i_data_bus[46]), .B2(n1914), .ZN(n1580) );
  AOI22D1BWP30P140LVT U1959 ( .A1(i_data_bus[590]), .A2(n1912), .B1(
        i_data_bus[238]), .B2(n1911), .ZN(n1579) );
  AOI22D1BWP30P140LVT U1960 ( .A1(i_data_bus[110]), .A2(n1936), .B1(
        i_data_bus[142]), .B2(n1935), .ZN(n1578) );
  ND4D1BWP30P140LVT U1961 ( .A1(n1580), .A2(n1581), .A3(n1579), .A4(n1578), 
        .ZN(n1592) );
  AOI22D1BWP30P140LVT U1962 ( .A1(i_data_bus[942]), .A2(n127), .B1(
        i_data_bus[462]), .B2(n1933), .ZN(n1585) );
  AOI22D1BWP30P140LVT U1963 ( .A1(i_data_bus[1006]), .A2(n1934), .B1(
        i_data_bus[430]), .B2(n1921), .ZN(n1584) );
  AOI22D1BWP30P140LVT U1964 ( .A1(i_data_bus[206]), .A2(n1916), .B1(
        i_data_bus[494]), .B2(n1932), .ZN(n1583) );
  AOI22D1BWP30P140LVT U1965 ( .A1(i_data_bus[526]), .A2(n1927), .B1(
        i_data_bus[366]), .B2(n1926), .ZN(n1582) );
  ND4D1BWP30P140LVT U1966 ( .A1(n1585), .A2(n1584), .A3(n1583), .A4(n1582), 
        .ZN(n1591) );
  AOI22D1BWP30P140LVT U1967 ( .A1(i_data_bus[846]), .A2(n1948), .B1(
        i_data_bus[750]), .B2(n1945), .ZN(n1589) );
  AOI22D1BWP30P140LVT U1968 ( .A1(i_data_bus[782]), .A2(n1946), .B1(
        i_data_bus[878]), .B2(n1941), .ZN(n1588) );
  AOI22D1BWP30P140LVT U1969 ( .A1(i_data_bus[686]), .A2(n1947), .B1(
        i_data_bus[654]), .B2(n1944), .ZN(n1587) );
  AOI22D1BWP30P140LVT U1970 ( .A1(i_data_bus[814]), .A2(n1943), .B1(
        i_data_bus[718]), .B2(n1942), .ZN(n1586) );
  ND4D1BWP30P140LVT U1971 ( .A1(n1589), .A2(n1588), .A3(n1587), .A4(n1586), 
        .ZN(n1590) );
  OR4D1BWP30P140LVT U1972 ( .A1(n1593), .A2(n1590), .A3(n1591), .A4(n1592), 
        .Z(o_data_bus[110]) );
  AOI22D1BWP30P140LVT U1973 ( .A1(i_data_bus[911]), .A2(n128), .B1(
        i_data_bus[1007]), .B2(n1934), .ZN(n1597) );
  AOI22D1BWP30P140LVT U1974 ( .A1(i_data_bus[111]), .A2(n1936), .B1(
        i_data_bus[175]), .B2(n1915), .ZN(n1596) );
  AOI22D1BWP30P140LVT U1975 ( .A1(i_data_bus[591]), .A2(n1912), .B1(
        i_data_bus[239]), .B2(n1911), .ZN(n1595) );
  AOI22D1BWP30P140LVT U1976 ( .A1(i_data_bus[975]), .A2(n1923), .B1(
        i_data_bus[79]), .B2(n1925), .ZN(n1594) );
  AOI22D1BWP30P140LVT U1977 ( .A1(i_data_bus[47]), .A2(n1914), .B1(
        i_data_bus[303]), .B2(n1922), .ZN(n1601) );
  AOI22D1BWP30P140LVT U1978 ( .A1(i_data_bus[527]), .A2(n1927), .B1(
        i_data_bus[335]), .B2(n1913), .ZN(n1600) );
  AOI22D1BWP30P140LVT U1979 ( .A1(i_data_bus[207]), .A2(n1916), .B1(
        i_data_bus[367]), .B2(n1926), .ZN(n1599) );
  AOI22D1BWP30P140LVT U1980 ( .A1(i_data_bus[271]), .A2(n1293), .B1(
        i_data_bus[143]), .B2(n1935), .ZN(n1598) );
  AOI22D1BWP30P140LVT U1981 ( .A1(i_data_bus[559]), .A2(n1924), .B1(
        i_data_bus[15]), .B2(n2), .ZN(n1605) );
  AOI22D1BWP30P140LVT U1982 ( .A1(i_data_bus[431]), .A2(n1921), .B1(
        i_data_bus[463]), .B2(n1933), .ZN(n1604) );
  AOI22D1BWP30P140LVT U1983 ( .A1(i_data_bus[943]), .A2(n127), .B1(
        i_data_bus[399]), .B2(n1279), .ZN(n1603) );
  AOI22D1BWP30P140LVT U1984 ( .A1(i_data_bus[623]), .A2(n1910), .B1(
        i_data_bus[495]), .B2(n1932), .ZN(n1602) );
  AOI22D1BWP30P140LVT U1985 ( .A1(i_data_bus[655]), .A2(n1944), .B1(
        i_data_bus[879]), .B2(n1941), .ZN(n1609) );
  AOI22D1BWP30P140LVT U1986 ( .A1(i_data_bus[719]), .A2(n1942), .B1(
        i_data_bus[687]), .B2(n1947), .ZN(n1608) );
  AOI22D1BWP30P140LVT U1987 ( .A1(i_data_bus[847]), .A2(n1948), .B1(
        i_data_bus[783]), .B2(n1946), .ZN(n1607) );
  AOI22D1BWP30P140LVT U1988 ( .A1(i_data_bus[751]), .A2(n1945), .B1(
        i_data_bus[815]), .B2(n1943), .ZN(n1606) );
  AOI22D1BWP30P140LVT U1989 ( .A1(i_data_bus[80]), .A2(n1925), .B1(
        i_data_bus[368]), .B2(n1926), .ZN(n1614) );
  AOI22D1BWP30P140LVT U1990 ( .A1(i_data_bus[1008]), .A2(n1934), .B1(
        i_data_bus[240]), .B2(n1911), .ZN(n1613) );
  AOI22D1BWP30P140LVT U1991 ( .A1(i_data_bus[560]), .A2(n1924), .B1(
        i_data_bus[528]), .B2(n1927), .ZN(n1611) );
  ND4D1BWP30P140LVT U1992 ( .A1(n1614), .A2(n1613), .A3(n1612), .A4(n1611), 
        .ZN(n1630) );
  AOI22D1BWP30P140LVT U1993 ( .A1(i_data_bus[48]), .A2(n1914), .B1(
        i_data_bus[208]), .B2(n1916), .ZN(n1618) );
  AOI22D1BWP30P140LVT U1994 ( .A1(i_data_bus[336]), .A2(n1913), .B1(
        i_data_bus[144]), .B2(n1935), .ZN(n1617) );
  AOI22D1BWP30P140LVT U1995 ( .A1(i_data_bus[592]), .A2(n1912), .B1(
        i_data_bus[304]), .B2(n1922), .ZN(n1616) );
  AOI22D1BWP30P140LVT U1996 ( .A1(i_data_bus[496]), .A2(n1932), .B1(
        i_data_bus[272]), .B2(n1293), .ZN(n1615) );
  ND4D1BWP30P140LVT U1997 ( .A1(n1618), .A2(n1617), .A3(n1616), .A4(n1615), 
        .ZN(n1629) );
  AOI22D1BWP30P140LVT U1998 ( .A1(i_data_bus[16]), .A2(n2), .B1(
        i_data_bus[464]), .B2(n1933), .ZN(n1622) );
  AOI22D1BWP30P140LVT U1999 ( .A1(i_data_bus[624]), .A2(n1910), .B1(
        i_data_bus[400]), .B2(n1279), .ZN(n1621) );
  AOI22D1BWP30P140LVT U2000 ( .A1(i_data_bus[944]), .A2(n127), .B1(
        i_data_bus[432]), .B2(n1921), .ZN(n1620) );
  AOI22D1BWP30P140LVT U2001 ( .A1(i_data_bus[976]), .A2(n1923), .B1(
        i_data_bus[176]), .B2(n1915), .ZN(n1619) );
  ND4D1BWP30P140LVT U2002 ( .A1(n1622), .A2(n1621), .A3(n1620), .A4(n1619), 
        .ZN(n1628) );
  AOI22D1BWP30P140LVT U2003 ( .A1(i_data_bus[656]), .A2(n1944), .B1(
        i_data_bus[848]), .B2(n1948), .ZN(n1626) );
  AOI22D1BWP30P140LVT U2004 ( .A1(i_data_bus[880]), .A2(n1941), .B1(
        i_data_bus[688]), .B2(n1947), .ZN(n1625) );
  AOI22D1BWP30P140LVT U2005 ( .A1(i_data_bus[752]), .A2(n1945), .B1(
        i_data_bus[720]), .B2(n1942), .ZN(n1624) );
  AOI22D1BWP30P140LVT U2006 ( .A1(i_data_bus[784]), .A2(n1946), .B1(
        i_data_bus[816]), .B2(n1943), .ZN(n1623) );
  ND4D1BWP30P140LVT U2007 ( .A1(n1626), .A2(n1625), .A3(n1624), .A4(n1623), 
        .ZN(n1627) );
  OR4D1BWP30P140LVT U2008 ( .A1(n1630), .A2(n1629), .A3(n1628), .A4(n1627), 
        .Z(o_data_bus[112]) );
  AOI22D1BWP30P140LVT U2009 ( .A1(i_data_bus[1009]), .A2(n1934), .B1(
        i_data_bus[593]), .B2(n1912), .ZN(n1634) );
  AOI22D1BWP30P140LVT U2010 ( .A1(i_data_bus[305]), .A2(n1922), .B1(
        i_data_bus[497]), .B2(n1932), .ZN(n1633) );
  AOI22D1BWP30P140LVT U2011 ( .A1(i_data_bus[113]), .A2(n1936), .B1(
        i_data_bus[273]), .B2(n1293), .ZN(n1632) );
  AOI22D1BWP30P140LVT U2012 ( .A1(i_data_bus[561]), .A2(n1924), .B1(
        i_data_bus[241]), .B2(n1911), .ZN(n1631) );
  ND4D1BWP30P140LVT U2013 ( .A1(n1634), .A2(n1633), .A3(n1632), .A4(n1631), 
        .ZN(n1650) );
  AOI22D1BWP30P140LVT U2014 ( .A1(i_data_bus[81]), .A2(n1925), .B1(
        i_data_bus[945]), .B2(n127), .ZN(n1638) );
  AOI22D1BWP30P140LVT U2015 ( .A1(i_data_bus[401]), .A2(n1279), .B1(
        i_data_bus[209]), .B2(n1916), .ZN(n1637) );
  AOI22D1BWP30P140LVT U2016 ( .A1(i_data_bus[977]), .A2(n1923), .B1(
        i_data_bus[433]), .B2(n1921), .ZN(n1636) );
  AOI22D1BWP30P140LVT U2017 ( .A1(i_data_bus[49]), .A2(n1914), .B1(
        i_data_bus[913]), .B2(n128), .ZN(n1635) );
  ND4D1BWP30P140LVT U2018 ( .A1(n1638), .A2(n1637), .A3(n1636), .A4(n1635), 
        .ZN(n1649) );
  AOI22D1BWP30P140LVT U2019 ( .A1(i_data_bus[145]), .A2(n1935), .B1(
        i_data_bus[177]), .B2(n1915), .ZN(n1642) );
  AOI22D1BWP30P140LVT U2020 ( .A1(i_data_bus[17]), .A2(n2), .B1(
        i_data_bus[465]), .B2(n1933), .ZN(n1641) );
  AOI22D1BWP30P140LVT U2021 ( .A1(i_data_bus[625]), .A2(n1910), .B1(
        i_data_bus[529]), .B2(n1927), .ZN(n1640) );
  AOI22D1BWP30P140LVT U2022 ( .A1(i_data_bus[337]), .A2(n1913), .B1(
        i_data_bus[369]), .B2(n1926), .ZN(n1639) );
  ND4D1BWP30P140LVT U2023 ( .A1(n1642), .A2(n1641), .A3(n1640), .A4(n1639), 
        .ZN(n1648) );
  AOI22D1BWP30P140LVT U2024 ( .A1(i_data_bus[881]), .A2(n1941), .B1(
        i_data_bus[817]), .B2(n1943), .ZN(n1646) );
  AOI22D1BWP30P140LVT U2025 ( .A1(i_data_bus[785]), .A2(n1946), .B1(
        i_data_bus[657]), .B2(n1944), .ZN(n1645) );
  AOI22D1BWP30P140LVT U2026 ( .A1(i_data_bus[689]), .A2(n1947), .B1(
        i_data_bus[753]), .B2(n1945), .ZN(n1644) );
  AOI22D1BWP30P140LVT U2027 ( .A1(i_data_bus[849]), .A2(n1948), .B1(
        i_data_bus[721]), .B2(n1942), .ZN(n1643) );
  ND4D1BWP30P140LVT U2028 ( .A1(n1646), .A2(n1645), .A3(n1644), .A4(n1643), 
        .ZN(n1647) );
  OR4D1BWP30P140LVT U2029 ( .A1(n1650), .A2(n1649), .A3(n1648), .A4(n1647), 
        .Z(o_data_bus[113]) );
  AOI22D1BWP30P140LVT U2030 ( .A1(i_data_bus[402]), .A2(n1279), .B1(
        i_data_bus[146]), .B2(n1935), .ZN(n1654) );
  AOI22D1BWP30P140LVT U2031 ( .A1(i_data_bus[242]), .A2(n1911), .B1(
        i_data_bus[210]), .B2(n1916), .ZN(n1653) );
  AOI22D1BWP30P140LVT U2032 ( .A1(i_data_bus[594]), .A2(n1912), .B1(
        i_data_bus[466]), .B2(n1933), .ZN(n1651) );
  ND4D1BWP30P140LVT U2033 ( .A1(n1654), .A2(n1653), .A3(n1652), .A4(n1651), 
        .ZN(n1670) );
  AOI22D1BWP30P140LVT U2034 ( .A1(i_data_bus[626]), .A2(n1910), .B1(
        i_data_bus[178]), .B2(n1915), .ZN(n1658) );
  AOI22D1BWP30P140LVT U2035 ( .A1(i_data_bus[914]), .A2(n128), .B1(
        i_data_bus[370]), .B2(n1926), .ZN(n1657) );
  AOI22D1BWP30P140LVT U2036 ( .A1(i_data_bus[562]), .A2(n1924), .B1(
        i_data_bus[338]), .B2(n1913), .ZN(n1656) );
  AOI22D1BWP30P140LVT U2037 ( .A1(i_data_bus[50]), .A2(n1914), .B1(
        i_data_bus[498]), .B2(n1932), .ZN(n1655) );
  ND4D1BWP30P140LVT U2038 ( .A1(n1658), .A2(n1657), .A3(n1656), .A4(n1655), 
        .ZN(n1669) );
  AOI22D1BWP30P140LVT U2039 ( .A1(i_data_bus[978]), .A2(n1923), .B1(
        i_data_bus[1010]), .B2(n1934), .ZN(n1662) );
  AOI22D1BWP30P140LVT U2040 ( .A1(i_data_bus[274]), .A2(n1293), .B1(
        i_data_bus[434]), .B2(n1921), .ZN(n1661) );
  AOI22D1BWP30P140LVT U2041 ( .A1(i_data_bus[18]), .A2(n2), .B1(
        i_data_bus[306]), .B2(n1922), .ZN(n1660) );
  AOI22D1BWP30P140LVT U2042 ( .A1(i_data_bus[114]), .A2(n1936), .B1(
        i_data_bus[946]), .B2(n127), .ZN(n1659) );
  ND4D1BWP30P140LVT U2043 ( .A1(n1662), .A2(n1661), .A3(n1660), .A4(n1659), 
        .ZN(n1668) );
  AOI22D1BWP30P140LVT U2044 ( .A1(i_data_bus[882]), .A2(n1941), .B1(
        i_data_bus[850]), .B2(n1948), .ZN(n1666) );
  AOI22D1BWP30P140LVT U2045 ( .A1(i_data_bus[722]), .A2(n1942), .B1(
        i_data_bus[818]), .B2(n1943), .ZN(n1665) );
  AOI22D1BWP30P140LVT U2046 ( .A1(i_data_bus[690]), .A2(n1947), .B1(
        i_data_bus[754]), .B2(n1945), .ZN(n1664) );
  AOI22D1BWP30P140LVT U2047 ( .A1(i_data_bus[658]), .A2(n1944), .B1(
        i_data_bus[786]), .B2(n1946), .ZN(n1663) );
  ND4D1BWP30P140LVT U2048 ( .A1(n1666), .A2(n1665), .A3(n1664), .A4(n1663), 
        .ZN(n1667) );
  OR4D1BWP30P140LVT U2049 ( .A1(n1670), .A2(n1669), .A3(n1668), .A4(n1667), 
        .Z(o_data_bus[114]) );
  AOI22D1BWP30P140LVT U2050 ( .A1(i_data_bus[147]), .A2(n1935), .B1(
        i_data_bus[275]), .B2(n1293), .ZN(n1674) );
  AOI22D1BWP30P140LVT U2051 ( .A1(i_data_bus[595]), .A2(n1912), .B1(
        i_data_bus[179]), .B2(n1915), .ZN(n1673) );
  AOI22D1BWP30P140LVT U2052 ( .A1(i_data_bus[339]), .A2(n1913), .B1(
        i_data_bus[435]), .B2(n1921), .ZN(n1672) );
  AOI22D1BWP30P140LVT U2053 ( .A1(i_data_bus[1011]), .A2(n1934), .B1(
        i_data_bus[947]), .B2(n127), .ZN(n1671) );
  ND4D1BWP30P140LVT U2054 ( .A1(n1674), .A2(n1673), .A3(n1672), .A4(n1671), 
        .ZN(n1690) );
  AOI22D1BWP30P140LVT U2055 ( .A1(i_data_bus[979]), .A2(n1923), .B1(
        i_data_bus[211]), .B2(n1916), .ZN(n1678) );
  AOI22D1BWP30P140LVT U2056 ( .A1(i_data_bus[83]), .A2(n1925), .B1(
        i_data_bus[915]), .B2(n128), .ZN(n1677) );
  AOI22D1BWP30P140LVT U2057 ( .A1(i_data_bus[627]), .A2(n1910), .B1(
        i_data_bus[371]), .B2(n1926), .ZN(n1676) );
  AOI22D1BWP30P140LVT U2058 ( .A1(i_data_bus[307]), .A2(n1922), .B1(
        i_data_bus[403]), .B2(n1279), .ZN(n1675) );
  ND4D1BWP30P140LVT U2059 ( .A1(n1678), .A2(n1677), .A3(n1676), .A4(n1675), 
        .ZN(n1689) );
  AOI22D1BWP30P140LVT U2060 ( .A1(i_data_bus[563]), .A2(n1924), .B1(
        i_data_bus[531]), .B2(n1927), .ZN(n1682) );
  AOI22D1BWP30P140LVT U2061 ( .A1(i_data_bus[243]), .A2(n1911), .B1(
        i_data_bus[467]), .B2(n1933), .ZN(n1681) );
  AOI22D1BWP30P140LVT U2062 ( .A1(i_data_bus[51]), .A2(n1914), .B1(
        i_data_bus[115]), .B2(n1936), .ZN(n1680) );
  AOI22D1BWP30P140LVT U2063 ( .A1(i_data_bus[19]), .A2(n2), .B1(
        i_data_bus[499]), .B2(n1932), .ZN(n1679) );
  ND4D1BWP30P140LVT U2064 ( .A1(n1680), .A2(n1681), .A3(n1682), .A4(n1679), 
        .ZN(n1688) );
  AOI22D1BWP30P140LVT U2065 ( .A1(i_data_bus[883]), .A2(n1941), .B1(
        i_data_bus[851]), .B2(n1948), .ZN(n1686) );
  AOI22D1BWP30P140LVT U2066 ( .A1(i_data_bus[819]), .A2(n1943), .B1(
        i_data_bus[787]), .B2(n1946), .ZN(n1685) );
  AOI22D1BWP30P140LVT U2067 ( .A1(i_data_bus[755]), .A2(n1945), .B1(
        i_data_bus[659]), .B2(n1944), .ZN(n1684) );
  AOI22D1BWP30P140LVT U2068 ( .A1(i_data_bus[691]), .A2(n1947), .B1(
        i_data_bus[723]), .B2(n1942), .ZN(n1683) );
  ND4D1BWP30P140LVT U2069 ( .A1(n1686), .A2(n1685), .A3(n1684), .A4(n1683), 
        .ZN(n1687) );
  OR4D1BWP30P140LVT U2070 ( .A1(n1690), .A2(n1689), .A3(n1687), .A4(n1688), 
        .Z(o_data_bus[115]) );
  AOI22D1BWP30P140LVT U2071 ( .A1(i_data_bus[916]), .A2(n128), .B1(
        i_data_bus[276]), .B2(n1293), .ZN(n1694) );
  AOI22D1BWP30P140LVT U2072 ( .A1(i_data_bus[980]), .A2(n1923), .B1(
        i_data_bus[436]), .B2(n1921), .ZN(n1693) );
  AOI22D1BWP30P140LVT U2073 ( .A1(i_data_bus[340]), .A2(n1913), .B1(
        i_data_bus[468]), .B2(n1933), .ZN(n1692) );
  AOI22D1BWP30P140LVT U2074 ( .A1(i_data_bus[116]), .A2(n1936), .B1(
        i_data_bus[404]), .B2(n1279), .ZN(n1691) );
  ND4D1BWP30P140LVT U2075 ( .A1(n1694), .A2(n1693), .A3(n1692), .A4(n1691), 
        .ZN(n1710) );
  AOI22D1BWP30P140LVT U2076 ( .A1(i_data_bus[20]), .A2(n2), .B1(
        i_data_bus[180]), .B2(n1915), .ZN(n1698) );
  AOI22D1BWP30P140LVT U2077 ( .A1(i_data_bus[564]), .A2(n1924), .B1(
        i_data_bus[212]), .B2(n1916), .ZN(n1697) );
  AOI22D1BWP30P140LVT U2078 ( .A1(i_data_bus[628]), .A2(n1910), .B1(
        i_data_bus[948]), .B2(n127), .ZN(n1696) );
  AOI22D1BWP30P140LVT U2079 ( .A1(i_data_bus[84]), .A2(n1925), .B1(
        i_data_bus[372]), .B2(n1926), .ZN(n1695) );
  ND4D1BWP30P140LVT U2080 ( .A1(n1698), .A2(n1697), .A3(n1696), .A4(n1695), 
        .ZN(n1709) );
  AOI22D1BWP30P140LVT U2081 ( .A1(i_data_bus[244]), .A2(n1911), .B1(
        i_data_bus[148]), .B2(n1935), .ZN(n1702) );
  AOI22D1BWP30P140LVT U2082 ( .A1(i_data_bus[532]), .A2(n1927), .B1(
        i_data_bus[308]), .B2(n1922), .ZN(n1701) );
  AOI22D1BWP30P140LVT U2083 ( .A1(i_data_bus[52]), .A2(n1914), .B1(
        i_data_bus[1012]), .B2(n1934), .ZN(n1700) );
  AOI22D1BWP30P140LVT U2084 ( .A1(i_data_bus[596]), .A2(n1912), .B1(
        i_data_bus[500]), .B2(n1932), .ZN(n1699) );
  ND4D1BWP30P140LVT U2085 ( .A1(n1702), .A2(n1701), .A3(n1700), .A4(n1699), 
        .ZN(n1708) );
  AOI22D1BWP30P140LVT U2086 ( .A1(i_data_bus[756]), .A2(n1945), .B1(
        i_data_bus[884]), .B2(n1941), .ZN(n1706) );
  AOI22D1BWP30P140LVT U2087 ( .A1(i_data_bus[660]), .A2(n1944), .B1(
        i_data_bus[692]), .B2(n1947), .ZN(n1705) );
  AOI22D1BWP30P140LVT U2088 ( .A1(i_data_bus[724]), .A2(n1942), .B1(
        i_data_bus[820]), .B2(n1943), .ZN(n1704) );
  AOI22D1BWP30P140LVT U2089 ( .A1(i_data_bus[788]), .A2(n1946), .B1(
        i_data_bus[852]), .B2(n1948), .ZN(n1703) );
  ND4D1BWP30P140LVT U2090 ( .A1(n1706), .A2(n1705), .A3(n1704), .A4(n1703), 
        .ZN(n1707) );
  OR4D1BWP30P140LVT U2091 ( .A1(n1710), .A2(n1709), .A3(n1708), .A4(n1707), 
        .Z(o_data_bus[116]) );
  AOI22D1BWP30P140LVT U2092 ( .A1(i_data_bus[533]), .A2(n1927), .B1(
        i_data_bus[373]), .B2(n1926), .ZN(n1714) );
  AOI22D1BWP30P140LVT U2093 ( .A1(i_data_bus[1013]), .A2(n1934), .B1(
        i_data_bus[469]), .B2(n1933), .ZN(n1713) );
  AOI22D1BWP30P140LVT U2094 ( .A1(i_data_bus[181]), .A2(n1915), .B1(
        i_data_bus[501]), .B2(n1932), .ZN(n1712) );
  AOI22D1BWP30P140LVT U2095 ( .A1(i_data_bus[277]), .A2(n1293), .B1(
        i_data_bus[405]), .B2(n1279), .ZN(n1711) );
  ND4D1BWP30P140LVT U2096 ( .A1(n1714), .A2(n1713), .A3(n1712), .A4(n1711), 
        .ZN(n1730) );
  AOI22D1BWP30P140LVT U2097 ( .A1(i_data_bus[213]), .A2(n1916), .B1(
        i_data_bus[245]), .B2(n1911), .ZN(n1718) );
  AOI22D1BWP30P140LVT U2098 ( .A1(i_data_bus[917]), .A2(n128), .B1(
        i_data_bus[21]), .B2(n2), .ZN(n1717) );
  AOI22D1BWP30P140LVT U2099 ( .A1(i_data_bus[117]), .A2(n1936), .B1(
        i_data_bus[149]), .B2(n1935), .ZN(n1715) );
  ND4D1BWP30P140LVT U2100 ( .A1(n1716), .A2(n1717), .A3(n1718), .A4(n1715), 
        .ZN(n1729) );
  AOI22D1BWP30P140LVT U2101 ( .A1(i_data_bus[53]), .A2(n1914), .B1(
        i_data_bus[341]), .B2(n1913), .ZN(n1722) );
  AOI22D1BWP30P140LVT U2102 ( .A1(i_data_bus[949]), .A2(n127), .B1(
        i_data_bus[981]), .B2(n1923), .ZN(n1721) );
  AOI22D1BWP30P140LVT U2103 ( .A1(i_data_bus[597]), .A2(n1912), .B1(
        i_data_bus[309]), .B2(n1922), .ZN(n1720) );
  AOI22D1BWP30P140LVT U2104 ( .A1(i_data_bus[565]), .A2(n1924), .B1(
        i_data_bus[437]), .B2(n1921), .ZN(n1719) );
  ND4D1BWP30P140LVT U2105 ( .A1(n1722), .A2(n1721), .A3(n1720), .A4(n1719), 
        .ZN(n1728) );
  AOI22D1BWP30P140LVT U2106 ( .A1(i_data_bus[789]), .A2(n1946), .B1(
        i_data_bus[725]), .B2(n1942), .ZN(n1726) );
  AOI22D1BWP30P140LVT U2107 ( .A1(i_data_bus[821]), .A2(n1943), .B1(
        i_data_bus[693]), .B2(n1947), .ZN(n1725) );
  AOI22D1BWP30P140LVT U2108 ( .A1(i_data_bus[757]), .A2(n1945), .B1(
        i_data_bus[853]), .B2(n1948), .ZN(n1724) );
  AOI22D1BWP30P140LVT U2109 ( .A1(i_data_bus[661]), .A2(n1944), .B1(
        i_data_bus[885]), .B2(n1941), .ZN(n1723) );
  ND4D1BWP30P140LVT U2110 ( .A1(n1726), .A2(n1725), .A3(n1724), .A4(n1723), 
        .ZN(n1727) );
  OR4D1BWP30P140LVT U2111 ( .A1(n1730), .A2(n1729), .A3(n1728), .A4(n1727), 
        .Z(o_data_bus[117]) );
  AOI22D1BWP30P140LVT U2112 ( .A1(i_data_bus[502]), .A2(n1932), .B1(
        i_data_bus[214]), .B2(n1916), .ZN(n1734) );
  AOI22D1BWP30P140LVT U2113 ( .A1(i_data_bus[406]), .A2(n1279), .B1(
        i_data_bus[342]), .B2(n1913), .ZN(n1733) );
  AOI22D1BWP30P140LVT U2114 ( .A1(i_data_bus[150]), .A2(n1935), .B1(
        i_data_bus[278]), .B2(n1293), .ZN(n1732) );
  AOI22D1BWP30P140LVT U2115 ( .A1(i_data_bus[630]), .A2(n1910), .B1(
        i_data_bus[982]), .B2(n1923), .ZN(n1731) );
  ND4D1BWP30P140LVT U2116 ( .A1(n1734), .A2(n1733), .A3(n1732), .A4(n1731), 
        .ZN(n1750) );
  AOI22D1BWP30P140LVT U2117 ( .A1(i_data_bus[118]), .A2(n1936), .B1(
        i_data_bus[950]), .B2(n127), .ZN(n1738) );
  AOI22D1BWP30P140LVT U2118 ( .A1(i_data_bus[1014]), .A2(n1934), .B1(
        i_data_bus[534]), .B2(n1927), .ZN(n1736) );
  AOI22D1BWP30P140LVT U2119 ( .A1(i_data_bus[566]), .A2(n1924), .B1(
        i_data_bus[374]), .B2(n1926), .ZN(n1735) );
  ND4D1BWP30P140LVT U2120 ( .A1(n1738), .A2(n1737), .A3(n1736), .A4(n1735), 
        .ZN(n1749) );
  AOI22D1BWP30P140LVT U2121 ( .A1(i_data_bus[54]), .A2(n1914), .B1(
        i_data_bus[438]), .B2(n1921), .ZN(n1742) );
  AOI22D1BWP30P140LVT U2122 ( .A1(i_data_bus[22]), .A2(n2), .B1(
        i_data_bus[470]), .B2(n1933), .ZN(n1741) );
  AOI22D1BWP30P140LVT U2123 ( .A1(i_data_bus[246]), .A2(n1911), .B1(
        i_data_bus[182]), .B2(n1915), .ZN(n1740) );
  AOI22D1BWP30P140LVT U2124 ( .A1(i_data_bus[918]), .A2(n128), .B1(
        i_data_bus[310]), .B2(n1922), .ZN(n1739) );
  ND4D1BWP30P140LVT U2125 ( .A1(n1742), .A2(n1741), .A3(n1740), .A4(n1739), 
        .ZN(n1748) );
  AOI22D1BWP30P140LVT U2126 ( .A1(i_data_bus[694]), .A2(n1947), .B1(
        i_data_bus[758]), .B2(n1945), .ZN(n1746) );
  AOI22D1BWP30P140LVT U2127 ( .A1(i_data_bus[726]), .A2(n1942), .B1(
        i_data_bus[854]), .B2(n1948), .ZN(n1745) );
  AOI22D1BWP30P140LVT U2128 ( .A1(i_data_bus[886]), .A2(n1941), .B1(
        i_data_bus[662]), .B2(n1944), .ZN(n1744) );
  AOI22D1BWP30P140LVT U2129 ( .A1(i_data_bus[822]), .A2(n1943), .B1(
        i_data_bus[790]), .B2(n1946), .ZN(n1743) );
  ND4D1BWP30P140LVT U2130 ( .A1(n1746), .A2(n1745), .A3(n1744), .A4(n1743), 
        .ZN(n1747) );
  OR4D1BWP30P140LVT U2131 ( .A1(n1750), .A2(n1749), .A3(n1748), .A4(n1747), 
        .Z(o_data_bus[118]) );
  AOI22D1BWP30P140LVT U2132 ( .A1(i_data_bus[471]), .A2(n1933), .B1(
        i_data_bus[439]), .B2(n1921), .ZN(n1754) );
  AOI22D1BWP30P140LVT U2133 ( .A1(i_data_bus[311]), .A2(n1922), .B1(
        i_data_bus[279]), .B2(n1293), .ZN(n1753) );
  AOI22D1BWP30P140LVT U2134 ( .A1(i_data_bus[599]), .A2(n1912), .B1(
        i_data_bus[343]), .B2(n1913), .ZN(n1751) );
  ND4D1BWP30P140LVT U2135 ( .A1(n1754), .A2(n1753), .A3(n1752), .A4(n1751), 
        .ZN(n1770) );
  AOI22D1BWP30P140LVT U2136 ( .A1(i_data_bus[247]), .A2(n1911), .B1(
        i_data_bus[375]), .B2(n1926), .ZN(n1758) );
  AOI22D1BWP30P140LVT U2137 ( .A1(i_data_bus[119]), .A2(n1936), .B1(
        i_data_bus[567]), .B2(n1924), .ZN(n1757) );
  AOI22D1BWP30P140LVT U2138 ( .A1(i_data_bus[151]), .A2(n1935), .B1(
        i_data_bus[407]), .B2(n1279), .ZN(n1756) );
  AOI22D1BWP30P140LVT U2139 ( .A1(i_data_bus[951]), .A2(n127), .B1(
        i_data_bus[919]), .B2(n128), .ZN(n1755) );
  ND4D1BWP30P140LVT U2140 ( .A1(n1758), .A2(n1757), .A3(n1756), .A4(n1755), 
        .ZN(n1769) );
  AOI22D1BWP30P140LVT U2141 ( .A1(i_data_bus[23]), .A2(n2), .B1(
        i_data_bus[535]), .B2(n1927), .ZN(n1762) );
  AOI22D1BWP30P140LVT U2142 ( .A1(i_data_bus[983]), .A2(n1923), .B1(
        i_data_bus[215]), .B2(n1916), .ZN(n1761) );
  AOI22D1BWP30P140LVT U2143 ( .A1(i_data_bus[631]), .A2(n1910), .B1(
        i_data_bus[183]), .B2(n1915), .ZN(n1760) );
  AOI22D1BWP30P140LVT U2144 ( .A1(i_data_bus[55]), .A2(n1914), .B1(
        i_data_bus[503]), .B2(n1932), .ZN(n1759) );
  ND4D1BWP30P140LVT U2145 ( .A1(n1762), .A2(n1761), .A3(n1760), .A4(n1759), 
        .ZN(n1768) );
  AOI22D1BWP30P140LVT U2146 ( .A1(i_data_bus[887]), .A2(n1941), .B1(
        i_data_bus[663]), .B2(n1944), .ZN(n1766) );
  AOI22D1BWP30P140LVT U2147 ( .A1(i_data_bus[759]), .A2(n1945), .B1(
        i_data_bus[855]), .B2(n1948), .ZN(n1765) );
  AOI22D1BWP30P140LVT U2148 ( .A1(i_data_bus[727]), .A2(n1942), .B1(
        i_data_bus[823]), .B2(n1943), .ZN(n1764) );
  AOI22D1BWP30P140LVT U2149 ( .A1(i_data_bus[695]), .A2(n1947), .B1(
        i_data_bus[791]), .B2(n1946), .ZN(n1763) );
  ND4D1BWP30P140LVT U2150 ( .A1(n1766), .A2(n1765), .A3(n1764), .A4(n1763), 
        .ZN(n1767) );
  OR4D1BWP30P140LVT U2151 ( .A1(n1770), .A2(n1769), .A3(n1768), .A4(n1767), 
        .Z(o_data_bus[119]) );
  AOI22D1BWP30P140LVT U2152 ( .A1(i_data_bus[600]), .A2(n1912), .B1(
        i_data_bus[952]), .B2(n127), .ZN(n1774) );
  AOI22D1BWP30P140LVT U2153 ( .A1(i_data_bus[536]), .A2(n1927), .B1(
        i_data_bus[248]), .B2(n1911), .ZN(n1773) );
  AOI22D1BWP30P140LVT U2154 ( .A1(i_data_bus[920]), .A2(n128), .B1(
        i_data_bus[376]), .B2(n1926), .ZN(n1772) );
  AOI22D1BWP30P140LVT U2155 ( .A1(i_data_bus[88]), .A2(n1925), .B1(
        i_data_bus[344]), .B2(n1913), .ZN(n1771) );
  ND4D1BWP30P140LVT U2156 ( .A1(n1774), .A2(n1773), .A3(n1772), .A4(n1771), 
        .ZN(n1790) );
  AOI22D1BWP30P140LVT U2157 ( .A1(i_data_bus[56]), .A2(n1914), .B1(
        i_data_bus[216]), .B2(n1916), .ZN(n1778) );
  AOI22D1BWP30P140LVT U2158 ( .A1(i_data_bus[440]), .A2(n1921), .B1(
        i_data_bus[152]), .B2(n1935), .ZN(n1777) );
  AOI22D1BWP30P140LVT U2159 ( .A1(i_data_bus[280]), .A2(n1293), .B1(
        i_data_bus[504]), .B2(n1932), .ZN(n1776) );
  AOI22D1BWP30P140LVT U2160 ( .A1(i_data_bus[1016]), .A2(n1934), .B1(
        i_data_bus[184]), .B2(n1915), .ZN(n1775) );
  ND4D1BWP30P140LVT U2161 ( .A1(n1778), .A2(n1777), .A3(n1776), .A4(n1775), 
        .ZN(n1789) );
  AOI22D1BWP30P140LVT U2162 ( .A1(i_data_bus[24]), .A2(n2), .B1(
        i_data_bus[568]), .B2(n1924), .ZN(n1782) );
  AOI22D1BWP30P140LVT U2163 ( .A1(i_data_bus[984]), .A2(n1923), .B1(
        i_data_bus[472]), .B2(n1933), .ZN(n1781) );
  AOI22D1BWP30P140LVT U2164 ( .A1(i_data_bus[632]), .A2(n1910), .B1(
        i_data_bus[408]), .B2(n1279), .ZN(n1780) );
  AOI22D1BWP30P140LVT U2165 ( .A1(i_data_bus[120]), .A2(n1936), .B1(
        i_data_bus[312]), .B2(n1922), .ZN(n1779) );
  ND4D1BWP30P140LVT U2166 ( .A1(n1782), .A2(n1781), .A3(n1780), .A4(n1779), 
        .ZN(n1788) );
  AOI22D1BWP30P140LVT U2167 ( .A1(i_data_bus[824]), .A2(n1943), .B1(
        i_data_bus[760]), .B2(n1945), .ZN(n1786) );
  AOI22D1BWP30P140LVT U2168 ( .A1(i_data_bus[856]), .A2(n1948), .B1(
        i_data_bus[664]), .B2(n1944), .ZN(n1785) );
  AOI22D1BWP30P140LVT U2169 ( .A1(i_data_bus[728]), .A2(n1942), .B1(
        i_data_bus[888]), .B2(n1941), .ZN(n1784) );
  AOI22D1BWP30P140LVT U2170 ( .A1(i_data_bus[792]), .A2(n1946), .B1(
        i_data_bus[696]), .B2(n1947), .ZN(n1783) );
  ND4D1BWP30P140LVT U2171 ( .A1(n1786), .A2(n1785), .A3(n1784), .A4(n1783), 
        .ZN(n1787) );
  OR4D1BWP30P140LVT U2172 ( .A1(n1790), .A2(n1789), .A3(n1788), .A4(n1787), 
        .Z(o_data_bus[120]) );
  AOI22D1BWP30P140LVT U2173 ( .A1(i_data_bus[345]), .A2(n1913), .B1(
        i_data_bus[441]), .B2(n1921), .ZN(n1793) );
  AOI22D1BWP30P140LVT U2174 ( .A1(i_data_bus[1017]), .A2(n1934), .B1(
        i_data_bus[313]), .B2(n1922), .ZN(n1792) );
  AOI22D1BWP30P140LVT U2175 ( .A1(i_data_bus[921]), .A2(n128), .B1(
        i_data_bus[121]), .B2(n1936), .ZN(n1791) );
  AOI22D1BWP30P140LVT U2176 ( .A1(i_data_bus[89]), .A2(n1925), .B1(
        i_data_bus[217]), .B2(n1916), .ZN(n1797) );
  AOI22D1BWP30P140LVT U2177 ( .A1(i_data_bus[953]), .A2(n127), .B1(
        i_data_bus[185]), .B2(n1915), .ZN(n1796) );
  AOI22D1BWP30P140LVT U2178 ( .A1(i_data_bus[57]), .A2(n1914), .B1(
        i_data_bus[601]), .B2(n1912), .ZN(n1795) );
  AOI22D1BWP30P140LVT U2179 ( .A1(i_data_bus[537]), .A2(n1927), .B1(
        i_data_bus[153]), .B2(n1935), .ZN(n1794) );
  ND4D1BWP30P140LVT U2180 ( .A1(n1797), .A2(n1796), .A3(n1795), .A4(n1794), 
        .ZN(n1808) );
  AOI22D1BWP30P140LVT U2181 ( .A1(i_data_bus[377]), .A2(n1926), .B1(
        i_data_bus[505]), .B2(n1932), .ZN(n1801) );
  AOI22D1BWP30P140LVT U2182 ( .A1(i_data_bus[633]), .A2(n1910), .B1(
        i_data_bus[473]), .B2(n1933), .ZN(n1800) );
  AOI22D1BWP30P140LVT U2183 ( .A1(i_data_bus[985]), .A2(n1923), .B1(
        i_data_bus[25]), .B2(n2), .ZN(n1799) );
  AOI22D1BWP30P140LVT U2184 ( .A1(i_data_bus[569]), .A2(n1924), .B1(
        i_data_bus[409]), .B2(n1279), .ZN(n1798) );
  ND4D1BWP30P140LVT U2185 ( .A1(n1801), .A2(n1800), .A3(n1799), .A4(n1798), 
        .ZN(n1807) );
  AOI22D1BWP30P140LVT U2186 ( .A1(i_data_bus[825]), .A2(n1943), .B1(
        i_data_bus[793]), .B2(n1946), .ZN(n1805) );
  AOI22D1BWP30P140LVT U2187 ( .A1(i_data_bus[761]), .A2(n1945), .B1(
        i_data_bus[857]), .B2(n1948), .ZN(n1804) );
  AOI22D1BWP30P140LVT U2188 ( .A1(i_data_bus[729]), .A2(n1942), .B1(
        i_data_bus[665]), .B2(n1944), .ZN(n1803) );
  AOI22D1BWP30P140LVT U2189 ( .A1(i_data_bus[697]), .A2(n1947), .B1(
        i_data_bus[889]), .B2(n1941), .ZN(n1802) );
  ND4D1BWP30P140LVT U2190 ( .A1(n1805), .A2(n1804), .A3(n1803), .A4(n1802), 
        .ZN(n1806) );
  OR4D1BWP30P140LVT U2191 ( .A1(n1807), .A2(n1808), .A3(n1809), .A4(n1806), 
        .Z(o_data_bus[121]) );
  AOI22D1BWP30P140LVT U2192 ( .A1(i_data_bus[634]), .A2(n1910), .B1(
        i_data_bus[314]), .B2(n1922), .ZN(n1813) );
  AOI22D1BWP30P140LVT U2193 ( .A1(i_data_bus[954]), .A2(n127), .B1(
        i_data_bus[506]), .B2(n1932), .ZN(n1812) );
  AOI22D1BWP30P140LVT U2194 ( .A1(i_data_bus[442]), .A2(n1921), .B1(
        i_data_bus[378]), .B2(n1926), .ZN(n1811) );
  AOI22D1BWP30P140LVT U2195 ( .A1(i_data_bus[570]), .A2(n1924), .B1(
        i_data_bus[218]), .B2(n1916), .ZN(n1810) );
  ND4D1BWP30P140LVT U2196 ( .A1(n1813), .A2(n1812), .A3(n1811), .A4(n1810), 
        .ZN(n1829) );
  AOI22D1BWP30P140LVT U2197 ( .A1(i_data_bus[90]), .A2(n1925), .B1(
        i_data_bus[474]), .B2(n1933), .ZN(n1817) );
  AOI22D1BWP30P140LVT U2198 ( .A1(i_data_bus[122]), .A2(n1936), .B1(
        i_data_bus[538]), .B2(n1927), .ZN(n1816) );
  AOI22D1BWP30P140LVT U2199 ( .A1(i_data_bus[602]), .A2(n1912), .B1(
        i_data_bus[986]), .B2(n1923), .ZN(n1815) );
  AOI22D1BWP30P140LVT U2200 ( .A1(i_data_bus[58]), .A2(n1914), .B1(
        i_data_bus[186]), .B2(n1915), .ZN(n1814) );
  ND4D1BWP30P140LVT U2201 ( .A1(n1817), .A2(n1816), .A3(n1815), .A4(n1814), 
        .ZN(n1828) );
  AOI22D1BWP30P140LVT U2202 ( .A1(i_data_bus[26]), .A2(n2), .B1(
        i_data_bus[346]), .B2(n1913), .ZN(n1821) );
  AOI22D1BWP30P140LVT U2203 ( .A1(i_data_bus[922]), .A2(n128), .B1(
        i_data_bus[282]), .B2(n1293), .ZN(n1820) );
  AOI22D1BWP30P140LVT U2204 ( .A1(i_data_bus[1018]), .A2(n1934), .B1(
        i_data_bus[154]), .B2(n1935), .ZN(n1819) );
  AOI22D1BWP30P140LVT U2205 ( .A1(i_data_bus[250]), .A2(n1911), .B1(
        i_data_bus[410]), .B2(n1279), .ZN(n1818) );
  ND4D1BWP30P140LVT U2206 ( .A1(n1821), .A2(n1820), .A3(n1819), .A4(n1818), 
        .ZN(n1827) );
  AOI22D1BWP30P140LVT U2207 ( .A1(i_data_bus[858]), .A2(n1948), .B1(
        i_data_bus[762]), .B2(n1945), .ZN(n1825) );
  AOI22D1BWP30P140LVT U2208 ( .A1(i_data_bus[826]), .A2(n1943), .B1(
        i_data_bus[730]), .B2(n1942), .ZN(n1824) );
  AOI22D1BWP30P140LVT U2209 ( .A1(i_data_bus[890]), .A2(n1941), .B1(
        i_data_bus[698]), .B2(n1947), .ZN(n1823) );
  AOI22D1BWP30P140LVT U2210 ( .A1(i_data_bus[794]), .A2(n1946), .B1(
        i_data_bus[666]), .B2(n1944), .ZN(n1822) );
  ND4D1BWP30P140LVT U2211 ( .A1(n1825), .A2(n1824), .A3(n1823), .A4(n1822), 
        .ZN(n1826) );
  OR4D1BWP30P140LVT U2212 ( .A1(n1829), .A2(n1828), .A3(n1827), .A4(n1826), 
        .Z(o_data_bus[122]) );
  AOI22D1BWP30P140LVT U2213 ( .A1(i_data_bus[603]), .A2(n1912), .B1(
        i_data_bus[923]), .B2(n128), .ZN(n1833) );
  AOI22D1BWP30P140LVT U2214 ( .A1(i_data_bus[411]), .A2(n1279), .B1(
        i_data_bus[283]), .B2(n1293), .ZN(n1832) );
  AOI22D1BWP30P140LVT U2215 ( .A1(i_data_bus[123]), .A2(n1936), .B1(
        i_data_bus[475]), .B2(n1933), .ZN(n1831) );
  AOI22D1BWP30P140LVT U2216 ( .A1(i_data_bus[987]), .A2(n1923), .B1(
        i_data_bus[347]), .B2(n1913), .ZN(n1830) );
  ND4D1BWP30P140LVT U2217 ( .A1(n1833), .A2(n1832), .A3(n1831), .A4(n1830), 
        .ZN(n1849) );
  AOI22D1BWP30P140LVT U2218 ( .A1(i_data_bus[635]), .A2(n1910), .B1(
        i_data_bus[219]), .B2(n1916), .ZN(n1837) );
  AOI22D1BWP30P140LVT U2219 ( .A1(i_data_bus[1019]), .A2(n1934), .B1(
        i_data_bus[155]), .B2(n1935), .ZN(n1836) );
  AOI22D1BWP30P140LVT U2220 ( .A1(i_data_bus[91]), .A2(n1925), .B1(
        i_data_bus[379]), .B2(n1926), .ZN(n1835) );
  AOI22D1BWP30P140LVT U2221 ( .A1(i_data_bus[571]), .A2(n1924), .B1(
        i_data_bus[443]), .B2(n1921), .ZN(n1834) );
  ND4D1BWP30P140LVT U2222 ( .A1(n1837), .A2(n1836), .A3(n1835), .A4(n1834), 
        .ZN(n1848) );
  AOI22D1BWP30P140LVT U2223 ( .A1(i_data_bus[27]), .A2(n2), .B1(i_data_bus[59]), .B2(n1914), .ZN(n1841) );
  AOI22D1BWP30P140LVT U2224 ( .A1(i_data_bus[539]), .A2(n1927), .B1(
        i_data_bus[955]), .B2(n127), .ZN(n1840) );
  AOI22D1BWP30P140LVT U2225 ( .A1(i_data_bus[507]), .A2(n1932), .B1(
        i_data_bus[187]), .B2(n1915), .ZN(n1839) );
  AOI22D1BWP30P140LVT U2226 ( .A1(i_data_bus[315]), .A2(n1922), .B1(
        i_data_bus[251]), .B2(n1911), .ZN(n1838) );
  ND4D1BWP30P140LVT U2227 ( .A1(n1841), .A2(n1840), .A3(n1839), .A4(n1838), 
        .ZN(n1847) );
  AOI22D1BWP30P140LVT U2228 ( .A1(i_data_bus[827]), .A2(n1943), .B1(
        i_data_bus[763]), .B2(n1945), .ZN(n1845) );
  AOI22D1BWP30P140LVT U2229 ( .A1(i_data_bus[731]), .A2(n1942), .B1(
        i_data_bus[699]), .B2(n1947), .ZN(n1844) );
  AOI22D1BWP30P140LVT U2230 ( .A1(i_data_bus[891]), .A2(n1941), .B1(
        i_data_bus[667]), .B2(n1944), .ZN(n1843) );
  AOI22D1BWP30P140LVT U2231 ( .A1(i_data_bus[795]), .A2(n1946), .B1(
        i_data_bus[859]), .B2(n1948), .ZN(n1842) );
  ND4D1BWP30P140LVT U2232 ( .A1(n1845), .A2(n1844), .A3(n1843), .A4(n1842), 
        .ZN(n1846) );
  OR4D1BWP30P140LVT U2233 ( .A1(n1849), .A2(n1848), .A3(n1847), .A4(n1846), 
        .Z(o_data_bus[123]) );
  AOI22D1BWP30P140LVT U2234 ( .A1(i_data_bus[124]), .A2(n1936), .B1(
        i_data_bus[1020]), .B2(n1934), .ZN(n1853) );
  AOI22D1BWP30P140LVT U2235 ( .A1(i_data_bus[636]), .A2(n1910), .B1(
        i_data_bus[444]), .B2(n1921), .ZN(n1852) );
  AOI22D1BWP30P140LVT U2236 ( .A1(i_data_bus[92]), .A2(n1925), .B1(
        i_data_bus[28]), .B2(n2), .ZN(n1851) );
  AOI22D1BWP30P140LVT U2237 ( .A1(i_data_bus[988]), .A2(n1923), .B1(
        i_data_bus[316]), .B2(n1922), .ZN(n1850) );
  ND4D1BWP30P140LVT U2238 ( .A1(n1853), .A2(n1852), .A3(n1851), .A4(n1850), 
        .ZN(n1869) );
  AOI22D1BWP30P140LVT U2239 ( .A1(i_data_bus[572]), .A2(n1924), .B1(
        i_data_bus[380]), .B2(n1926), .ZN(n1857) );
  AOI22D1BWP30P140LVT U2240 ( .A1(i_data_bus[956]), .A2(n127), .B1(
        i_data_bus[412]), .B2(n1279), .ZN(n1856) );
  AOI22D1BWP30P140LVT U2241 ( .A1(i_data_bus[60]), .A2(n1914), .B1(
        i_data_bus[188]), .B2(n1915), .ZN(n1855) );
  AOI22D1BWP30P140LVT U2242 ( .A1(i_data_bus[252]), .A2(n1911), .B1(
        i_data_bus[284]), .B2(n1293), .ZN(n1854) );
  ND4D1BWP30P140LVT U2243 ( .A1(n1857), .A2(n1856), .A3(n1855), .A4(n1854), 
        .ZN(n1868) );
  AOI22D1BWP30P140LVT U2244 ( .A1(i_data_bus[156]), .A2(n1935), .B1(
        i_data_bus[220]), .B2(n1916), .ZN(n1861) );
  AOI22D1BWP30P140LVT U2245 ( .A1(i_data_bus[540]), .A2(n1927), .B1(
        i_data_bus[348]), .B2(n1913), .ZN(n1860) );
  AOI22D1BWP30P140LVT U2246 ( .A1(i_data_bus[924]), .A2(n128), .B1(
        i_data_bus[476]), .B2(n1933), .ZN(n1859) );
  AOI22D1BWP30P140LVT U2247 ( .A1(i_data_bus[604]), .A2(n1912), .B1(
        i_data_bus[508]), .B2(n1932), .ZN(n1858) );
  ND4D1BWP30P140LVT U2248 ( .A1(n1861), .A2(n1860), .A3(n1859), .A4(n1858), 
        .ZN(n1867) );
  AOI22D1BWP30P140LVT U2249 ( .A1(i_data_bus[764]), .A2(n1945), .B1(
        i_data_bus[860]), .B2(n1948), .ZN(n1865) );
  AOI22D1BWP30P140LVT U2250 ( .A1(i_data_bus[796]), .A2(n1946), .B1(
        i_data_bus[828]), .B2(n1943), .ZN(n1864) );
  AOI22D1BWP30P140LVT U2251 ( .A1(i_data_bus[892]), .A2(n1941), .B1(
        i_data_bus[700]), .B2(n1947), .ZN(n1863) );
  AOI22D1BWP30P140LVT U2252 ( .A1(i_data_bus[732]), .A2(n1942), .B1(
        i_data_bus[668]), .B2(n1944), .ZN(n1862) );
  ND4D1BWP30P140LVT U2253 ( .A1(n1865), .A2(n1864), .A3(n1863), .A4(n1862), 
        .ZN(n1866) );
  OR4D1BWP30P140LVT U2254 ( .A1(n1869), .A2(n1868), .A3(n1867), .A4(n1866), 
        .Z(o_data_bus[124]) );
  AOI22D1BWP30P140LVT U2255 ( .A1(i_data_bus[93]), .A2(n1925), .B1(
        i_data_bus[189]), .B2(n1915), .ZN(n1873) );
  AOI22D1BWP30P140LVT U2256 ( .A1(i_data_bus[29]), .A2(n2), .B1(
        i_data_bus[477]), .B2(n1933), .ZN(n1872) );
  AOI22D1BWP30P140LVT U2257 ( .A1(i_data_bus[125]), .A2(n1936), .B1(
        i_data_bus[157]), .B2(n1935), .ZN(n1871) );
  AOI22D1BWP30P140LVT U2258 ( .A1(i_data_bus[637]), .A2(n1910), .B1(
        i_data_bus[221]), .B2(n1916), .ZN(n1870) );
  ND4D1BWP30P140LVT U2259 ( .A1(n1873), .A2(n1872), .A3(n1871), .A4(n1870), 
        .ZN(n1889) );
  AOI22D1BWP30P140LVT U2260 ( .A1(i_data_bus[573]), .A2(n1924), .B1(
        i_data_bus[1021]), .B2(n1934), .ZN(n1877) );
  AOI22D1BWP30P140LVT U2261 ( .A1(i_data_bus[989]), .A2(n1923), .B1(
        i_data_bus[285]), .B2(n1293), .ZN(n1876) );
  AOI22D1BWP30P140LVT U2262 ( .A1(i_data_bus[349]), .A2(n1913), .B1(
        i_data_bus[253]), .B2(n1911), .ZN(n1875) );
  AOI22D1BWP30P140LVT U2263 ( .A1(i_data_bus[605]), .A2(n1912), .B1(
        i_data_bus[317]), .B2(n1922), .ZN(n1874) );
  ND4D1BWP30P140LVT U2264 ( .A1(n1877), .A2(n1876), .A3(n1875), .A4(n1874), 
        .ZN(n1888) );
  AOI22D1BWP30P140LVT U2265 ( .A1(i_data_bus[61]), .A2(n1914), .B1(
        i_data_bus[413]), .B2(n1279), .ZN(n1881) );
  AOI22D1BWP30P140LVT U2266 ( .A1(i_data_bus[445]), .A2(n1921), .B1(
        i_data_bus[509]), .B2(n1932), .ZN(n1880) );
  AOI22D1BWP30P140LVT U2267 ( .A1(i_data_bus[957]), .A2(n127), .B1(
        i_data_bus[541]), .B2(n1927), .ZN(n1879) );
  AOI22D1BWP30P140LVT U2268 ( .A1(i_data_bus[925]), .A2(n128), .B1(
        i_data_bus[381]), .B2(n1926), .ZN(n1878) );
  ND4D1BWP30P140LVT U2269 ( .A1(n1881), .A2(n1880), .A3(n1879), .A4(n1878), 
        .ZN(n1887) );
  AOI22D1BWP30P140LVT U2270 ( .A1(i_data_bus[669]), .A2(n1944), .B1(
        i_data_bus[797]), .B2(n1946), .ZN(n1885) );
  AOI22D1BWP30P140LVT U2271 ( .A1(i_data_bus[829]), .A2(n1943), .B1(
        i_data_bus[861]), .B2(n1948), .ZN(n1884) );
  AOI22D1BWP30P140LVT U2272 ( .A1(i_data_bus[765]), .A2(n1945), .B1(
        i_data_bus[733]), .B2(n1942), .ZN(n1883) );
  AOI22D1BWP30P140LVT U2273 ( .A1(i_data_bus[701]), .A2(n1947), .B1(
        i_data_bus[893]), .B2(n1941), .ZN(n1882) );
  ND4D1BWP30P140LVT U2274 ( .A1(n1885), .A2(n1884), .A3(n1883), .A4(n1882), 
        .ZN(n1886) );
  OR4D1BWP30P140LVT U2275 ( .A1(n1889), .A2(n1888), .A3(n1887), .A4(n1886), 
        .Z(o_data_bus[125]) );
  AOI22D1BWP30P140LVT U2276 ( .A1(i_data_bus[958]), .A2(n127), .B1(
        i_data_bus[606]), .B2(n1912), .ZN(n1893) );
  AOI22D1BWP30P140LVT U2277 ( .A1(i_data_bus[62]), .A2(n1914), .B1(
        i_data_bus[574]), .B2(n1924), .ZN(n1892) );
  AOI22D1BWP30P140LVT U2278 ( .A1(i_data_bus[126]), .A2(n1936), .B1(
        i_data_bus[478]), .B2(n1933), .ZN(n1891) );
  AOI22D1BWP30P140LVT U2279 ( .A1(i_data_bus[638]), .A2(n1910), .B1(
        i_data_bus[446]), .B2(n1921), .ZN(n1890) );
  ND4D1BWP30P140LVT U2280 ( .A1(n1893), .A2(n1892), .A3(n1891), .A4(n1890), 
        .ZN(n1909) );
  AOI22D1BWP30P140LVT U2281 ( .A1(i_data_bus[542]), .A2(n1927), .B1(
        i_data_bus[382]), .B2(n1926), .ZN(n1897) );
  AOI22D1BWP30P140LVT U2282 ( .A1(i_data_bus[222]), .A2(n1916), .B1(
        i_data_bus[510]), .B2(n1932), .ZN(n1896) );
  AOI22D1BWP30P140LVT U2283 ( .A1(i_data_bus[30]), .A2(n2), .B1(
        i_data_bus[158]), .B2(n1935), .ZN(n1895) );
  AOI22D1BWP30P140LVT U2284 ( .A1(i_data_bus[990]), .A2(n1923), .B1(
        i_data_bus[350]), .B2(n1913), .ZN(n1894) );
  ND4D1BWP30P140LVT U2285 ( .A1(n1897), .A2(n1896), .A3(n1895), .A4(n1894), 
        .ZN(n1908) );
  AOI22D1BWP30P140LVT U2286 ( .A1(i_data_bus[318]), .A2(n1922), .B1(
        i_data_bus[190]), .B2(n1915), .ZN(n1901) );
  AOI22D1BWP30P140LVT U2287 ( .A1(i_data_bus[1022]), .A2(n1934), .B1(
        i_data_bus[254]), .B2(n1911), .ZN(n1900) );
  AOI22D1BWP30P140LVT U2288 ( .A1(i_data_bus[94]), .A2(n1925), .B1(
        i_data_bus[286]), .B2(n1293), .ZN(n1899) );
  AOI22D1BWP30P140LVT U2289 ( .A1(i_data_bus[926]), .A2(n128), .B1(
        i_data_bus[414]), .B2(n1279), .ZN(n1898) );
  ND4D1BWP30P140LVT U2290 ( .A1(n1901), .A2(n1900), .A3(n1899), .A4(n1898), 
        .ZN(n1907) );
  AOI22D1BWP30P140LVT U2291 ( .A1(i_data_bus[670]), .A2(n1944), .B1(
        i_data_bus[894]), .B2(n1941), .ZN(n1905) );
  AOI22D1BWP30P140LVT U2292 ( .A1(i_data_bus[798]), .A2(n1946), .B1(
        i_data_bus[830]), .B2(n1943), .ZN(n1904) );
  AOI22D1BWP30P140LVT U2293 ( .A1(i_data_bus[766]), .A2(n1945), .B1(
        i_data_bus[702]), .B2(n1947), .ZN(n1903) );
  AOI22D1BWP30P140LVT U2294 ( .A1(i_data_bus[862]), .A2(n1948), .B1(
        i_data_bus[734]), .B2(n1942), .ZN(n1902) );
  ND4D1BWP30P140LVT U2295 ( .A1(n1905), .A2(n1904), .A3(n1903), .A4(n1902), 
        .ZN(n1906) );
  OR4D1BWP30P140LVT U2296 ( .A1(n1909), .A2(n1908), .A3(n1907), .A4(n1906), 
        .Z(o_data_bus[126]) );
  AOI22D1BWP30P140LVT U2297 ( .A1(i_data_bus[639]), .A2(n1910), .B1(
        i_data_bus[415]), .B2(n1279), .ZN(n1920) );
  AOI22D1BWP30P140LVT U2298 ( .A1(i_data_bus[607]), .A2(n1912), .B1(
        i_data_bus[255]), .B2(n1911), .ZN(n1919) );
  AOI22D1BWP30P140LVT U2299 ( .A1(i_data_bus[63]), .A2(n1914), .B1(
        i_data_bus[351]), .B2(n1913), .ZN(n1918) );
  AOI22D1BWP30P140LVT U2300 ( .A1(i_data_bus[223]), .A2(n1916), .B1(
        i_data_bus[191]), .B2(n1915), .ZN(n1917) );
  ND4D1BWP30P140LVT U2301 ( .A1(n1920), .A2(n1919), .A3(n1918), .A4(n1917), 
        .ZN(n1956) );
  AOI22D1BWP30P140LVT U2302 ( .A1(i_data_bus[319]), .A2(n1922), .B1(
        i_data_bus[447]), .B2(n1921), .ZN(n1931) );
  AOI22D1BWP30P140LVT U2303 ( .A1(i_data_bus[991]), .A2(n1923), .B1(
        i_data_bus[959]), .B2(n127), .ZN(n1930) );
  AOI22D1BWP30P140LVT U2304 ( .A1(i_data_bus[95]), .A2(n1925), .B1(
        i_data_bus[575]), .B2(n1924), .ZN(n1929) );
  AOI22D1BWP30P140LVT U2305 ( .A1(i_data_bus[543]), .A2(n1927), .B1(
        i_data_bus[383]), .B2(n1926), .ZN(n1928) );
  ND4D1BWP30P140LVT U2306 ( .A1(n1931), .A2(n1930), .A3(n1929), .A4(n1928), 
        .ZN(n1955) );
  AOI22D1BWP30P140LVT U2307 ( .A1(i_data_bus[511]), .A2(n1932), .B1(
        i_data_bus[287]), .B2(n1293), .ZN(n1940) );
  AOI22D1BWP30P140LVT U2308 ( .A1(i_data_bus[927]), .A2(n128), .B1(
        i_data_bus[479]), .B2(n1933), .ZN(n1939) );
  AOI22D1BWP30P140LVT U2309 ( .A1(i_data_bus[1023]), .A2(n1934), .B1(
        i_data_bus[31]), .B2(n2), .ZN(n1938) );
  AOI22D1BWP30P140LVT U2310 ( .A1(i_data_bus[127]), .A2(n1936), .B1(
        i_data_bus[159]), .B2(n1935), .ZN(n1937) );
  ND4D1BWP30P140LVT U2311 ( .A1(n1940), .A2(n1939), .A3(n1938), .A4(n1937), 
        .ZN(n1954) );
  AOI22D1BWP30P140LVT U2312 ( .A1(i_data_bus[735]), .A2(n1942), .B1(
        i_data_bus[895]), .B2(n1941), .ZN(n1952) );
  AOI22D1BWP30P140LVT U2313 ( .A1(i_data_bus[671]), .A2(n1944), .B1(
        i_data_bus[831]), .B2(n1943), .ZN(n1951) );
  AOI22D1BWP30P140LVT U2314 ( .A1(i_data_bus[799]), .A2(n1946), .B1(
        i_data_bus[767]), .B2(n1945), .ZN(n1950) );
  AOI22D1BWP30P140LVT U2315 ( .A1(i_data_bus[863]), .A2(n1948), .B1(
        i_data_bus[703]), .B2(n1947), .ZN(n1949) );
  ND4D1BWP30P140LVT U2316 ( .A1(n1952), .A2(n1951), .A3(n1950), .A4(n1949), 
        .ZN(n1953) );
  OR4D1BWP30P140LVT U2317 ( .A1(n1956), .A2(n1955), .A3(n1954), .A4(n1953), 
        .Z(o_data_bus[127]) );
  NR3D0P7BWP30P140LVT U2318 ( .A1(n5490), .A2(n1957), .A3(n1978), .ZN(n2626)
         );
  INVD1BWP30P140LVT U2319 ( .I(i_cmd[36]), .ZN(n1958) );
  AOI22D1BWP30P140LVT U2320 ( .A1(i_data_bus[960]), .A2(n2626), .B1(
        i_data_bus[128]), .B2(n2600), .ZN(n1962) );
  INR3D2BWP30P140LVT U2321 ( .A1(i_cmd[140]), .B1(n5479), .B2(n1975), .ZN(
        n2618) );
  INR3D2BWP30P140LVT U2322 ( .A1(i_cmd[156]), .B1(n5478), .B2(n1975), .ZN(
        n2617) );
  AOI22D1BWP30P140LVT U2323 ( .A1(i_data_bus[544]), .A2(n2618), .B1(
        i_data_bus[608]), .B2(n2617), .ZN(n1961) );
  INR3D2BWP30P140LVT U2324 ( .A1(i_cmd[60]), .B1(n5471), .B2(n1980), .ZN(n2603) );
  INR3D2BWP30P140LVT U2325 ( .A1(i_cmd[76]), .B1(n4095), .B2(n1977), .ZN(n2604) );
  AOI22D1BWP30P140LVT U2326 ( .A1(i_data_bus[224]), .A2(n2603), .B1(
        i_data_bus[288]), .B2(n2604), .ZN(n1960) );
  INR3D2BWP30P140LVT U2327 ( .A1(i_cmd[124]), .B1(n4110), .B2(n1966), .ZN(
        n2629) );
  INR3D2BWP30P140LVT U2328 ( .A1(i_cmd[108]), .B1(n4085), .B2(n1966), .ZN(
        n2615) );
  AOI22D1BWP30P140LVT U2329 ( .A1(i_data_bus[480]), .A2(n2629), .B1(
        i_data_bus[416]), .B2(n2615), .ZN(n1959) );
  ND4D1BWP30P140LVT U2330 ( .A1(n1962), .A2(n1961), .A3(n1960), .A4(n1959), 
        .ZN(n1998) );
  INR3D2BWP30P140LVT U2331 ( .A1(i_cmd[84]), .B1(n4084), .B2(n1977), .ZN(n2625) );
  INVD1BWP30P140LVT U2332 ( .I(i_cmd[68]), .ZN(n1963) );
  NR3D0P7BWP30P140LVT U2333 ( .A1(n5497), .A2(n1963), .A3(n1977), .ZN(n1964)
         );
  AOI22D1BWP30P140LVT U2334 ( .A1(i_data_bus[320]), .A2(n2625), .B1(
        i_data_bus[256]), .B2(n2606), .ZN(n1974) );
  NR3D0P7BWP30P140LVT U2335 ( .A1(n5476), .A2(n140), .A3(n1966), .ZN(n1965) );
  INR3D2BWP30P140LVT U2336 ( .A1(i_cmd[116]), .B1(n4083), .B2(n1966), .ZN(
        n2599) );
  AOI22D1BWP30P140LVT U2337 ( .A1(i_data_bus[384]), .A2(n2614), .B1(
        i_data_bus[448]), .B2(n2599), .ZN(n1973) );
  NR3D0P7BWP30P140LVT U2338 ( .A1(n5470), .A2(n1967), .A3(n1978), .ZN(n2616)
         );
  NR3D0P7BWP30P140LVT U2339 ( .A1(n5486), .A2(n1968), .A3(n1978), .ZN(n2611)
         );
  AOI22D1BWP30P140LVT U2340 ( .A1(i_data_bus[992]), .A2(n2616), .B1(
        i_data_bus[928]), .B2(n2611), .ZN(n1972) );
  INVD1BWP30P140LVT U2341 ( .I(i_cmd[4]), .ZN(n1970) );
  AOI22D1BWP30P140LVT U2342 ( .A1(i_data_bus[0]), .A2(n2624), .B1(
        i_data_bus[64]), .B2(n2602), .ZN(n1971) );
  ND4D1BWP30P140LVT U2343 ( .A1(n1974), .A2(n1973), .A3(n1972), .A4(n1971), 
        .ZN(n1997) );
  INR3D2BWP30P140LVT U2344 ( .A1(i_cmd[52]), .B1(n5494), .B2(n1980), .ZN(n2627) );
  AOI22D1BWP30P140LVT U2345 ( .A1(i_data_bus[512]), .A2(n2601), .B1(
        i_data_bus[192]), .B2(n2627), .ZN(n1984) );
  INR3D2BWP30P140LVT U2346 ( .A1(i_cmd[148]), .B1(n5481), .B2(n1975), .ZN(
        n2630) );
  AOI22D1BWP30P140LVT U2347 ( .A1(i_data_bus[96]), .A2(n2623), .B1(
        i_data_bus[576]), .B2(n2630), .ZN(n1983) );
  INR3D2BWP30P140LVT U2348 ( .A1(i_cmd[92]), .B1(n4074), .B2(n1977), .ZN(n2613) );
  AOI22D1BWP30P140LVT U2349 ( .A1(i_data_bus[32]), .A2(n2628), .B1(
        i_data_bus[352]), .B2(n2613), .ZN(n1982) );
  NR3D0P7BWP30P140LVT U2350 ( .A1(n5473), .A2(n1979), .A3(n1978), .ZN(n2612)
         );
  INR3D2BWP30P140LVT U2351 ( .A1(i_cmd[44]), .B1(n5487), .B2(n1980), .ZN(n2605) );
  AOI22D1BWP30P140LVT U2352 ( .A1(i_data_bus[896]), .A2(n2612), .B1(
        i_data_bus[160]), .B2(n2605), .ZN(n1981) );
  ND4D1BWP30P140LVT U2353 ( .A1(n1984), .A2(n1983), .A3(n1982), .A4(n1981), 
        .ZN(n1996) );
  INR3D2BWP30P140LVT U2354 ( .A1(i_cmd[172]), .B1(n5463), .B2(n1990), .ZN(
        n2637) );
  AOI22D1BWP30P140LVT U2355 ( .A1(i_data_bus[672]), .A2(n2637), .B1(
        i_data_bus[800]), .B2(n2635), .ZN(n1994) );
  INVD1BWP30P140LVT U2356 ( .I(i_cmd[196]), .ZN(n1985) );
  AOI22D1BWP30P140LVT U2357 ( .A1(i_data_bus[768]), .A2(n1986), .B1(
        i_data_bus[864]), .B2(n2639), .ZN(n1993) );
  INR3D2BWP30P140LVT U2358 ( .A1(i_cmd[180]), .B1(n5448), .B2(n1990), .ZN(
        n2640) );
  AOI22D1BWP30P140LVT U2359 ( .A1(i_data_bus[832]), .A2(n2638), .B1(
        i_data_bus[704]), .B2(n2640), .ZN(n1992) );
  INVD1BWP30P140LVT U2360 ( .I(i_cmd[164]), .ZN(n1988) );
  INR3D2BWP30P140LVT U2361 ( .A1(i_cmd[188]), .B1(n5458), .B2(n1990), .ZN(
        n2636) );
  AOI22D1BWP30P140LVT U2362 ( .A1(i_data_bus[640]), .A2(n1989), .B1(
        i_data_bus[736]), .B2(n2636), .ZN(n1991) );
  ND4D1BWP30P140LVT U2363 ( .A1(n1994), .A2(n1993), .A3(n1992), .A4(n1991), 
        .ZN(n1995) );
  OR4D1BWP30P140LVT U2364 ( .A1(n1998), .A2(n1997), .A3(n1996), .A4(n1995), 
        .Z(o_data_bus[128]) );
  AOI22D1BWP30P140LVT U2365 ( .A1(i_data_bus[65]), .A2(n2602), .B1(
        i_data_bus[449]), .B2(n2599), .ZN(n2002) );
  AOI22D1BWP30P140LVT U2366 ( .A1(i_data_bus[33]), .A2(n2628), .B1(
        i_data_bus[161]), .B2(n2605), .ZN(n2001) );
  AOI22D1BWP30P140LVT U2367 ( .A1(i_data_bus[257]), .A2(n2606), .B1(
        i_data_bus[289]), .B2(n2604), .ZN(n2000) );
  AOI22D1BWP30P140LVT U2368 ( .A1(i_data_bus[609]), .A2(n2617), .B1(
        i_data_bus[1]), .B2(n2624), .ZN(n1999) );
  ND4D1BWP30P140LVT U2369 ( .A1(n2002), .A2(n2001), .A3(n2000), .A4(n1999), 
        .ZN(n2018) );
  AOI22D1BWP30P140LVT U2370 ( .A1(i_data_bus[225]), .A2(n2603), .B1(
        i_data_bus[129]), .B2(n2600), .ZN(n2006) );
  AOI22D1BWP30P140LVT U2371 ( .A1(i_data_bus[545]), .A2(n2618), .B1(
        i_data_bus[193]), .B2(n2627), .ZN(n2005) );
  AOI22D1BWP30P140LVT U2372 ( .A1(i_data_bus[577]), .A2(n2630), .B1(
        i_data_bus[321]), .B2(n2625), .ZN(n2004) );
  AOI22D1BWP30P140LVT U2373 ( .A1(i_data_bus[385]), .A2(n2614), .B1(
        i_data_bus[481]), .B2(n2629), .ZN(n2003) );
  ND4D1BWP30P140LVT U2374 ( .A1(n2006), .A2(n2005), .A3(n2004), .A4(n2003), 
        .ZN(n2017) );
  AOI22D1BWP30P140LVT U2375 ( .A1(i_data_bus[97]), .A2(n2623), .B1(
        i_data_bus[993]), .B2(n2616), .ZN(n2010) );
  AOI22D1BWP30P140LVT U2376 ( .A1(i_data_bus[353]), .A2(n2613), .B1(
        i_data_bus[417]), .B2(n2615), .ZN(n2009) );
  AOI22D1BWP30P140LVT U2377 ( .A1(i_data_bus[961]), .A2(n2626), .B1(
        i_data_bus[513]), .B2(n2601), .ZN(n2008) );
  AOI22D1BWP30P140LVT U2378 ( .A1(i_data_bus[897]), .A2(n2612), .B1(
        i_data_bus[929]), .B2(n2611), .ZN(n2007) );
  ND4D1BWP30P140LVT U2379 ( .A1(n2010), .A2(n2009), .A3(n2008), .A4(n2007), 
        .ZN(n2016) );
  AOI22D1BWP30P140LVT U2380 ( .A1(i_data_bus[865]), .A2(n2639), .B1(
        i_data_bus[737]), .B2(n2636), .ZN(n2014) );
  AOI22D1BWP30P140LVT U2381 ( .A1(i_data_bus[641]), .A2(n1989), .B1(
        i_data_bus[801]), .B2(n2635), .ZN(n2013) );
  AOI22D1BWP30P140LVT U2382 ( .A1(i_data_bus[705]), .A2(n2640), .B1(
        i_data_bus[769]), .B2(n1986), .ZN(n2012) );
  AOI22D1BWP30P140LVT U2383 ( .A1(i_data_bus[673]), .A2(n2637), .B1(
        i_data_bus[833]), .B2(n2638), .ZN(n2011) );
  ND4D1BWP30P140LVT U2384 ( .A1(n2014), .A2(n2013), .A3(n2012), .A4(n2011), 
        .ZN(n2015) );
  OR4D1BWP30P140LVT U2385 ( .A1(n2018), .A2(n2017), .A3(n2016), .A4(n2015), 
        .Z(o_data_bus[129]) );
  AOI22D1BWP30P140LVT U2386 ( .A1(i_data_bus[578]), .A2(n2630), .B1(
        i_data_bus[962]), .B2(n2626), .ZN(n2022) );
  AOI22D1BWP30P140LVT U2387 ( .A1(i_data_bus[418]), .A2(n2615), .B1(
        i_data_bus[450]), .B2(n2599), .ZN(n2021) );
  AOI22D1BWP30P140LVT U2388 ( .A1(i_data_bus[66]), .A2(n2602), .B1(
        i_data_bus[930]), .B2(n2611), .ZN(n2020) );
  AOI22D1BWP30P140LVT U2389 ( .A1(i_data_bus[994]), .A2(n2616), .B1(
        i_data_bus[258]), .B2(n2606), .ZN(n2019) );
  ND4D1BWP30P140LVT U2390 ( .A1(n2022), .A2(n2021), .A3(n2020), .A4(n2019), 
        .ZN(n2038) );
  AOI22D1BWP30P140LVT U2391 ( .A1(i_data_bus[290]), .A2(n2604), .B1(
        i_data_bus[354]), .B2(n2613), .ZN(n2026) );
  AOI22D1BWP30P140LVT U2392 ( .A1(i_data_bus[162]), .A2(n2605), .B1(
        i_data_bus[130]), .B2(n2600), .ZN(n2025) );
  AOI22D1BWP30P140LVT U2393 ( .A1(i_data_bus[194]), .A2(n2627), .B1(
        i_data_bus[482]), .B2(n2629), .ZN(n2024) );
  AOI22D1BWP30P140LVT U2394 ( .A1(i_data_bus[546]), .A2(n2618), .B1(
        i_data_bus[386]), .B2(n2614), .ZN(n2023) );
  ND4D1BWP30P140LVT U2395 ( .A1(n2026), .A2(n2025), .A3(n2024), .A4(n2023), 
        .ZN(n2037) );
  AOI22D1BWP30P140LVT U2396 ( .A1(i_data_bus[34]), .A2(n2628), .B1(
        i_data_bus[322]), .B2(n2625), .ZN(n2030) );
  AOI22D1BWP30P140LVT U2397 ( .A1(i_data_bus[2]), .A2(n2624), .B1(
        i_data_bus[514]), .B2(n2601), .ZN(n2029) );
  AOI22D1BWP30P140LVT U2398 ( .A1(i_data_bus[610]), .A2(n2617), .B1(
        i_data_bus[226]), .B2(n2603), .ZN(n2028) );
  AOI22D1BWP30P140LVT U2399 ( .A1(i_data_bus[898]), .A2(n2612), .B1(
        i_data_bus[98]), .B2(n2623), .ZN(n2027) );
  ND4D1BWP30P140LVT U2400 ( .A1(n2030), .A2(n2029), .A3(n2028), .A4(n2027), 
        .ZN(n2036) );
  AOI22D1BWP30P140LVT U2401 ( .A1(i_data_bus[674]), .A2(n2637), .B1(
        i_data_bus[834]), .B2(n2638), .ZN(n2034) );
  AOI22D1BWP30P140LVT U2402 ( .A1(i_data_bus[738]), .A2(n2636), .B1(
        i_data_bus[642]), .B2(n1989), .ZN(n2033) );
  AOI22D1BWP30P140LVT U2403 ( .A1(i_data_bus[866]), .A2(n2639), .B1(
        i_data_bus[706]), .B2(n2640), .ZN(n2032) );
  AOI22D1BWP30P140LVT U2404 ( .A1(i_data_bus[802]), .A2(n2635), .B1(
        i_data_bus[770]), .B2(n1986), .ZN(n2031) );
  ND4D1BWP30P140LVT U2405 ( .A1(n2034), .A2(n2033), .A3(n2032), .A4(n2031), 
        .ZN(n2035) );
  OR4D1BWP30P140LVT U2406 ( .A1(n2038), .A2(n2037), .A3(n2036), .A4(n2035), 
        .Z(o_data_bus[130]) );
  AOI22D1BWP30P140LVT U2407 ( .A1(i_data_bus[67]), .A2(n2602), .B1(
        i_data_bus[515]), .B2(n2601), .ZN(n2042) );
  AOI22D1BWP30P140LVT U2408 ( .A1(i_data_bus[579]), .A2(n2630), .B1(
        i_data_bus[547]), .B2(n2618), .ZN(n2041) );
  AOI22D1BWP30P140LVT U2409 ( .A1(i_data_bus[963]), .A2(n2626), .B1(
        i_data_bus[419]), .B2(n2615), .ZN(n2040) );
  AOI22D1BWP30P140LVT U2410 ( .A1(i_data_bus[899]), .A2(n2612), .B1(
        i_data_bus[35]), .B2(n2628), .ZN(n2039) );
  ND4D1BWP30P140LVT U2411 ( .A1(n2042), .A2(n2041), .A3(n2040), .A4(n2039), 
        .ZN(n2058) );
  AOI22D1BWP30P140LVT U2412 ( .A1(i_data_bus[3]), .A2(n2624), .B1(
        i_data_bus[99]), .B2(n2623), .ZN(n2046) );
  AOI22D1BWP30P140LVT U2413 ( .A1(i_data_bus[931]), .A2(n2611), .B1(
        i_data_bus[355]), .B2(n2613), .ZN(n2045) );
  AOI22D1BWP30P140LVT U2414 ( .A1(i_data_bus[483]), .A2(n2629), .B1(
        i_data_bus[227]), .B2(n2603), .ZN(n2044) );
  AOI22D1BWP30P140LVT U2415 ( .A1(i_data_bus[995]), .A2(n2616), .B1(
        i_data_bus[195]), .B2(n2627), .ZN(n2043) );
  ND4D1BWP30P140LVT U2416 ( .A1(n2046), .A2(n2045), .A3(n2044), .A4(n2043), 
        .ZN(n2057) );
  AOI22D1BWP30P140LVT U2417 ( .A1(i_data_bus[131]), .A2(n2600), .B1(
        i_data_bus[163]), .B2(n2605), .ZN(n2050) );
  AOI22D1BWP30P140LVT U2418 ( .A1(i_data_bus[611]), .A2(n2617), .B1(
        i_data_bus[259]), .B2(n2606), .ZN(n2049) );
  AOI22D1BWP30P140LVT U2419 ( .A1(i_data_bus[387]), .A2(n2614), .B1(
        i_data_bus[291]), .B2(n2604), .ZN(n2048) );
  AOI22D1BWP30P140LVT U2420 ( .A1(i_data_bus[323]), .A2(n2625), .B1(
        i_data_bus[451]), .B2(n2599), .ZN(n2047) );
  ND4D1BWP30P140LVT U2421 ( .A1(n2050), .A2(n2049), .A3(n2048), .A4(n2047), 
        .ZN(n2056) );
  AOI22D1BWP30P140LVT U2422 ( .A1(i_data_bus[835]), .A2(n2638), .B1(
        i_data_bus[867]), .B2(n2639), .ZN(n2054) );
  AOI22D1BWP30P140LVT U2423 ( .A1(i_data_bus[771]), .A2(n1986), .B1(
        i_data_bus[675]), .B2(n2637), .ZN(n2053) );
  AOI22D1BWP30P140LVT U2424 ( .A1(i_data_bus[739]), .A2(n2636), .B1(
        i_data_bus[803]), .B2(n2635), .ZN(n2052) );
  AOI22D1BWP30P140LVT U2425 ( .A1(i_data_bus[643]), .A2(n1989), .B1(
        i_data_bus[707]), .B2(n2640), .ZN(n2051) );
  ND4D1BWP30P140LVT U2426 ( .A1(n2054), .A2(n2053), .A3(n2052), .A4(n2051), 
        .ZN(n2055) );
  OR4D1BWP30P140LVT U2427 ( .A1(n2058), .A2(n2057), .A3(n2056), .A4(n2055), 
        .Z(o_data_bus[131]) );
  AOI22D1BWP30P140LVT U2428 ( .A1(i_data_bus[324]), .A2(n2625), .B1(
        i_data_bus[388]), .B2(n2614), .ZN(n2062) );
  AOI22D1BWP30P140LVT U2429 ( .A1(i_data_bus[516]), .A2(n2601), .B1(
        i_data_bus[36]), .B2(n2628), .ZN(n2061) );
  AOI22D1BWP30P140LVT U2430 ( .A1(i_data_bus[132]), .A2(n2600), .B1(
        i_data_bus[484]), .B2(n2629), .ZN(n2060) );
  AOI22D1BWP30P140LVT U2431 ( .A1(i_data_bus[580]), .A2(n2630), .B1(
        i_data_bus[420]), .B2(n2615), .ZN(n2059) );
  ND4D1BWP30P140LVT U2432 ( .A1(n2062), .A2(n2061), .A3(n2060), .A4(n2059), 
        .ZN(n2078) );
  AOI22D1BWP30P140LVT U2433 ( .A1(i_data_bus[4]), .A2(n2624), .B1(
        i_data_bus[452]), .B2(n2599), .ZN(n2066) );
  AOI22D1BWP30P140LVT U2434 ( .A1(i_data_bus[932]), .A2(n2611), .B1(
        i_data_bus[228]), .B2(n2603), .ZN(n2065) );
  AOI22D1BWP30P140LVT U2435 ( .A1(i_data_bus[100]), .A2(n2623), .B1(
        i_data_bus[164]), .B2(n2605), .ZN(n2064) );
  AOI22D1BWP30P140LVT U2436 ( .A1(i_data_bus[964]), .A2(n2626), .B1(
        i_data_bus[356]), .B2(n2613), .ZN(n2063) );
  ND4D1BWP30P140LVT U2437 ( .A1(n2066), .A2(n2065), .A3(n2064), .A4(n2063), 
        .ZN(n2077) );
  AOI22D1BWP30P140LVT U2438 ( .A1(i_data_bus[68]), .A2(n2602), .B1(
        i_data_bus[292]), .B2(n2604), .ZN(n2070) );
  AOI22D1BWP30P140LVT U2439 ( .A1(i_data_bus[612]), .A2(n2617), .B1(
        i_data_bus[900]), .B2(n2612), .ZN(n2069) );
  AOI22D1BWP30P140LVT U2440 ( .A1(i_data_bus[548]), .A2(n2618), .B1(
        i_data_bus[196]), .B2(n2627), .ZN(n2068) );
  AOI22D1BWP30P140LVT U2441 ( .A1(i_data_bus[996]), .A2(n2616), .B1(
        i_data_bus[260]), .B2(n2606), .ZN(n2067) );
  ND4D1BWP30P140LVT U2442 ( .A1(n2070), .A2(n2069), .A3(n2068), .A4(n2067), 
        .ZN(n2076) );
  AOI22D1BWP30P140LVT U2443 ( .A1(i_data_bus[868]), .A2(n2639), .B1(
        i_data_bus[644]), .B2(n1989), .ZN(n2074) );
  AOI22D1BWP30P140LVT U2444 ( .A1(i_data_bus[772]), .A2(n1986), .B1(
        i_data_bus[836]), .B2(n2638), .ZN(n2073) );
  AOI22D1BWP30P140LVT U2445 ( .A1(i_data_bus[740]), .A2(n2636), .B1(
        i_data_bus[676]), .B2(n2637), .ZN(n2072) );
  AOI22D1BWP30P140LVT U2446 ( .A1(i_data_bus[708]), .A2(n2640), .B1(
        i_data_bus[804]), .B2(n2635), .ZN(n2071) );
  ND4D1BWP30P140LVT U2447 ( .A1(n2074), .A2(n2073), .A3(n2072), .A4(n2071), 
        .ZN(n2075) );
  OR4D1BWP30P140LVT U2448 ( .A1(n2078), .A2(n2077), .A3(n2076), .A4(n2075), 
        .Z(o_data_bus[132]) );
  AOI22D1BWP30P140LVT U2449 ( .A1(i_data_bus[5]), .A2(n2624), .B1(
        i_data_bus[197]), .B2(n2627), .ZN(n2082) );
  AOI22D1BWP30P140LVT U2450 ( .A1(i_data_bus[997]), .A2(n2616), .B1(
        i_data_bus[69]), .B2(n2602), .ZN(n2081) );
  AOI22D1BWP30P140LVT U2451 ( .A1(i_data_bus[357]), .A2(n2613), .B1(
        i_data_bus[293]), .B2(n2604), .ZN(n2080) );
  AOI22D1BWP30P140LVT U2452 ( .A1(i_data_bus[517]), .A2(n2601), .B1(
        i_data_bus[229]), .B2(n2603), .ZN(n2079) );
  ND4D1BWP30P140LVT U2453 ( .A1(n2082), .A2(n2081), .A3(n2080), .A4(n2079), 
        .ZN(n2098) );
  AOI22D1BWP30P140LVT U2454 ( .A1(i_data_bus[581]), .A2(n2630), .B1(
        i_data_bus[389]), .B2(n2614), .ZN(n2086) );
  AOI22D1BWP30P140LVT U2455 ( .A1(i_data_bus[101]), .A2(n2623), .B1(
        i_data_bus[133]), .B2(n2600), .ZN(n2085) );
  AOI22D1BWP30P140LVT U2456 ( .A1(i_data_bus[453]), .A2(n2599), .B1(
        i_data_bus[325]), .B2(n2625), .ZN(n2084) );
  AOI22D1BWP30P140LVT U2457 ( .A1(i_data_bus[965]), .A2(n2626), .B1(
        i_data_bus[485]), .B2(n2629), .ZN(n2083) );
  ND4D1BWP30P140LVT U2458 ( .A1(n2086), .A2(n2085), .A3(n2084), .A4(n2083), 
        .ZN(n2097) );
  AOI22D1BWP30P140LVT U2459 ( .A1(i_data_bus[613]), .A2(n2617), .B1(
        i_data_bus[421]), .B2(n2615), .ZN(n2090) );
  AOI22D1BWP30P140LVT U2460 ( .A1(i_data_bus[165]), .A2(n2605), .B1(
        i_data_bus[261]), .B2(n2606), .ZN(n2089) );
  AOI22D1BWP30P140LVT U2461 ( .A1(i_data_bus[901]), .A2(n2612), .B1(
        i_data_bus[37]), .B2(n2628), .ZN(n2088) );
  AOI22D1BWP30P140LVT U2462 ( .A1(i_data_bus[549]), .A2(n2618), .B1(
        i_data_bus[933]), .B2(n2611), .ZN(n2087) );
  ND4D1BWP30P140LVT U2463 ( .A1(n2090), .A2(n2089), .A3(n2088), .A4(n2087), 
        .ZN(n2096) );
  AOI22D1BWP30P140LVT U2464 ( .A1(i_data_bus[805]), .A2(n2635), .B1(
        i_data_bus[709]), .B2(n2640), .ZN(n2094) );
  AOI22D1BWP30P140LVT U2465 ( .A1(i_data_bus[677]), .A2(n2637), .B1(
        i_data_bus[837]), .B2(n2638), .ZN(n2093) );
  AOI22D1BWP30P140LVT U2466 ( .A1(i_data_bus[645]), .A2(n1989), .B1(
        i_data_bus[869]), .B2(n2639), .ZN(n2092) );
  AOI22D1BWP30P140LVT U2467 ( .A1(i_data_bus[773]), .A2(n1986), .B1(
        i_data_bus[741]), .B2(n2636), .ZN(n2091) );
  ND4D1BWP30P140LVT U2468 ( .A1(n2094), .A2(n2093), .A3(n2092), .A4(n2091), 
        .ZN(n2095) );
  OR4D1BWP30P140LVT U2469 ( .A1(n2098), .A2(n2097), .A3(n2096), .A4(n2095), 
        .Z(o_data_bus[133]) );
  AOI22D1BWP30P140LVT U2470 ( .A1(i_data_bus[902]), .A2(n2612), .B1(
        i_data_bus[166]), .B2(n2605), .ZN(n2102) );
  AOI22D1BWP30P140LVT U2471 ( .A1(i_data_bus[390]), .A2(n2614), .B1(
        i_data_bus[454]), .B2(n2599), .ZN(n2101) );
  AOI22D1BWP30P140LVT U2472 ( .A1(i_data_bus[582]), .A2(n2630), .B1(
        i_data_bus[550]), .B2(n2618), .ZN(n2100) );
  AOI22D1BWP30P140LVT U2473 ( .A1(i_data_bus[422]), .A2(n2615), .B1(
        i_data_bus[294]), .B2(n2604), .ZN(n2099) );
  ND4D1BWP30P140LVT U2474 ( .A1(n2102), .A2(n2101), .A3(n2100), .A4(n2099), 
        .ZN(n2118) );
  AOI22D1BWP30P140LVT U2475 ( .A1(i_data_bus[70]), .A2(n2602), .B1(
        i_data_bus[102]), .B2(n2623), .ZN(n2106) );
  AOI22D1BWP30P140LVT U2476 ( .A1(i_data_bus[358]), .A2(n2613), .B1(
        i_data_bus[198]), .B2(n2627), .ZN(n2105) );
  AOI22D1BWP30P140LVT U2477 ( .A1(i_data_bus[38]), .A2(n2628), .B1(
        i_data_bus[326]), .B2(n2625), .ZN(n2104) );
  AOI22D1BWP30P140LVT U2478 ( .A1(i_data_bus[934]), .A2(n2611), .B1(
        i_data_bus[486]), .B2(n2629), .ZN(n2103) );
  ND4D1BWP30P140LVT U2479 ( .A1(n2106), .A2(n2105), .A3(n2104), .A4(n2103), 
        .ZN(n2117) );
  AOI22D1BWP30P140LVT U2480 ( .A1(i_data_bus[6]), .A2(n2624), .B1(
        i_data_bus[518]), .B2(n2601), .ZN(n2110) );
  AOI22D1BWP30P140LVT U2481 ( .A1(i_data_bus[614]), .A2(n2617), .B1(
        i_data_bus[998]), .B2(n2616), .ZN(n2109) );
  AOI22D1BWP30P140LVT U2482 ( .A1(i_data_bus[966]), .A2(n2626), .B1(
        i_data_bus[262]), .B2(n2606), .ZN(n2108) );
  AOI22D1BWP30P140LVT U2483 ( .A1(i_data_bus[230]), .A2(n2603), .B1(
        i_data_bus[134]), .B2(n2600), .ZN(n2107) );
  ND4D1BWP30P140LVT U2484 ( .A1(n2110), .A2(n2109), .A3(n2108), .A4(n2107), 
        .ZN(n2116) );
  AOI22D1BWP30P140LVT U2485 ( .A1(i_data_bus[646]), .A2(n1989), .B1(
        i_data_bus[678]), .B2(n2637), .ZN(n2114) );
  AOI22D1BWP30P140LVT U2486 ( .A1(i_data_bus[870]), .A2(n2639), .B1(
        i_data_bus[838]), .B2(n2638), .ZN(n2113) );
  AOI22D1BWP30P140LVT U2487 ( .A1(i_data_bus[710]), .A2(n2640), .B1(
        i_data_bus[774]), .B2(n1986), .ZN(n2112) );
  AOI22D1BWP30P140LVT U2488 ( .A1(i_data_bus[806]), .A2(n2635), .B1(
        i_data_bus[742]), .B2(n2636), .ZN(n2111) );
  ND4D1BWP30P140LVT U2489 ( .A1(n2114), .A2(n2113), .A3(n2112), .A4(n2111), 
        .ZN(n2115) );
  OR4D1BWP30P140LVT U2490 ( .A1(n2118), .A2(n2117), .A3(n2116), .A4(n2115), 
        .Z(o_data_bus[134]) );
  AOI22D1BWP30P140LVT U2491 ( .A1(i_data_bus[967]), .A2(n2626), .B1(
        i_data_bus[359]), .B2(n2613), .ZN(n2122) );
  AOI22D1BWP30P140LVT U2492 ( .A1(i_data_bus[615]), .A2(n2617), .B1(
        i_data_bus[519]), .B2(n2601), .ZN(n2121) );
  AOI22D1BWP30P140LVT U2493 ( .A1(i_data_bus[935]), .A2(n2611), .B1(
        i_data_bus[135]), .B2(n2600), .ZN(n2120) );
  AOI22D1BWP30P140LVT U2494 ( .A1(i_data_bus[487]), .A2(n2629), .B1(
        i_data_bus[167]), .B2(n2605), .ZN(n2119) );
  ND4D1BWP30P140LVT U2495 ( .A1(n2122), .A2(n2121), .A3(n2120), .A4(n2119), 
        .ZN(n2138) );
  AOI22D1BWP30P140LVT U2496 ( .A1(i_data_bus[103]), .A2(n2623), .B1(
        i_data_bus[7]), .B2(n2624), .ZN(n2126) );
  AOI22D1BWP30P140LVT U2497 ( .A1(i_data_bus[39]), .A2(n2628), .B1(
        i_data_bus[199]), .B2(n2627), .ZN(n2125) );
  AOI22D1BWP30P140LVT U2498 ( .A1(i_data_bus[263]), .A2(n2606), .B1(
        i_data_bus[295]), .B2(n2604), .ZN(n2124) );
  AOI22D1BWP30P140LVT U2499 ( .A1(i_data_bus[903]), .A2(n2612), .B1(
        i_data_bus[231]), .B2(n2603), .ZN(n2123) );
  ND4D1BWP30P140LVT U2500 ( .A1(n2126), .A2(n2125), .A3(n2124), .A4(n2123), 
        .ZN(n2137) );
  AOI22D1BWP30P140LVT U2501 ( .A1(i_data_bus[999]), .A2(n2616), .B1(
        i_data_bus[71]), .B2(n2602), .ZN(n2130) );
  AOI22D1BWP30P140LVT U2502 ( .A1(i_data_bus[423]), .A2(n2615), .B1(
        i_data_bus[327]), .B2(n2625), .ZN(n2129) );
  AOI22D1BWP30P140LVT U2503 ( .A1(i_data_bus[455]), .A2(n2599), .B1(
        i_data_bus[391]), .B2(n2614), .ZN(n2128) );
  AOI22D1BWP30P140LVT U2504 ( .A1(i_data_bus[551]), .A2(n2618), .B1(
        i_data_bus[583]), .B2(n2630), .ZN(n2127) );
  ND4D1BWP30P140LVT U2505 ( .A1(n2130), .A2(n2129), .A3(n2128), .A4(n2127), 
        .ZN(n2136) );
  AOI22D1BWP30P140LVT U2506 ( .A1(i_data_bus[871]), .A2(n2639), .B1(
        i_data_bus[711]), .B2(n2640), .ZN(n2134) );
  AOI22D1BWP30P140LVT U2507 ( .A1(i_data_bus[839]), .A2(n2638), .B1(
        i_data_bus[647]), .B2(n1989), .ZN(n2133) );
  AOI22D1BWP30P140LVT U2508 ( .A1(i_data_bus[679]), .A2(n2637), .B1(
        i_data_bus[775]), .B2(n1986), .ZN(n2132) );
  AOI22D1BWP30P140LVT U2509 ( .A1(i_data_bus[807]), .A2(n2635), .B1(
        i_data_bus[743]), .B2(n2636), .ZN(n2131) );
  ND4D1BWP30P140LVT U2510 ( .A1(n2134), .A2(n2133), .A3(n2132), .A4(n2131), 
        .ZN(n2135) );
  OR4D1BWP30P140LVT U2511 ( .A1(n2138), .A2(n2137), .A3(n2136), .A4(n2135), 
        .Z(o_data_bus[135]) );
  AOI22D1BWP30P140LVT U2512 ( .A1(i_data_bus[424]), .A2(n2615), .B1(
        i_data_bus[360]), .B2(n2613), .ZN(n2142) );
  AOI22D1BWP30P140LVT U2513 ( .A1(i_data_bus[552]), .A2(n2618), .B1(
        i_data_bus[40]), .B2(n2628), .ZN(n2141) );
  AOI22D1BWP30P140LVT U2514 ( .A1(i_data_bus[104]), .A2(n2623), .B1(
        i_data_bus[1000]), .B2(n2616), .ZN(n2140) );
  AOI22D1BWP30P140LVT U2515 ( .A1(i_data_bus[520]), .A2(n2601), .B1(
        i_data_bus[72]), .B2(n2602), .ZN(n2139) );
  ND4D1BWP30P140LVT U2516 ( .A1(n2142), .A2(n2141), .A3(n2140), .A4(n2139), 
        .ZN(n2158) );
  AOI22D1BWP30P140LVT U2517 ( .A1(i_data_bus[936]), .A2(n2611), .B1(
        i_data_bus[328]), .B2(n2625), .ZN(n2146) );
  AOI22D1BWP30P140LVT U2518 ( .A1(i_data_bus[8]), .A2(n2624), .B1(
        i_data_bus[488]), .B2(n2629), .ZN(n2145) );
  AOI22D1BWP30P140LVT U2519 ( .A1(i_data_bus[968]), .A2(n2626), .B1(
        i_data_bus[296]), .B2(n2604), .ZN(n2144) );
  AOI22D1BWP30P140LVT U2520 ( .A1(i_data_bus[264]), .A2(n2606), .B1(
        i_data_bus[136]), .B2(n2600), .ZN(n2143) );
  ND4D1BWP30P140LVT U2521 ( .A1(n2146), .A2(n2145), .A3(n2144), .A4(n2143), 
        .ZN(n2157) );
  AOI22D1BWP30P140LVT U2522 ( .A1(i_data_bus[456]), .A2(n2599), .B1(
        i_data_bus[200]), .B2(n2627), .ZN(n2150) );
  AOI22D1BWP30P140LVT U2523 ( .A1(i_data_bus[584]), .A2(n2630), .B1(
        i_data_bus[392]), .B2(n2614), .ZN(n2149) );
  AOI22D1BWP30P140LVT U2524 ( .A1(i_data_bus[904]), .A2(n2612), .B1(
        i_data_bus[168]), .B2(n2605), .ZN(n2148) );
  AOI22D1BWP30P140LVT U2525 ( .A1(i_data_bus[616]), .A2(n2617), .B1(
        i_data_bus[232]), .B2(n2603), .ZN(n2147) );
  ND4D1BWP30P140LVT U2526 ( .A1(n2150), .A2(n2149), .A3(n2148), .A4(n2147), 
        .ZN(n2156) );
  AOI22D1BWP30P140LVT U2527 ( .A1(i_data_bus[680]), .A2(n2637), .B1(
        i_data_bus[872]), .B2(n2639), .ZN(n2154) );
  AOI22D1BWP30P140LVT U2528 ( .A1(i_data_bus[840]), .A2(n2638), .B1(
        i_data_bus[776]), .B2(n1986), .ZN(n2153) );
  AOI22D1BWP30P140LVT U2529 ( .A1(i_data_bus[744]), .A2(n2636), .B1(
        i_data_bus[808]), .B2(n2635), .ZN(n2152) );
  AOI22D1BWP30P140LVT U2530 ( .A1(i_data_bus[712]), .A2(n2640), .B1(
        i_data_bus[648]), .B2(n1989), .ZN(n2151) );
  ND4D1BWP30P140LVT U2531 ( .A1(n2154), .A2(n2153), .A3(n2152), .A4(n2151), 
        .ZN(n2155) );
  OR4D1BWP30P140LVT U2532 ( .A1(n2158), .A2(n2157), .A3(n2156), .A4(n2155), 
        .Z(o_data_bus[136]) );
  AOI22D1BWP30P140LVT U2533 ( .A1(i_data_bus[553]), .A2(n2618), .B1(
        i_data_bus[361]), .B2(n2613), .ZN(n2162) );
  AOI22D1BWP30P140LVT U2534 ( .A1(i_data_bus[201]), .A2(n2627), .B1(
        i_data_bus[329]), .B2(n2625), .ZN(n2161) );
  AOI22D1BWP30P140LVT U2535 ( .A1(i_data_bus[233]), .A2(n2603), .B1(
        i_data_bus[137]), .B2(n2600), .ZN(n2160) );
  AOI22D1BWP30P140LVT U2536 ( .A1(i_data_bus[297]), .A2(n2604), .B1(
        i_data_bus[457]), .B2(n2599), .ZN(n2159) );
  ND4D1BWP30P140LVT U2537 ( .A1(n2162), .A2(n2161), .A3(n2160), .A4(n2159), 
        .ZN(n2178) );
  AOI22D1BWP30P140LVT U2538 ( .A1(i_data_bus[9]), .A2(n2624), .B1(
        i_data_bus[585]), .B2(n2630), .ZN(n2166) );
  AOI22D1BWP30P140LVT U2539 ( .A1(i_data_bus[73]), .A2(n2602), .B1(
        i_data_bus[969]), .B2(n2626), .ZN(n2165) );
  AOI22D1BWP30P140LVT U2540 ( .A1(i_data_bus[489]), .A2(n2629), .B1(
        i_data_bus[393]), .B2(n2614), .ZN(n2164) );
  AOI22D1BWP30P140LVT U2541 ( .A1(i_data_bus[105]), .A2(n2623), .B1(
        i_data_bus[1001]), .B2(n2616), .ZN(n2163) );
  ND4D1BWP30P140LVT U2542 ( .A1(n2166), .A2(n2165), .A3(n2164), .A4(n2163), 
        .ZN(n2177) );
  AOI22D1BWP30P140LVT U2543 ( .A1(i_data_bus[41]), .A2(n2628), .B1(
        i_data_bus[265]), .B2(n2606), .ZN(n2170) );
  AOI22D1BWP30P140LVT U2544 ( .A1(i_data_bus[905]), .A2(n2612), .B1(
        i_data_bus[937]), .B2(n2611), .ZN(n2169) );
  AOI22D1BWP30P140LVT U2545 ( .A1(i_data_bus[521]), .A2(n2601), .B1(
        i_data_bus[617]), .B2(n2617), .ZN(n2168) );
  AOI22D1BWP30P140LVT U2546 ( .A1(i_data_bus[169]), .A2(n2605), .B1(
        i_data_bus[425]), .B2(n2615), .ZN(n2167) );
  ND4D1BWP30P140LVT U2547 ( .A1(n2170), .A2(n2169), .A3(n2168), .A4(n2167), 
        .ZN(n2176) );
  AOI22D1BWP30P140LVT U2548 ( .A1(i_data_bus[745]), .A2(n2636), .B1(
        i_data_bus[873]), .B2(n2639), .ZN(n2174) );
  AOI22D1BWP30P140LVT U2549 ( .A1(i_data_bus[681]), .A2(n2637), .B1(
        i_data_bus[649]), .B2(n1989), .ZN(n2173) );
  AOI22D1BWP30P140LVT U2550 ( .A1(i_data_bus[777]), .A2(n1986), .B1(
        i_data_bus[841]), .B2(n2638), .ZN(n2172) );
  AOI22D1BWP30P140LVT U2551 ( .A1(i_data_bus[713]), .A2(n2640), .B1(
        i_data_bus[809]), .B2(n2635), .ZN(n2171) );
  ND4D1BWP30P140LVT U2552 ( .A1(n2174), .A2(n2173), .A3(n2172), .A4(n2171), 
        .ZN(n2175) );
  OR4D1BWP30P140LVT U2553 ( .A1(n2178), .A2(n2177), .A3(n2176), .A4(n2175), 
        .Z(o_data_bus[137]) );
  AOI22D1BWP30P140LVT U2554 ( .A1(i_data_bus[906]), .A2(n2612), .B1(
        i_data_bus[522]), .B2(n2601), .ZN(n2182) );
  AOI22D1BWP30P140LVT U2555 ( .A1(i_data_bus[618]), .A2(n2617), .B1(
        i_data_bus[426]), .B2(n2615), .ZN(n2181) );
  AOI22D1BWP30P140LVT U2556 ( .A1(i_data_bus[970]), .A2(n2626), .B1(
        i_data_bus[266]), .B2(n2606), .ZN(n2180) );
  AOI22D1BWP30P140LVT U2557 ( .A1(i_data_bus[106]), .A2(n2623), .B1(
        i_data_bus[586]), .B2(n2630), .ZN(n2179) );
  ND4D1BWP30P140LVT U2558 ( .A1(n2182), .A2(n2181), .A3(n2180), .A4(n2179), 
        .ZN(n2198) );
  AOI22D1BWP30P140LVT U2559 ( .A1(i_data_bus[74]), .A2(n2602), .B1(
        i_data_bus[394]), .B2(n2614), .ZN(n2186) );
  AOI22D1BWP30P140LVT U2560 ( .A1(i_data_bus[202]), .A2(n2627), .B1(
        i_data_bus[234]), .B2(n2603), .ZN(n2185) );
  AOI22D1BWP30P140LVT U2561 ( .A1(i_data_bus[554]), .A2(n2618), .B1(
        i_data_bus[298]), .B2(n2604), .ZN(n2184) );
  AOI22D1BWP30P140LVT U2562 ( .A1(i_data_bus[42]), .A2(n2628), .B1(
        i_data_bus[362]), .B2(n2613), .ZN(n2183) );
  ND4D1BWP30P140LVT U2563 ( .A1(n2186), .A2(n2185), .A3(n2184), .A4(n2183), 
        .ZN(n2197) );
  AOI22D1BWP30P140LVT U2564 ( .A1(i_data_bus[10]), .A2(n2624), .B1(
        i_data_bus[138]), .B2(n2600), .ZN(n2190) );
  AOI22D1BWP30P140LVT U2565 ( .A1(i_data_bus[1002]), .A2(n2616), .B1(
        i_data_bus[170]), .B2(n2605), .ZN(n2189) );
  AOI22D1BWP30P140LVT U2566 ( .A1(i_data_bus[330]), .A2(n2625), .B1(
        i_data_bus[458]), .B2(n2599), .ZN(n2188) );
  AOI22D1BWP30P140LVT U2567 ( .A1(i_data_bus[938]), .A2(n2611), .B1(
        i_data_bus[490]), .B2(n2629), .ZN(n2187) );
  ND4D1BWP30P140LVT U2568 ( .A1(n2190), .A2(n2189), .A3(n2188), .A4(n2187), 
        .ZN(n2196) );
  AOI22D1BWP30P140LVT U2569 ( .A1(i_data_bus[650]), .A2(n1989), .B1(
        i_data_bus[842]), .B2(n2638), .ZN(n2194) );
  AOI22D1BWP30P140LVT U2570 ( .A1(i_data_bus[778]), .A2(n1986), .B1(
        i_data_bus[874]), .B2(n2639), .ZN(n2193) );
  AOI22D1BWP30P140LVT U2571 ( .A1(i_data_bus[714]), .A2(n2640), .B1(
        i_data_bus[810]), .B2(n2635), .ZN(n2192) );
  AOI22D1BWP30P140LVT U2572 ( .A1(i_data_bus[746]), .A2(n2636), .B1(
        i_data_bus[682]), .B2(n2637), .ZN(n2191) );
  ND4D1BWP30P140LVT U2573 ( .A1(n2194), .A2(n2193), .A3(n2192), .A4(n2191), 
        .ZN(n2195) );
  OR4D1BWP30P140LVT U2574 ( .A1(n2198), .A2(n2197), .A3(n2196), .A4(n2195), 
        .Z(o_data_bus[138]) );
  AOI22D1BWP30P140LVT U2575 ( .A1(i_data_bus[523]), .A2(n2601), .B1(
        i_data_bus[235]), .B2(n2603), .ZN(n2202) );
  AOI22D1BWP30P140LVT U2576 ( .A1(i_data_bus[203]), .A2(n2627), .B1(
        i_data_bus[171]), .B2(n2605), .ZN(n2201) );
  AOI22D1BWP30P140LVT U2577 ( .A1(i_data_bus[971]), .A2(n2626), .B1(
        i_data_bus[587]), .B2(n2630), .ZN(n2200) );
  AOI22D1BWP30P140LVT U2578 ( .A1(i_data_bus[907]), .A2(n2612), .B1(
        i_data_bus[619]), .B2(n2617), .ZN(n2199) );
  ND4D1BWP30P140LVT U2579 ( .A1(n2202), .A2(n2201), .A3(n2200), .A4(n2199), 
        .ZN(n2218) );
  AOI22D1BWP30P140LVT U2580 ( .A1(i_data_bus[107]), .A2(n2623), .B1(
        i_data_bus[427]), .B2(n2615), .ZN(n2206) );
  AOI22D1BWP30P140LVT U2581 ( .A1(i_data_bus[75]), .A2(n2602), .B1(
        i_data_bus[139]), .B2(n2600), .ZN(n2205) );
  AOI22D1BWP30P140LVT U2582 ( .A1(i_data_bus[555]), .A2(n2618), .B1(
        i_data_bus[299]), .B2(n2604), .ZN(n2204) );
  AOI22D1BWP30P140LVT U2583 ( .A1(i_data_bus[939]), .A2(n2611), .B1(
        i_data_bus[267]), .B2(n2606), .ZN(n2203) );
  ND4D1BWP30P140LVT U2584 ( .A1(n2206), .A2(n2205), .A3(n2204), .A4(n2203), 
        .ZN(n2217) );
  AOI22D1BWP30P140LVT U2585 ( .A1(i_data_bus[43]), .A2(n2628), .B1(
        i_data_bus[363]), .B2(n2613), .ZN(n2210) );
  AOI22D1BWP30P140LVT U2586 ( .A1(i_data_bus[11]), .A2(n2624), .B1(
        i_data_bus[459]), .B2(n2599), .ZN(n2209) );
  AOI22D1BWP30P140LVT U2587 ( .A1(i_data_bus[1003]), .A2(n2616), .B1(
        i_data_bus[491]), .B2(n2629), .ZN(n2208) );
  AOI22D1BWP30P140LVT U2588 ( .A1(i_data_bus[395]), .A2(n2614), .B1(
        i_data_bus[331]), .B2(n2625), .ZN(n2207) );
  ND4D1BWP30P140LVT U2589 ( .A1(n2210), .A2(n2209), .A3(n2208), .A4(n2207), 
        .ZN(n2216) );
  AOI22D1BWP30P140LVT U2590 ( .A1(i_data_bus[811]), .A2(n2635), .B1(
        i_data_bus[779]), .B2(n1986), .ZN(n2214) );
  AOI22D1BWP30P140LVT U2591 ( .A1(i_data_bus[843]), .A2(n2638), .B1(
        i_data_bus[683]), .B2(n2637), .ZN(n2213) );
  AOI22D1BWP30P140LVT U2592 ( .A1(i_data_bus[651]), .A2(n1989), .B1(
        i_data_bus[715]), .B2(n2640), .ZN(n2212) );
  AOI22D1BWP30P140LVT U2593 ( .A1(i_data_bus[875]), .A2(n2639), .B1(
        i_data_bus[747]), .B2(n2636), .ZN(n2211) );
  ND4D1BWP30P140LVT U2594 ( .A1(n2214), .A2(n2213), .A3(n2212), .A4(n2211), 
        .ZN(n2215) );
  OR4D1BWP30P140LVT U2595 ( .A1(n2218), .A2(n2217), .A3(n2216), .A4(n2215), 
        .Z(o_data_bus[139]) );
  AOI22D1BWP30P140LVT U2596 ( .A1(i_data_bus[524]), .A2(n2601), .B1(
        i_data_bus[268]), .B2(n2606), .ZN(n2222) );
  AOI22D1BWP30P140LVT U2597 ( .A1(i_data_bus[460]), .A2(n2599), .B1(
        i_data_bus[332]), .B2(n2625), .ZN(n2221) );
  AOI22D1BWP30P140LVT U2598 ( .A1(i_data_bus[620]), .A2(n2617), .B1(
        i_data_bus[972]), .B2(n2626), .ZN(n2220) );
  AOI22D1BWP30P140LVT U2599 ( .A1(i_data_bus[492]), .A2(n2629), .B1(
        i_data_bus[172]), .B2(n2605), .ZN(n2219) );
  ND4D1BWP30P140LVT U2600 ( .A1(n2222), .A2(n2221), .A3(n2220), .A4(n2219), 
        .ZN(n2238) );
  AOI22D1BWP30P140LVT U2601 ( .A1(i_data_bus[76]), .A2(n2602), .B1(
        i_data_bus[204]), .B2(n2627), .ZN(n2226) );
  AOI22D1BWP30P140LVT U2602 ( .A1(i_data_bus[44]), .A2(n2628), .B1(
        i_data_bus[908]), .B2(n2612), .ZN(n2225) );
  AOI22D1BWP30P140LVT U2603 ( .A1(i_data_bus[12]), .A2(n2624), .B1(
        i_data_bus[396]), .B2(n2614), .ZN(n2224) );
  AOI22D1BWP30P140LVT U2604 ( .A1(i_data_bus[108]), .A2(n2623), .B1(
        i_data_bus[140]), .B2(n2600), .ZN(n2223) );
  ND4D1BWP30P140LVT U2605 ( .A1(n2226), .A2(n2225), .A3(n2224), .A4(n2223), 
        .ZN(n2237) );
  AOI22D1BWP30P140LVT U2606 ( .A1(i_data_bus[588]), .A2(n2630), .B1(
        i_data_bus[428]), .B2(n2615), .ZN(n2230) );
  AOI22D1BWP30P140LVT U2607 ( .A1(i_data_bus[556]), .A2(n2618), .B1(
        i_data_bus[364]), .B2(n2613), .ZN(n2229) );
  AOI22D1BWP30P140LVT U2608 ( .A1(i_data_bus[1004]), .A2(n2616), .B1(
        i_data_bus[300]), .B2(n2604), .ZN(n2228) );
  AOI22D1BWP30P140LVT U2609 ( .A1(i_data_bus[940]), .A2(n2611), .B1(
        i_data_bus[236]), .B2(n2603), .ZN(n2227) );
  ND4D1BWP30P140LVT U2610 ( .A1(n2230), .A2(n2229), .A3(n2228), .A4(n2227), 
        .ZN(n2236) );
  AOI22D1BWP30P140LVT U2611 ( .A1(i_data_bus[716]), .A2(n2640), .B1(
        i_data_bus[844]), .B2(n2638), .ZN(n2234) );
  AOI22D1BWP30P140LVT U2612 ( .A1(i_data_bus[780]), .A2(n1986), .B1(
        i_data_bus[748]), .B2(n2636), .ZN(n2233) );
  AOI22D1BWP30P140LVT U2613 ( .A1(i_data_bus[812]), .A2(n2635), .B1(
        i_data_bus[652]), .B2(n1989), .ZN(n2232) );
  AOI22D1BWP30P140LVT U2614 ( .A1(i_data_bus[684]), .A2(n2637), .B1(
        i_data_bus[876]), .B2(n2639), .ZN(n2231) );
  ND4D1BWP30P140LVT U2615 ( .A1(n2234), .A2(n2233), .A3(n2232), .A4(n2231), 
        .ZN(n2235) );
  OR4D1BWP30P140LVT U2616 ( .A1(n2238), .A2(n2237), .A3(n2236), .A4(n2235), 
        .Z(o_data_bus[140]) );
  AOI22D1BWP30P140LVT U2617 ( .A1(i_data_bus[397]), .A2(n2614), .B1(
        i_data_bus[461]), .B2(n2599), .ZN(n2242) );
  AOI22D1BWP30P140LVT U2618 ( .A1(i_data_bus[941]), .A2(n2611), .B1(
        i_data_bus[141]), .B2(n2600), .ZN(n2241) );
  AOI22D1BWP30P140LVT U2619 ( .A1(i_data_bus[525]), .A2(n2601), .B1(
        i_data_bus[557]), .B2(n2618), .ZN(n2240) );
  AOI22D1BWP30P140LVT U2620 ( .A1(i_data_bus[973]), .A2(n2626), .B1(
        i_data_bus[429]), .B2(n2615), .ZN(n2239) );
  ND4D1BWP30P140LVT U2621 ( .A1(n2242), .A2(n2241), .A3(n2240), .A4(n2239), 
        .ZN(n2258) );
  AOI22D1BWP30P140LVT U2622 ( .A1(i_data_bus[493]), .A2(n2629), .B1(
        i_data_bus[333]), .B2(n2625), .ZN(n2246) );
  AOI22D1BWP30P140LVT U2623 ( .A1(i_data_bus[621]), .A2(n2617), .B1(
        i_data_bus[109]), .B2(n2623), .ZN(n2245) );
  AOI22D1BWP30P140LVT U2624 ( .A1(i_data_bus[301]), .A2(n2604), .B1(
        i_data_bus[173]), .B2(n2605), .ZN(n2244) );
  AOI22D1BWP30P140LVT U2625 ( .A1(i_data_bus[589]), .A2(n2630), .B1(
        i_data_bus[269]), .B2(n2606), .ZN(n2243) );
  ND4D1BWP30P140LVT U2626 ( .A1(n2246), .A2(n2245), .A3(n2244), .A4(n2243), 
        .ZN(n2257) );
  AOI22D1BWP30P140LVT U2627 ( .A1(i_data_bus[45]), .A2(n2628), .B1(
        i_data_bus[1005]), .B2(n2616), .ZN(n2250) );
  AOI22D1BWP30P140LVT U2628 ( .A1(i_data_bus[13]), .A2(n2624), .B1(
        i_data_bus[205]), .B2(n2627), .ZN(n2249) );
  AOI22D1BWP30P140LVT U2629 ( .A1(i_data_bus[909]), .A2(n2612), .B1(
        i_data_bus[365]), .B2(n2613), .ZN(n2248) );
  AOI22D1BWP30P140LVT U2630 ( .A1(i_data_bus[77]), .A2(n2602), .B1(
        i_data_bus[237]), .B2(n2603), .ZN(n2247) );
  ND4D1BWP30P140LVT U2631 ( .A1(n2250), .A2(n2249), .A3(n2248), .A4(n2247), 
        .ZN(n2256) );
  AOI22D1BWP30P140LVT U2632 ( .A1(i_data_bus[749]), .A2(n2636), .B1(
        i_data_bus[845]), .B2(n2638), .ZN(n2254) );
  AOI22D1BWP30P140LVT U2633 ( .A1(i_data_bus[813]), .A2(n2635), .B1(
        i_data_bus[717]), .B2(n2640), .ZN(n2253) );
  AOI22D1BWP30P140LVT U2634 ( .A1(i_data_bus[685]), .A2(n2637), .B1(
        i_data_bus[653]), .B2(n1989), .ZN(n2252) );
  AOI22D1BWP30P140LVT U2635 ( .A1(i_data_bus[877]), .A2(n2639), .B1(
        i_data_bus[781]), .B2(n1986), .ZN(n2251) );
  ND4D1BWP30P140LVT U2636 ( .A1(n2254), .A2(n2253), .A3(n2252), .A4(n2251), 
        .ZN(n2255) );
  OR4D1BWP30P140LVT U2637 ( .A1(n2258), .A2(n2257), .A3(n2256), .A4(n2255), 
        .Z(o_data_bus[141]) );
  AOI22D1BWP30P140LVT U2638 ( .A1(i_data_bus[942]), .A2(n2611), .B1(
        i_data_bus[430]), .B2(n2615), .ZN(n2262) );
  AOI22D1BWP30P140LVT U2639 ( .A1(i_data_bus[270]), .A2(n2606), .B1(
        i_data_bus[142]), .B2(n2600), .ZN(n2261) );
  AOI22D1BWP30P140LVT U2640 ( .A1(i_data_bus[334]), .A2(n2625), .B1(
        i_data_bus[398]), .B2(n2614), .ZN(n2260) );
  AOI22D1BWP30P140LVT U2641 ( .A1(i_data_bus[622]), .A2(n2617), .B1(
        i_data_bus[302]), .B2(n2604), .ZN(n2259) );
  ND4D1BWP30P140LVT U2642 ( .A1(n2262), .A2(n2261), .A3(n2260), .A4(n2259), 
        .ZN(n2278) );
  AOI22D1BWP30P140LVT U2643 ( .A1(i_data_bus[558]), .A2(n2618), .B1(
        i_data_bus[174]), .B2(n2605), .ZN(n2266) );
  AOI22D1BWP30P140LVT U2644 ( .A1(i_data_bus[78]), .A2(n2602), .B1(
        i_data_bus[462]), .B2(n2599), .ZN(n2265) );
  AOI22D1BWP30P140LVT U2645 ( .A1(i_data_bus[590]), .A2(n2630), .B1(
        i_data_bus[494]), .B2(n2629), .ZN(n2264) );
  AOI22D1BWP30P140LVT U2646 ( .A1(i_data_bus[366]), .A2(n2613), .B1(
        i_data_bus[238]), .B2(n2603), .ZN(n2263) );
  ND4D1BWP30P140LVT U2647 ( .A1(n2266), .A2(n2265), .A3(n2264), .A4(n2263), 
        .ZN(n2277) );
  AOI22D1BWP30P140LVT U2648 ( .A1(i_data_bus[1006]), .A2(n2616), .B1(
        i_data_bus[526]), .B2(n2601), .ZN(n2270) );
  AOI22D1BWP30P140LVT U2649 ( .A1(i_data_bus[14]), .A2(n2624), .B1(
        i_data_bus[974]), .B2(n2626), .ZN(n2269) );
  AOI22D1BWP30P140LVT U2650 ( .A1(i_data_bus[910]), .A2(n2612), .B1(
        i_data_bus[46]), .B2(n2628), .ZN(n2268) );
  AOI22D1BWP30P140LVT U2651 ( .A1(i_data_bus[110]), .A2(n2623), .B1(
        i_data_bus[206]), .B2(n2627), .ZN(n2267) );
  ND4D1BWP30P140LVT U2652 ( .A1(n2270), .A2(n2269), .A3(n2268), .A4(n2267), 
        .ZN(n2276) );
  AOI22D1BWP30P140LVT U2653 ( .A1(i_data_bus[814]), .A2(n2635), .B1(
        i_data_bus[878]), .B2(n2639), .ZN(n2274) );
  AOI22D1BWP30P140LVT U2654 ( .A1(i_data_bus[750]), .A2(n2636), .B1(
        i_data_bus[718]), .B2(n2640), .ZN(n2273) );
  AOI22D1BWP30P140LVT U2655 ( .A1(i_data_bus[686]), .A2(n2637), .B1(
        i_data_bus[654]), .B2(n1989), .ZN(n2272) );
  AOI22D1BWP30P140LVT U2656 ( .A1(i_data_bus[846]), .A2(n2638), .B1(
        i_data_bus[782]), .B2(n1986), .ZN(n2271) );
  ND4D1BWP30P140LVT U2657 ( .A1(n2274), .A2(n2273), .A3(n2272), .A4(n2271), 
        .ZN(n2275) );
  OR4D1BWP30P140LVT U2658 ( .A1(n2278), .A2(n2277), .A3(n2276), .A4(n2275), 
        .Z(o_data_bus[142]) );
  AOI22D1BWP30P140LVT U2659 ( .A1(i_data_bus[79]), .A2(n2602), .B1(
        i_data_bus[911]), .B2(n2612), .ZN(n2282) );
  AOI22D1BWP30P140LVT U2660 ( .A1(i_data_bus[975]), .A2(n2626), .B1(
        i_data_bus[591]), .B2(n2630), .ZN(n2281) );
  AOI22D1BWP30P140LVT U2661 ( .A1(i_data_bus[559]), .A2(n2618), .B1(
        i_data_bus[495]), .B2(n2629), .ZN(n2280) );
  AOI22D1BWP30P140LVT U2662 ( .A1(i_data_bus[1007]), .A2(n2616), .B1(
        i_data_bus[207]), .B2(n2627), .ZN(n2279) );
  ND4D1BWP30P140LVT U2663 ( .A1(n2282), .A2(n2281), .A3(n2280), .A4(n2279), 
        .ZN(n2298) );
  AOI22D1BWP30P140LVT U2664 ( .A1(i_data_bus[399]), .A2(n2614), .B1(
        i_data_bus[367]), .B2(n2613), .ZN(n2286) );
  AOI22D1BWP30P140LVT U2665 ( .A1(i_data_bus[47]), .A2(n2628), .B1(
        i_data_bus[15]), .B2(n2624), .ZN(n2285) );
  AOI22D1BWP30P140LVT U2666 ( .A1(i_data_bus[111]), .A2(n2623), .B1(
        i_data_bus[143]), .B2(n2600), .ZN(n2284) );
  AOI22D1BWP30P140LVT U2667 ( .A1(i_data_bus[943]), .A2(n2611), .B1(
        i_data_bus[271]), .B2(n2606), .ZN(n2283) );
  ND4D1BWP30P140LVT U2668 ( .A1(n2286), .A2(n2285), .A3(n2284), .A4(n2283), 
        .ZN(n2297) );
  AOI22D1BWP30P140LVT U2669 ( .A1(i_data_bus[623]), .A2(n2617), .B1(
        i_data_bus[463]), .B2(n2599), .ZN(n2290) );
  AOI22D1BWP30P140LVT U2670 ( .A1(i_data_bus[239]), .A2(n2603), .B1(
        i_data_bus[335]), .B2(n2625), .ZN(n2289) );
  AOI22D1BWP30P140LVT U2671 ( .A1(i_data_bus[527]), .A2(n2601), .B1(
        i_data_bus[175]), .B2(n2605), .ZN(n2288) );
  AOI22D1BWP30P140LVT U2672 ( .A1(i_data_bus[431]), .A2(n2615), .B1(
        i_data_bus[303]), .B2(n2604), .ZN(n2287) );
  ND4D1BWP30P140LVT U2673 ( .A1(n2290), .A2(n2289), .A3(n2288), .A4(n2287), 
        .ZN(n2296) );
  AOI22D1BWP30P140LVT U2674 ( .A1(i_data_bus[847]), .A2(n2638), .B1(
        i_data_bus[655]), .B2(n1989), .ZN(n2294) );
  AOI22D1BWP30P140LVT U2675 ( .A1(i_data_bus[719]), .A2(n2640), .B1(
        i_data_bus[879]), .B2(n2639), .ZN(n2293) );
  AOI22D1BWP30P140LVT U2676 ( .A1(i_data_bus[751]), .A2(n2636), .B1(
        i_data_bus[815]), .B2(n2635), .ZN(n2292) );
  AOI22D1BWP30P140LVT U2677 ( .A1(i_data_bus[783]), .A2(n1986), .B1(
        i_data_bus[687]), .B2(n2637), .ZN(n2291) );
  ND4D1BWP30P140LVT U2678 ( .A1(n2294), .A2(n2293), .A3(n2292), .A4(n2291), 
        .ZN(n2295) );
  OR4D1BWP30P140LVT U2679 ( .A1(n2298), .A2(n2297), .A3(n2296), .A4(n2295), 
        .Z(o_data_bus[143]) );
  AOI22D1BWP30P140LVT U2680 ( .A1(i_data_bus[48]), .A2(n2628), .B1(
        i_data_bus[240]), .B2(n2603), .ZN(n2302) );
  AOI22D1BWP30P140LVT U2681 ( .A1(i_data_bus[592]), .A2(n2630), .B1(
        i_data_bus[304]), .B2(n2604), .ZN(n2301) );
  AOI22D1BWP30P140LVT U2682 ( .A1(i_data_bus[528]), .A2(n2601), .B1(
        i_data_bus[112]), .B2(n2623), .ZN(n2300) );
  AOI22D1BWP30P140LVT U2683 ( .A1(i_data_bus[912]), .A2(n2612), .B1(
        i_data_bus[208]), .B2(n2627), .ZN(n2299) );
  ND4D1BWP30P140LVT U2684 ( .A1(n2302), .A2(n2301), .A3(n2300), .A4(n2299), 
        .ZN(n2318) );
  AOI22D1BWP30P140LVT U2685 ( .A1(i_data_bus[80]), .A2(n2602), .B1(
        i_data_bus[624]), .B2(n2617), .ZN(n2306) );
  AOI22D1BWP30P140LVT U2686 ( .A1(i_data_bus[976]), .A2(n2626), .B1(
        i_data_bus[464]), .B2(n2599), .ZN(n2305) );
  AOI22D1BWP30P140LVT U2687 ( .A1(i_data_bus[944]), .A2(n2611), .B1(
        i_data_bus[496]), .B2(n2629), .ZN(n2304) );
  AOI22D1BWP30P140LVT U2688 ( .A1(i_data_bus[1008]), .A2(n2616), .B1(
        i_data_bus[432]), .B2(n2615), .ZN(n2303) );
  ND4D1BWP30P140LVT U2689 ( .A1(n2306), .A2(n2305), .A3(n2304), .A4(n2303), 
        .ZN(n2317) );
  AOI22D1BWP30P140LVT U2690 ( .A1(i_data_bus[560]), .A2(n2618), .B1(
        i_data_bus[272]), .B2(n2606), .ZN(n2310) );
  AOI22D1BWP30P140LVT U2691 ( .A1(i_data_bus[336]), .A2(n2625), .B1(
        i_data_bus[400]), .B2(n2614), .ZN(n2309) );
  AOI22D1BWP30P140LVT U2692 ( .A1(i_data_bus[144]), .A2(n2600), .B1(
        i_data_bus[176]), .B2(n2605), .ZN(n2308) );
  AOI22D1BWP30P140LVT U2693 ( .A1(i_data_bus[16]), .A2(n2624), .B1(
        i_data_bus[368]), .B2(n2613), .ZN(n2307) );
  ND4D1BWP30P140LVT U2694 ( .A1(n2310), .A2(n2309), .A3(n2308), .A4(n2307), 
        .ZN(n2316) );
  AOI22D1BWP30P140LVT U2695 ( .A1(i_data_bus[784]), .A2(n1986), .B1(
        i_data_bus[816]), .B2(n2635), .ZN(n2314) );
  AOI22D1BWP30P140LVT U2696 ( .A1(i_data_bus[720]), .A2(n2640), .B1(
        i_data_bus[848]), .B2(n2638), .ZN(n2313) );
  AOI22D1BWP30P140LVT U2697 ( .A1(i_data_bus[880]), .A2(n2639), .B1(
        i_data_bus[752]), .B2(n2636), .ZN(n2312) );
  AOI22D1BWP30P140LVT U2698 ( .A1(i_data_bus[656]), .A2(n1989), .B1(
        i_data_bus[688]), .B2(n2637), .ZN(n2311) );
  ND4D1BWP30P140LVT U2699 ( .A1(n2314), .A2(n2313), .A3(n2312), .A4(n2311), 
        .ZN(n2315) );
  OR4D1BWP30P140LVT U2700 ( .A1(n2318), .A2(n2317), .A3(n2316), .A4(n2315), 
        .Z(o_data_bus[144]) );
  AOI22D1BWP30P140LVT U2701 ( .A1(i_data_bus[465]), .A2(n2599), .B1(
        i_data_bus[369]), .B2(n2613), .ZN(n2322) );
  AOI22D1BWP30P140LVT U2702 ( .A1(i_data_bus[945]), .A2(n2611), .B1(
        i_data_bus[337]), .B2(n2625), .ZN(n2321) );
  AOI22D1BWP30P140LVT U2703 ( .A1(i_data_bus[241]), .A2(n2603), .B1(
        i_data_bus[273]), .B2(n2606), .ZN(n2320) );
  AOI22D1BWP30P140LVT U2704 ( .A1(i_data_bus[1009]), .A2(n2616), .B1(
        i_data_bus[401]), .B2(n2614), .ZN(n2319) );
  ND4D1BWP30P140LVT U2705 ( .A1(n2322), .A2(n2321), .A3(n2320), .A4(n2319), 
        .ZN(n2338) );
  AOI22D1BWP30P140LVT U2706 ( .A1(i_data_bus[17]), .A2(n2624), .B1(
        i_data_bus[529]), .B2(n2601), .ZN(n2326) );
  AOI22D1BWP30P140LVT U2707 ( .A1(i_data_bus[433]), .A2(n2615), .B1(
        i_data_bus[177]), .B2(n2605), .ZN(n2325) );
  AOI22D1BWP30P140LVT U2708 ( .A1(i_data_bus[593]), .A2(n2630), .B1(
        i_data_bus[305]), .B2(n2604), .ZN(n2324) );
  AOI22D1BWP30P140LVT U2709 ( .A1(i_data_bus[113]), .A2(n2623), .B1(
        i_data_bus[561]), .B2(n2618), .ZN(n2323) );
  ND4D1BWP30P140LVT U2710 ( .A1(n2326), .A2(n2325), .A3(n2324), .A4(n2323), 
        .ZN(n2337) );
  AOI22D1BWP30P140LVT U2711 ( .A1(i_data_bus[145]), .A2(n2600), .B1(
        i_data_bus[497]), .B2(n2629), .ZN(n2330) );
  AOI22D1BWP30P140LVT U2712 ( .A1(i_data_bus[625]), .A2(n2617), .B1(
        i_data_bus[209]), .B2(n2627), .ZN(n2329) );
  AOI22D1BWP30P140LVT U2713 ( .A1(i_data_bus[49]), .A2(n2628), .B1(
        i_data_bus[81]), .B2(n2602), .ZN(n2328) );
  AOI22D1BWP30P140LVT U2714 ( .A1(i_data_bus[913]), .A2(n2612), .B1(
        i_data_bus[977]), .B2(n2626), .ZN(n2327) );
  ND4D1BWP30P140LVT U2715 ( .A1(n2330), .A2(n2329), .A3(n2328), .A4(n2327), 
        .ZN(n2336) );
  AOI22D1BWP30P140LVT U2716 ( .A1(i_data_bus[785]), .A2(n1986), .B1(
        i_data_bus[817]), .B2(n2635), .ZN(n2334) );
  AOI22D1BWP30P140LVT U2717 ( .A1(i_data_bus[881]), .A2(n2639), .B1(
        i_data_bus[753]), .B2(n2636), .ZN(n2333) );
  AOI22D1BWP30P140LVT U2718 ( .A1(i_data_bus[689]), .A2(n2637), .B1(
        i_data_bus[721]), .B2(n2640), .ZN(n2332) );
  AOI22D1BWP30P140LVT U2719 ( .A1(i_data_bus[849]), .A2(n2638), .B1(
        i_data_bus[657]), .B2(n1989), .ZN(n2331) );
  ND4D1BWP30P140LVT U2720 ( .A1(n2334), .A2(n2333), .A3(n2332), .A4(n2331), 
        .ZN(n2335) );
  OR4D1BWP30P140LVT U2721 ( .A1(n2338), .A2(n2337), .A3(n2336), .A4(n2335), 
        .Z(o_data_bus[145]) );
  AOI22D1BWP30P140LVT U2722 ( .A1(i_data_bus[914]), .A2(n2612), .B1(
        i_data_bus[434]), .B2(n2615), .ZN(n2342) );
  AOI22D1BWP30P140LVT U2723 ( .A1(i_data_bus[562]), .A2(n2618), .B1(
        i_data_bus[338]), .B2(n2625), .ZN(n2341) );
  AOI22D1BWP30P140LVT U2724 ( .A1(i_data_bus[978]), .A2(n2626), .B1(
        i_data_bus[306]), .B2(n2604), .ZN(n2340) );
  AOI22D1BWP30P140LVT U2725 ( .A1(i_data_bus[50]), .A2(n2628), .B1(
        i_data_bus[146]), .B2(n2600), .ZN(n2339) );
  ND4D1BWP30P140LVT U2726 ( .A1(n2342), .A2(n2341), .A3(n2340), .A4(n2339), 
        .ZN(n2358) );
  AOI22D1BWP30P140LVT U2727 ( .A1(i_data_bus[18]), .A2(n2624), .B1(
        i_data_bus[178]), .B2(n2605), .ZN(n2346) );
  AOI22D1BWP30P140LVT U2728 ( .A1(i_data_bus[594]), .A2(n2630), .B1(
        i_data_bus[210]), .B2(n2627), .ZN(n2345) );
  AOI22D1BWP30P140LVT U2729 ( .A1(i_data_bus[626]), .A2(n2617), .B1(
        i_data_bus[370]), .B2(n2613), .ZN(n2344) );
  AOI22D1BWP30P140LVT U2730 ( .A1(i_data_bus[1010]), .A2(n2616), .B1(
        i_data_bus[82]), .B2(n2602), .ZN(n2343) );
  ND4D1BWP30P140LVT U2731 ( .A1(n2346), .A2(n2345), .A3(n2344), .A4(n2343), 
        .ZN(n2357) );
  AOI22D1BWP30P140LVT U2732 ( .A1(i_data_bus[114]), .A2(n2623), .B1(
        i_data_bus[402]), .B2(n2614), .ZN(n2350) );
  AOI22D1BWP30P140LVT U2733 ( .A1(i_data_bus[242]), .A2(n2603), .B1(
        i_data_bus[274]), .B2(n2606), .ZN(n2349) );
  AOI22D1BWP30P140LVT U2734 ( .A1(i_data_bus[946]), .A2(n2611), .B1(
        i_data_bus[498]), .B2(n2629), .ZN(n2348) );
  AOI22D1BWP30P140LVT U2735 ( .A1(i_data_bus[530]), .A2(n2601), .B1(
        i_data_bus[466]), .B2(n2599), .ZN(n2347) );
  ND4D1BWP30P140LVT U2736 ( .A1(n2350), .A2(n2349), .A3(n2348), .A4(n2347), 
        .ZN(n2356) );
  AOI22D1BWP30P140LVT U2737 ( .A1(i_data_bus[658]), .A2(n1989), .B1(
        i_data_bus[754]), .B2(n2636), .ZN(n2354) );
  AOI22D1BWP30P140LVT U2738 ( .A1(i_data_bus[882]), .A2(n2639), .B1(
        i_data_bus[850]), .B2(n2638), .ZN(n2353) );
  AOI22D1BWP30P140LVT U2739 ( .A1(i_data_bus[690]), .A2(n2637), .B1(
        i_data_bus[786]), .B2(n1986), .ZN(n2352) );
  AOI22D1BWP30P140LVT U2740 ( .A1(i_data_bus[722]), .A2(n2640), .B1(
        i_data_bus[818]), .B2(n2635), .ZN(n2351) );
  ND4D1BWP30P140LVT U2741 ( .A1(n2354), .A2(n2353), .A3(n2352), .A4(n2351), 
        .ZN(n2355) );
  OR4D1BWP30P140LVT U2742 ( .A1(n2358), .A2(n2357), .A3(n2356), .A4(n2355), 
        .Z(o_data_bus[146]) );
  AOI22D1BWP30P140LVT U2743 ( .A1(i_data_bus[339]), .A2(n2625), .B1(
        i_data_bus[275]), .B2(n2606), .ZN(n2362) );
  AOI22D1BWP30P140LVT U2744 ( .A1(i_data_bus[531]), .A2(n2601), .B1(
        i_data_bus[19]), .B2(n2624), .ZN(n2361) );
  AOI22D1BWP30P140LVT U2745 ( .A1(i_data_bus[947]), .A2(n2611), .B1(
        i_data_bus[499]), .B2(n2629), .ZN(n2360) );
  AOI22D1BWP30P140LVT U2746 ( .A1(i_data_bus[563]), .A2(n2618), .B1(
        i_data_bus[371]), .B2(n2613), .ZN(n2359) );
  ND4D1BWP30P140LVT U2747 ( .A1(n2362), .A2(n2361), .A3(n2360), .A4(n2359), 
        .ZN(n2378) );
  AOI22D1BWP30P140LVT U2748 ( .A1(i_data_bus[979]), .A2(n2626), .B1(
        i_data_bus[627]), .B2(n2617), .ZN(n2366) );
  AOI22D1BWP30P140LVT U2749 ( .A1(i_data_bus[211]), .A2(n2627), .B1(
        i_data_bus[147]), .B2(n2600), .ZN(n2365) );
  AOI22D1BWP30P140LVT U2750 ( .A1(i_data_bus[595]), .A2(n2630), .B1(
        i_data_bus[179]), .B2(n2605), .ZN(n2364) );
  AOI22D1BWP30P140LVT U2751 ( .A1(i_data_bus[51]), .A2(n2628), .B1(
        i_data_bus[243]), .B2(n2603), .ZN(n2363) );
  ND4D1BWP30P140LVT U2752 ( .A1(n2366), .A2(n2365), .A3(n2364), .A4(n2363), 
        .ZN(n2377) );
  AOI22D1BWP30P140LVT U2753 ( .A1(i_data_bus[915]), .A2(n2612), .B1(
        i_data_bus[403]), .B2(n2614), .ZN(n2370) );
  AOI22D1BWP30P140LVT U2754 ( .A1(i_data_bus[83]), .A2(n2602), .B1(
        i_data_bus[435]), .B2(n2615), .ZN(n2369) );
  AOI22D1BWP30P140LVT U2755 ( .A1(i_data_bus[1011]), .A2(n2616), .B1(
        i_data_bus[307]), .B2(n2604), .ZN(n2368) );
  AOI22D1BWP30P140LVT U2756 ( .A1(i_data_bus[115]), .A2(n2623), .B1(
        i_data_bus[467]), .B2(n2599), .ZN(n2367) );
  ND4D1BWP30P140LVT U2757 ( .A1(n2370), .A2(n2369), .A3(n2368), .A4(n2367), 
        .ZN(n2376) );
  AOI22D1BWP30P140LVT U2758 ( .A1(i_data_bus[755]), .A2(n2636), .B1(
        i_data_bus[691]), .B2(n2637), .ZN(n2374) );
  AOI22D1BWP30P140LVT U2759 ( .A1(i_data_bus[787]), .A2(n1986), .B1(
        i_data_bus[851]), .B2(n2638), .ZN(n2373) );
  AOI22D1BWP30P140LVT U2760 ( .A1(i_data_bus[819]), .A2(n2635), .B1(
        i_data_bus[723]), .B2(n2640), .ZN(n2372) );
  AOI22D1BWP30P140LVT U2761 ( .A1(i_data_bus[659]), .A2(n1989), .B1(
        i_data_bus[883]), .B2(n2639), .ZN(n2371) );
  ND4D1BWP30P140LVT U2762 ( .A1(n2374), .A2(n2373), .A3(n2372), .A4(n2371), 
        .ZN(n2375) );
  OR4D1BWP30P140LVT U2763 ( .A1(n2378), .A2(n2377), .A3(n2376), .A4(n2375), 
        .Z(o_data_bus[147]) );
  AOI22D1BWP30P140LVT U2764 ( .A1(i_data_bus[980]), .A2(n2626), .B1(
        i_data_bus[1012]), .B2(n2616), .ZN(n2382) );
  AOI22D1BWP30P140LVT U2765 ( .A1(i_data_bus[244]), .A2(n2603), .B1(
        i_data_bus[180]), .B2(n2605), .ZN(n2381) );
  AOI22D1BWP30P140LVT U2766 ( .A1(i_data_bus[20]), .A2(n2624), .B1(
        i_data_bus[372]), .B2(n2613), .ZN(n2380) );
  AOI22D1BWP30P140LVT U2767 ( .A1(i_data_bus[628]), .A2(n2617), .B1(
        i_data_bus[404]), .B2(n2614), .ZN(n2379) );
  ND4D1BWP30P140LVT U2768 ( .A1(n2382), .A2(n2381), .A3(n2380), .A4(n2379), 
        .ZN(n2398) );
  AOI22D1BWP30P140LVT U2769 ( .A1(i_data_bus[52]), .A2(n2628), .B1(
        i_data_bus[500]), .B2(n2629), .ZN(n2386) );
  AOI22D1BWP30P140LVT U2770 ( .A1(i_data_bus[340]), .A2(n2625), .B1(
        i_data_bus[276]), .B2(n2606), .ZN(n2385) );
  AOI22D1BWP30P140LVT U2771 ( .A1(i_data_bus[948]), .A2(n2611), .B1(
        i_data_bus[148]), .B2(n2600), .ZN(n2384) );
  AOI22D1BWP30P140LVT U2772 ( .A1(i_data_bus[596]), .A2(n2630), .B1(
        i_data_bus[436]), .B2(n2615), .ZN(n2383) );
  ND4D1BWP30P140LVT U2773 ( .A1(n2386), .A2(n2385), .A3(n2384), .A4(n2383), 
        .ZN(n2397) );
  AOI22D1BWP30P140LVT U2774 ( .A1(i_data_bus[532]), .A2(n2601), .B1(
        i_data_bus[308]), .B2(n2604), .ZN(n2390) );
  AOI22D1BWP30P140LVT U2775 ( .A1(i_data_bus[564]), .A2(n2618), .B1(
        i_data_bus[212]), .B2(n2627), .ZN(n2389) );
  AOI22D1BWP30P140LVT U2776 ( .A1(i_data_bus[84]), .A2(n2602), .B1(
        i_data_bus[116]), .B2(n2623), .ZN(n2388) );
  AOI22D1BWP30P140LVT U2777 ( .A1(i_data_bus[916]), .A2(n2612), .B1(
        i_data_bus[468]), .B2(n2599), .ZN(n2387) );
  ND4D1BWP30P140LVT U2778 ( .A1(n2390), .A2(n2389), .A3(n2388), .A4(n2387), 
        .ZN(n2396) );
  AOI22D1BWP30P140LVT U2779 ( .A1(i_data_bus[884]), .A2(n2639), .B1(
        i_data_bus[692]), .B2(n2637), .ZN(n2394) );
  AOI22D1BWP30P140LVT U2780 ( .A1(i_data_bus[724]), .A2(n2640), .B1(
        i_data_bus[820]), .B2(n2635), .ZN(n2393) );
  AOI22D1BWP30P140LVT U2781 ( .A1(i_data_bus[852]), .A2(n2638), .B1(
        i_data_bus[660]), .B2(n1989), .ZN(n2392) );
  AOI22D1BWP30P140LVT U2782 ( .A1(i_data_bus[788]), .A2(n1986), .B1(
        i_data_bus[756]), .B2(n2636), .ZN(n2391) );
  ND4D1BWP30P140LVT U2783 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), 
        .ZN(n2395) );
  OR4D1BWP30P140LVT U2784 ( .A1(n2398), .A2(n2397), .A3(n2396), .A4(n2395), 
        .Z(o_data_bus[148]) );
  AOI22D1BWP30P140LVT U2785 ( .A1(i_data_bus[917]), .A2(n2612), .B1(
        i_data_bus[565]), .B2(n2618), .ZN(n2402) );
  AOI22D1BWP30P140LVT U2786 ( .A1(i_data_bus[1013]), .A2(n2616), .B1(
        i_data_bus[149]), .B2(n2600), .ZN(n2401) );
  AOI22D1BWP30P140LVT U2787 ( .A1(i_data_bus[117]), .A2(n2623), .B1(
        i_data_bus[629]), .B2(n2617), .ZN(n2400) );
  AOI22D1BWP30P140LVT U2788 ( .A1(i_data_bus[277]), .A2(n2606), .B1(
        i_data_bus[373]), .B2(n2613), .ZN(n2399) );
  ND4D1BWP30P140LVT U2789 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), 
        .ZN(n2418) );
  AOI22D1BWP30P140LVT U2790 ( .A1(i_data_bus[53]), .A2(n2628), .B1(
        i_data_bus[533]), .B2(n2601), .ZN(n2406) );
  AOI22D1BWP30P140LVT U2791 ( .A1(i_data_bus[437]), .A2(n2615), .B1(
        i_data_bus[501]), .B2(n2629), .ZN(n2405) );
  AOI22D1BWP30P140LVT U2792 ( .A1(i_data_bus[341]), .A2(n2625), .B1(
        i_data_bus[309]), .B2(n2604), .ZN(n2404) );
  AOI22D1BWP30P140LVT U2793 ( .A1(i_data_bus[597]), .A2(n2630), .B1(
        i_data_bus[181]), .B2(n2605), .ZN(n2403) );
  ND4D1BWP30P140LVT U2794 ( .A1(n2406), .A2(n2405), .A3(n2404), .A4(n2403), 
        .ZN(n2417) );
  AOI22D1BWP30P140LVT U2795 ( .A1(i_data_bus[85]), .A2(n2602), .B1(
        i_data_bus[245]), .B2(n2603), .ZN(n2410) );
  AOI22D1BWP30P140LVT U2796 ( .A1(i_data_bus[21]), .A2(n2624), .B1(
        i_data_bus[469]), .B2(n2599), .ZN(n2409) );
  AOI22D1BWP30P140LVT U2797 ( .A1(i_data_bus[981]), .A2(n2626), .B1(
        i_data_bus[213]), .B2(n2627), .ZN(n2408) );
  AOI22D1BWP30P140LVT U2798 ( .A1(i_data_bus[949]), .A2(n2611), .B1(
        i_data_bus[405]), .B2(n2614), .ZN(n2407) );
  ND4D1BWP30P140LVT U2799 ( .A1(n2410), .A2(n2409), .A3(n2408), .A4(n2407), 
        .ZN(n2416) );
  AOI22D1BWP30P140LVT U2800 ( .A1(i_data_bus[853]), .A2(n2638), .B1(
        i_data_bus[693]), .B2(n2637), .ZN(n2414) );
  AOI22D1BWP30P140LVT U2801 ( .A1(i_data_bus[661]), .A2(n1989), .B1(
        i_data_bus[725]), .B2(n2640), .ZN(n2413) );
  AOI22D1BWP30P140LVT U2802 ( .A1(i_data_bus[821]), .A2(n2635), .B1(
        i_data_bus[885]), .B2(n2639), .ZN(n2412) );
  AOI22D1BWP30P140LVT U2803 ( .A1(i_data_bus[757]), .A2(n2636), .B1(
        i_data_bus[789]), .B2(n1986), .ZN(n2411) );
  ND4D1BWP30P140LVT U2804 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), 
        .ZN(n2415) );
  OR4D1BWP30P140LVT U2805 ( .A1(n2418), .A2(n2417), .A3(n2416), .A4(n2415), 
        .Z(o_data_bus[149]) );
  AOI22D1BWP30P140LVT U2806 ( .A1(i_data_bus[118]), .A2(n2623), .B1(
        i_data_bus[470]), .B2(n2599), .ZN(n2422) );
  AOI22D1BWP30P140LVT U2807 ( .A1(i_data_bus[1014]), .A2(n2616), .B1(
        i_data_bus[982]), .B2(n2626), .ZN(n2421) );
  AOI22D1BWP30P140LVT U2808 ( .A1(i_data_bus[534]), .A2(n2601), .B1(
        i_data_bus[150]), .B2(n2600), .ZN(n2420) );
  AOI22D1BWP30P140LVT U2809 ( .A1(i_data_bus[22]), .A2(n2624), .B1(
        i_data_bus[214]), .B2(n2627), .ZN(n2419) );
  ND4D1BWP30P140LVT U2810 ( .A1(n2422), .A2(n2421), .A3(n2420), .A4(n2419), 
        .ZN(n2438) );
  AOI22D1BWP30P140LVT U2811 ( .A1(i_data_bus[54]), .A2(n2628), .B1(
        i_data_bus[502]), .B2(n2629), .ZN(n2426) );
  AOI22D1BWP30P140LVT U2812 ( .A1(i_data_bus[566]), .A2(n2618), .B1(
        i_data_bus[310]), .B2(n2604), .ZN(n2425) );
  AOI22D1BWP30P140LVT U2813 ( .A1(i_data_bus[598]), .A2(n2630), .B1(
        i_data_bus[246]), .B2(n2603), .ZN(n2424) );
  AOI22D1BWP30P140LVT U2814 ( .A1(i_data_bus[438]), .A2(n2615), .B1(
        i_data_bus[278]), .B2(n2606), .ZN(n2423) );
  ND4D1BWP30P140LVT U2815 ( .A1(n2426), .A2(n2425), .A3(n2424), .A4(n2423), 
        .ZN(n2437) );
  AOI22D1BWP30P140LVT U2816 ( .A1(i_data_bus[86]), .A2(n2602), .B1(
        i_data_bus[630]), .B2(n2617), .ZN(n2430) );
  AOI22D1BWP30P140LVT U2817 ( .A1(i_data_bus[918]), .A2(n2612), .B1(
        i_data_bus[182]), .B2(n2605), .ZN(n2429) );
  AOI22D1BWP30P140LVT U2818 ( .A1(i_data_bus[406]), .A2(n2614), .B1(
        i_data_bus[342]), .B2(n2625), .ZN(n2428) );
  AOI22D1BWP30P140LVT U2819 ( .A1(i_data_bus[950]), .A2(n2611), .B1(
        i_data_bus[374]), .B2(n2613), .ZN(n2427) );
  ND4D1BWP30P140LVT U2820 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), 
        .ZN(n2436) );
  AOI22D1BWP30P140LVT U2821 ( .A1(i_data_bus[694]), .A2(n2637), .B1(
        i_data_bus[758]), .B2(n2636), .ZN(n2434) );
  AOI22D1BWP30P140LVT U2822 ( .A1(i_data_bus[822]), .A2(n2635), .B1(
        i_data_bus[886]), .B2(n2639), .ZN(n2433) );
  AOI22D1BWP30P140LVT U2823 ( .A1(i_data_bus[790]), .A2(n1986), .B1(
        i_data_bus[854]), .B2(n2638), .ZN(n2432) );
  AOI22D1BWP30P140LVT U2824 ( .A1(i_data_bus[726]), .A2(n2640), .B1(
        i_data_bus[662]), .B2(n1989), .ZN(n2431) );
  ND4D1BWP30P140LVT U2825 ( .A1(n2434), .A2(n2433), .A3(n2432), .A4(n2431), 
        .ZN(n2435) );
  OR4D1BWP30P140LVT U2826 ( .A1(n2438), .A2(n2437), .A3(n2436), .A4(n2435), 
        .Z(o_data_bus[150]) );
  AOI22D1BWP30P140LVT U2827 ( .A1(i_data_bus[567]), .A2(n2618), .B1(
        i_data_bus[151]), .B2(n2600), .ZN(n2442) );
  AOI22D1BWP30P140LVT U2828 ( .A1(i_data_bus[919]), .A2(n2612), .B1(
        i_data_bus[503]), .B2(n2629), .ZN(n2441) );
  AOI22D1BWP30P140LVT U2829 ( .A1(i_data_bus[87]), .A2(n2602), .B1(
        i_data_bus[535]), .B2(n2601), .ZN(n2440) );
  AOI22D1BWP30P140LVT U2830 ( .A1(i_data_bus[599]), .A2(n2630), .B1(
        i_data_bus[407]), .B2(n2614), .ZN(n2439) );
  ND4D1BWP30P140LVT U2831 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2439), 
        .ZN(n2458) );
  AOI22D1BWP30P140LVT U2832 ( .A1(i_data_bus[279]), .A2(n2606), .B1(
        i_data_bus[215]), .B2(n2627), .ZN(n2446) );
  AOI22D1BWP30P140LVT U2833 ( .A1(i_data_bus[951]), .A2(n2611), .B1(
        i_data_bus[183]), .B2(n2605), .ZN(n2445) );
  AOI22D1BWP30P140LVT U2834 ( .A1(i_data_bus[471]), .A2(n2599), .B1(
        i_data_bus[375]), .B2(n2613), .ZN(n2444) );
  AOI22D1BWP30P140LVT U2835 ( .A1(i_data_bus[119]), .A2(n2623), .B1(
        i_data_bus[343]), .B2(n2625), .ZN(n2443) );
  ND4D1BWP30P140LVT U2836 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), 
        .ZN(n2457) );
  AOI22D1BWP30P140LVT U2837 ( .A1(i_data_bus[247]), .A2(n2603), .B1(
        i_data_bus[439]), .B2(n2615), .ZN(n2450) );
  AOI22D1BWP30P140LVT U2838 ( .A1(i_data_bus[1015]), .A2(n2616), .B1(
        i_data_bus[311]), .B2(n2604), .ZN(n2449) );
  AOI22D1BWP30P140LVT U2839 ( .A1(i_data_bus[23]), .A2(n2624), .B1(
        i_data_bus[55]), .B2(n2628), .ZN(n2448) );
  AOI22D1BWP30P140LVT U2840 ( .A1(i_data_bus[631]), .A2(n2617), .B1(
        i_data_bus[983]), .B2(n2626), .ZN(n2447) );
  ND4D1BWP30P140LVT U2841 ( .A1(n2450), .A2(n2449), .A3(n2448), .A4(n2447), 
        .ZN(n2456) );
  AOI22D1BWP30P140LVT U2842 ( .A1(i_data_bus[887]), .A2(n2639), .B1(
        i_data_bus[855]), .B2(n2638), .ZN(n2454) );
  AOI22D1BWP30P140LVT U2843 ( .A1(i_data_bus[695]), .A2(n2637), .B1(
        i_data_bus[663]), .B2(n1989), .ZN(n2453) );
  AOI22D1BWP30P140LVT U2844 ( .A1(i_data_bus[759]), .A2(n2636), .B1(
        i_data_bus[823]), .B2(n2635), .ZN(n2452) );
  AOI22D1BWP30P140LVT U2845 ( .A1(i_data_bus[727]), .A2(n2640), .B1(
        i_data_bus[791]), .B2(n1986), .ZN(n2451) );
  ND4D1BWP30P140LVT U2846 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), 
        .ZN(n2455) );
  OR4D1BWP30P140LVT U2847 ( .A1(n2458), .A2(n2457), .A3(n2456), .A4(n2455), 
        .Z(o_data_bus[151]) );
  AOI22D1BWP30P140LVT U2848 ( .A1(i_data_bus[24]), .A2(n2624), .B1(
        i_data_bus[344]), .B2(n2625), .ZN(n2462) );
  AOI22D1BWP30P140LVT U2849 ( .A1(i_data_bus[88]), .A2(n2602), .B1(
        i_data_bus[248]), .B2(n2603), .ZN(n2461) );
  AOI22D1BWP30P140LVT U2850 ( .A1(i_data_bus[920]), .A2(n2612), .B1(
        i_data_bus[472]), .B2(n2599), .ZN(n2460) );
  AOI22D1BWP30P140LVT U2851 ( .A1(i_data_bus[280]), .A2(n2606), .B1(
        i_data_bus[504]), .B2(n2629), .ZN(n2459) );
  ND4D1BWP30P140LVT U2852 ( .A1(n2462), .A2(n2461), .A3(n2460), .A4(n2459), 
        .ZN(n2478) );
  AOI22D1BWP30P140LVT U2853 ( .A1(i_data_bus[984]), .A2(n2626), .B1(
        i_data_bus[184]), .B2(n2605), .ZN(n2466) );
  AOI22D1BWP30P140LVT U2854 ( .A1(i_data_bus[536]), .A2(n2601), .B1(
        i_data_bus[440]), .B2(n2615), .ZN(n2465) );
  AOI22D1BWP30P140LVT U2855 ( .A1(i_data_bus[568]), .A2(n2618), .B1(
        i_data_bus[376]), .B2(n2613), .ZN(n2464) );
  AOI22D1BWP30P140LVT U2856 ( .A1(i_data_bus[632]), .A2(n2617), .B1(
        i_data_bus[600]), .B2(n2630), .ZN(n2463) );
  ND4D1BWP30P140LVT U2857 ( .A1(n2466), .A2(n2465), .A3(n2464), .A4(n2463), 
        .ZN(n2477) );
  AOI22D1BWP30P140LVT U2858 ( .A1(i_data_bus[952]), .A2(n2611), .B1(
        i_data_bus[56]), .B2(n2628), .ZN(n2470) );
  AOI22D1BWP30P140LVT U2859 ( .A1(i_data_bus[120]), .A2(n2623), .B1(
        i_data_bus[152]), .B2(n2600), .ZN(n2469) );
  AOI22D1BWP30P140LVT U2860 ( .A1(i_data_bus[408]), .A2(n2614), .B1(
        i_data_bus[216]), .B2(n2627), .ZN(n2468) );
  AOI22D1BWP30P140LVT U2861 ( .A1(i_data_bus[1016]), .A2(n2616), .B1(
        i_data_bus[312]), .B2(n2604), .ZN(n2467) );
  ND4D1BWP30P140LVT U2862 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), 
        .ZN(n2476) );
  AOI22D1BWP30P140LVT U2863 ( .A1(i_data_bus[792]), .A2(n1986), .B1(
        i_data_bus[728]), .B2(n2640), .ZN(n2474) );
  AOI22D1BWP30P140LVT U2864 ( .A1(i_data_bus[856]), .A2(n2638), .B1(
        i_data_bus[888]), .B2(n2639), .ZN(n2473) );
  AOI22D1BWP30P140LVT U2865 ( .A1(i_data_bus[696]), .A2(n2637), .B1(
        i_data_bus[760]), .B2(n2636), .ZN(n2472) );
  AOI22D1BWP30P140LVT U2866 ( .A1(i_data_bus[824]), .A2(n2635), .B1(
        i_data_bus[664]), .B2(n1989), .ZN(n2471) );
  ND4D1BWP30P140LVT U2867 ( .A1(n2474), .A2(n2473), .A3(n2472), .A4(n2471), 
        .ZN(n2475) );
  OR4D1BWP30P140LVT U2868 ( .A1(n2478), .A2(n2477), .A3(n2476), .A4(n2475), 
        .Z(o_data_bus[152]) );
  AOI22D1BWP30P140LVT U2869 ( .A1(i_data_bus[985]), .A2(n2626), .B1(
        i_data_bus[409]), .B2(n2614), .ZN(n2482) );
  AOI22D1BWP30P140LVT U2870 ( .A1(i_data_bus[377]), .A2(n2613), .B1(
        i_data_bus[441]), .B2(n2615), .ZN(n2481) );
  AOI22D1BWP30P140LVT U2871 ( .A1(i_data_bus[281]), .A2(n2606), .B1(
        i_data_bus[217]), .B2(n2627), .ZN(n2480) );
  AOI22D1BWP30P140LVT U2872 ( .A1(i_data_bus[1017]), .A2(n2616), .B1(
        i_data_bus[89]), .B2(n2602), .ZN(n2479) );
  ND4D1BWP30P140LVT U2873 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), 
        .ZN(n2498) );
  AOI22D1BWP30P140LVT U2874 ( .A1(i_data_bus[601]), .A2(n2630), .B1(
        i_data_bus[313]), .B2(n2604), .ZN(n2486) );
  AOI22D1BWP30P140LVT U2875 ( .A1(i_data_bus[185]), .A2(n2605), .B1(
        i_data_bus[505]), .B2(n2629), .ZN(n2485) );
  AOI22D1BWP30P140LVT U2876 ( .A1(i_data_bus[57]), .A2(n2628), .B1(
        i_data_bus[121]), .B2(n2623), .ZN(n2484) );
  AOI22D1BWP30P140LVT U2877 ( .A1(i_data_bus[537]), .A2(n2601), .B1(
        i_data_bus[473]), .B2(n2599), .ZN(n2483) );
  ND4D1BWP30P140LVT U2878 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), 
        .ZN(n2497) );
  AOI22D1BWP30P140LVT U2879 ( .A1(i_data_bus[25]), .A2(n2624), .B1(
        i_data_bus[249]), .B2(n2603), .ZN(n2490) );
  AOI22D1BWP30P140LVT U2880 ( .A1(i_data_bus[569]), .A2(n2618), .B1(
        i_data_bus[153]), .B2(n2600), .ZN(n2489) );
  AOI22D1BWP30P140LVT U2881 ( .A1(i_data_bus[633]), .A2(n2617), .B1(
        i_data_bus[953]), .B2(n2611), .ZN(n2488) );
  AOI22D1BWP30P140LVT U2882 ( .A1(i_data_bus[921]), .A2(n2612), .B1(
        i_data_bus[345]), .B2(n2625), .ZN(n2487) );
  ND4D1BWP30P140LVT U2883 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), 
        .ZN(n2496) );
  AOI22D1BWP30P140LVT U2884 ( .A1(i_data_bus[825]), .A2(n2635), .B1(
        i_data_bus[729]), .B2(n2640), .ZN(n2494) );
  AOI22D1BWP30P140LVT U2885 ( .A1(i_data_bus[761]), .A2(n2636), .B1(
        i_data_bus[889]), .B2(n2639), .ZN(n2493) );
  AOI22D1BWP30P140LVT U2886 ( .A1(i_data_bus[665]), .A2(n1989), .B1(
        i_data_bus[793]), .B2(n1986), .ZN(n2492) );
  AOI22D1BWP30P140LVT U2887 ( .A1(i_data_bus[697]), .A2(n2637), .B1(
        i_data_bus[857]), .B2(n2638), .ZN(n2491) );
  ND4D1BWP30P140LVT U2888 ( .A1(n2494), .A2(n2493), .A3(n2492), .A4(n2491), 
        .ZN(n2495) );
  OR4D1BWP30P140LVT U2889 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), 
        .Z(o_data_bus[153]) );
  AOI22D1BWP30P140LVT U2890 ( .A1(i_data_bus[602]), .A2(n2630), .B1(
        i_data_bus[506]), .B2(n2629), .ZN(n2502) );
  AOI22D1BWP30P140LVT U2891 ( .A1(i_data_bus[122]), .A2(n2623), .B1(
        i_data_bus[186]), .B2(n2605), .ZN(n2501) );
  AOI22D1BWP30P140LVT U2892 ( .A1(i_data_bus[90]), .A2(n2602), .B1(
        i_data_bus[218]), .B2(n2627), .ZN(n2500) );
  AOI22D1BWP30P140LVT U2893 ( .A1(i_data_bus[570]), .A2(n2618), .B1(
        i_data_bus[410]), .B2(n2614), .ZN(n2499) );
  ND4D1BWP30P140LVT U2894 ( .A1(n2502), .A2(n2501), .A3(n2500), .A4(n2499), 
        .ZN(n2518) );
  AOI22D1BWP30P140LVT U2895 ( .A1(i_data_bus[922]), .A2(n2612), .B1(
        i_data_bus[250]), .B2(n2603), .ZN(n2506) );
  AOI22D1BWP30P140LVT U2896 ( .A1(i_data_bus[954]), .A2(n2611), .B1(
        i_data_bus[634]), .B2(n2617), .ZN(n2505) );
  AOI22D1BWP30P140LVT U2897 ( .A1(i_data_bus[346]), .A2(n2625), .B1(
        i_data_bus[282]), .B2(n2606), .ZN(n2504) );
  AOI22D1BWP30P140LVT U2898 ( .A1(i_data_bus[1018]), .A2(n2616), .B1(
        i_data_bus[58]), .B2(n2628), .ZN(n2503) );
  ND4D1BWP30P140LVT U2899 ( .A1(n2506), .A2(n2505), .A3(n2504), .A4(n2503), 
        .ZN(n2517) );
  AOI22D1BWP30P140LVT U2900 ( .A1(i_data_bus[986]), .A2(n2626), .B1(
        i_data_bus[314]), .B2(n2604), .ZN(n2510) );
  AOI22D1BWP30P140LVT U2901 ( .A1(i_data_bus[154]), .A2(n2600), .B1(
        i_data_bus[378]), .B2(n2613), .ZN(n2509) );
  AOI22D1BWP30P140LVT U2902 ( .A1(i_data_bus[538]), .A2(n2601), .B1(
        i_data_bus[442]), .B2(n2615), .ZN(n2508) );
  AOI22D1BWP30P140LVT U2903 ( .A1(i_data_bus[26]), .A2(n2624), .B1(
        i_data_bus[474]), .B2(n2599), .ZN(n2507) );
  ND4D1BWP30P140LVT U2904 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), 
        .ZN(n2516) );
  AOI22D1BWP30P140LVT U2905 ( .A1(i_data_bus[826]), .A2(n2635), .B1(
        i_data_bus[890]), .B2(n2639), .ZN(n2514) );
  AOI22D1BWP30P140LVT U2906 ( .A1(i_data_bus[794]), .A2(n1986), .B1(
        i_data_bus[666]), .B2(n1989), .ZN(n2513) );
  AOI22D1BWP30P140LVT U2907 ( .A1(i_data_bus[858]), .A2(n2638), .B1(
        i_data_bus[762]), .B2(n2636), .ZN(n2512) );
  AOI22D1BWP30P140LVT U2908 ( .A1(i_data_bus[698]), .A2(n2637), .B1(
        i_data_bus[730]), .B2(n2640), .ZN(n2511) );
  ND4D1BWP30P140LVT U2909 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), 
        .ZN(n2515) );
  OR4D1BWP30P140LVT U2910 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), 
        .Z(o_data_bus[154]) );
  AOI22D1BWP30P140LVT U2911 ( .A1(i_data_bus[539]), .A2(n2601), .B1(
        i_data_bus[475]), .B2(n2599), .ZN(n2522) );
  AOI22D1BWP30P140LVT U2912 ( .A1(i_data_bus[635]), .A2(n2617), .B1(
        i_data_bus[27]), .B2(n2624), .ZN(n2521) );
  AOI22D1BWP30P140LVT U2913 ( .A1(i_data_bus[155]), .A2(n2600), .B1(
        i_data_bus[251]), .B2(n2603), .ZN(n2520) );
  AOI22D1BWP30P140LVT U2914 ( .A1(i_data_bus[379]), .A2(n2613), .B1(
        i_data_bus[347]), .B2(n2625), .ZN(n2519) );
  ND4D1BWP30P140LVT U2915 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), 
        .ZN(n2538) );
  AOI22D1BWP30P140LVT U2916 ( .A1(i_data_bus[59]), .A2(n2628), .B1(
        i_data_bus[315]), .B2(n2604), .ZN(n2526) );
  AOI22D1BWP30P140LVT U2917 ( .A1(i_data_bus[603]), .A2(n2630), .B1(
        i_data_bus[923]), .B2(n2612), .ZN(n2525) );
  AOI22D1BWP30P140LVT U2918 ( .A1(i_data_bus[571]), .A2(n2618), .B1(
        i_data_bus[283]), .B2(n2606), .ZN(n2524) );
  AOI22D1BWP30P140LVT U2919 ( .A1(i_data_bus[987]), .A2(n2626), .B1(
        i_data_bus[187]), .B2(n2605), .ZN(n2523) );
  ND4D1BWP30P140LVT U2920 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), 
        .ZN(n2537) );
  AOI22D1BWP30P140LVT U2921 ( .A1(i_data_bus[123]), .A2(n2623), .B1(
        i_data_bus[1019]), .B2(n2616), .ZN(n2530) );
  AOI22D1BWP30P140LVT U2922 ( .A1(i_data_bus[955]), .A2(n2611), .B1(
        i_data_bus[411]), .B2(n2614), .ZN(n2529) );
  AOI22D1BWP30P140LVT U2923 ( .A1(i_data_bus[91]), .A2(n2602), .B1(
        i_data_bus[443]), .B2(n2615), .ZN(n2528) );
  AOI22D1BWP30P140LVT U2924 ( .A1(i_data_bus[507]), .A2(n2629), .B1(
        i_data_bus[219]), .B2(n2627), .ZN(n2527) );
  ND4D1BWP30P140LVT U2925 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), 
        .ZN(n2536) );
  AOI22D1BWP30P140LVT U2926 ( .A1(i_data_bus[763]), .A2(n2636), .B1(
        i_data_bus[699]), .B2(n2637), .ZN(n2534) );
  AOI22D1BWP30P140LVT U2927 ( .A1(i_data_bus[795]), .A2(n1986), .B1(
        i_data_bus[859]), .B2(n2638), .ZN(n2533) );
  AOI22D1BWP30P140LVT U2928 ( .A1(i_data_bus[827]), .A2(n2635), .B1(
        i_data_bus[667]), .B2(n1989), .ZN(n2532) );
  AOI22D1BWP30P140LVT U2929 ( .A1(i_data_bus[731]), .A2(n2640), .B1(
        i_data_bus[891]), .B2(n2639), .ZN(n2531) );
  ND4D1BWP30P140LVT U2930 ( .A1(n2534), .A2(n2533), .A3(n2532), .A4(n2531), 
        .ZN(n2535) );
  OR4D1BWP30P140LVT U2931 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), 
        .Z(o_data_bus[155]) );
  AOI22D1BWP30P140LVT U2932 ( .A1(i_data_bus[1020]), .A2(n2616), .B1(
        i_data_bus[508]), .B2(n2629), .ZN(n2542) );
  AOI22D1BWP30P140LVT U2933 ( .A1(i_data_bus[92]), .A2(n2602), .B1(
        i_data_bus[412]), .B2(n2614), .ZN(n2541) );
  AOI22D1BWP30P140LVT U2934 ( .A1(i_data_bus[604]), .A2(n2630), .B1(
        i_data_bus[348]), .B2(n2625), .ZN(n2540) );
  AOI22D1BWP30P140LVT U2935 ( .A1(i_data_bus[540]), .A2(n2601), .B1(
        i_data_bus[220]), .B2(n2627), .ZN(n2539) );
  ND4D1BWP30P140LVT U2936 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), 
        .ZN(n2558) );
  AOI22D1BWP30P140LVT U2937 ( .A1(i_data_bus[636]), .A2(n2617), .B1(
        i_data_bus[252]), .B2(n2603), .ZN(n2546) );
  AOI22D1BWP30P140LVT U2938 ( .A1(i_data_bus[476]), .A2(n2599), .B1(
        i_data_bus[316]), .B2(n2604), .ZN(n2545) );
  AOI22D1BWP30P140LVT U2939 ( .A1(i_data_bus[956]), .A2(n2611), .B1(
        i_data_bus[284]), .B2(n2606), .ZN(n2544) );
  AOI22D1BWP30P140LVT U2940 ( .A1(i_data_bus[28]), .A2(n2624), .B1(
        i_data_bus[572]), .B2(n2618), .ZN(n2543) );
  ND4D1BWP30P140LVT U2941 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), 
        .ZN(n2557) );
  AOI22D1BWP30P140LVT U2942 ( .A1(i_data_bus[988]), .A2(n2626), .B1(
        i_data_bus[380]), .B2(n2613), .ZN(n2550) );
  AOI22D1BWP30P140LVT U2943 ( .A1(i_data_bus[60]), .A2(n2628), .B1(
        i_data_bus[156]), .B2(n2600), .ZN(n2549) );
  AOI22D1BWP30P140LVT U2944 ( .A1(i_data_bus[924]), .A2(n2612), .B1(
        i_data_bus[444]), .B2(n2615), .ZN(n2548) );
  AOI22D1BWP30P140LVT U2945 ( .A1(i_data_bus[124]), .A2(n2623), .B1(
        i_data_bus[188]), .B2(n2605), .ZN(n2547) );
  ND4D1BWP30P140LVT U2946 ( .A1(n2550), .A2(n2549), .A3(n2548), .A4(n2547), 
        .ZN(n2556) );
  AOI22D1BWP30P140LVT U2947 ( .A1(i_data_bus[732]), .A2(n2640), .B1(
        i_data_bus[764]), .B2(n2636), .ZN(n2554) );
  AOI22D1BWP30P140LVT U2948 ( .A1(i_data_bus[796]), .A2(n1986), .B1(
        i_data_bus[700]), .B2(n2637), .ZN(n2553) );
  AOI22D1BWP30P140LVT U2949 ( .A1(i_data_bus[828]), .A2(n2635), .B1(
        i_data_bus[860]), .B2(n2638), .ZN(n2552) );
  AOI22D1BWP30P140LVT U2950 ( .A1(i_data_bus[892]), .A2(n2639), .B1(
        i_data_bus[668]), .B2(n1989), .ZN(n2551) );
  ND4D1BWP30P140LVT U2951 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), 
        .ZN(n2555) );
  OR4D1BWP30P140LVT U2952 ( .A1(n2558), .A2(n2557), .A3(n2556), .A4(n2555), 
        .Z(o_data_bus[156]) );
  AOI22D1BWP30P140LVT U2953 ( .A1(i_data_bus[637]), .A2(n2617), .B1(
        i_data_bus[541]), .B2(n2601), .ZN(n2562) );
  AOI22D1BWP30P140LVT U2954 ( .A1(i_data_bus[29]), .A2(n2624), .B1(
        i_data_bus[285]), .B2(n2606), .ZN(n2561) );
  AOI22D1BWP30P140LVT U2955 ( .A1(i_data_bus[477]), .A2(n2599), .B1(
        i_data_bus[413]), .B2(n2614), .ZN(n2560) );
  AOI22D1BWP30P140LVT U2956 ( .A1(i_data_bus[957]), .A2(n2611), .B1(
        i_data_bus[93]), .B2(n2602), .ZN(n2559) );
  ND4D1BWP30P140LVT U2957 ( .A1(n2562), .A2(n2561), .A3(n2560), .A4(n2559), 
        .ZN(n2578) );
  AOI22D1BWP30P140LVT U2958 ( .A1(i_data_bus[61]), .A2(n2628), .B1(
        i_data_bus[157]), .B2(n2600), .ZN(n2566) );
  AOI22D1BWP30P140LVT U2959 ( .A1(i_data_bus[125]), .A2(n2623), .B1(
        i_data_bus[445]), .B2(n2615), .ZN(n2565) );
  AOI22D1BWP30P140LVT U2960 ( .A1(i_data_bus[1021]), .A2(n2616), .B1(
        i_data_bus[349]), .B2(n2625), .ZN(n2564) );
  AOI22D1BWP30P140LVT U2961 ( .A1(i_data_bus[381]), .A2(n2613), .B1(
        i_data_bus[253]), .B2(n2603), .ZN(n2563) );
  ND4D1BWP30P140LVT U2962 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), 
        .ZN(n2577) );
  AOI22D1BWP30P140LVT U2963 ( .A1(i_data_bus[925]), .A2(n2612), .B1(
        i_data_bus[189]), .B2(n2605), .ZN(n2570) );
  AOI22D1BWP30P140LVT U2964 ( .A1(i_data_bus[573]), .A2(n2618), .B1(
        i_data_bus[317]), .B2(n2604), .ZN(n2569) );
  AOI22D1BWP30P140LVT U2965 ( .A1(i_data_bus[509]), .A2(n2629), .B1(
        i_data_bus[221]), .B2(n2627), .ZN(n2568) );
  AOI22D1BWP30P140LVT U2966 ( .A1(i_data_bus[989]), .A2(n2626), .B1(
        i_data_bus[605]), .B2(n2630), .ZN(n2567) );
  ND4D1BWP30P140LVT U2967 ( .A1(n2570), .A2(n2569), .A3(n2568), .A4(n2567), 
        .ZN(n2576) );
  AOI22D1BWP30P140LVT U2968 ( .A1(i_data_bus[765]), .A2(n2636), .B1(
        i_data_bus[797]), .B2(n1986), .ZN(n2574) );
  AOI22D1BWP30P140LVT U2969 ( .A1(i_data_bus[733]), .A2(n2640), .B1(
        i_data_bus[829]), .B2(n2635), .ZN(n2573) );
  AOI22D1BWP30P140LVT U2970 ( .A1(i_data_bus[861]), .A2(n2638), .B1(
        i_data_bus[893]), .B2(n2639), .ZN(n2572) );
  AOI22D1BWP30P140LVT U2971 ( .A1(i_data_bus[701]), .A2(n2637), .B1(
        i_data_bus[669]), .B2(n1989), .ZN(n2571) );
  ND4D1BWP30P140LVT U2972 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), 
        .ZN(n2575) );
  OR4D1BWP30P140LVT U2973 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), 
        .Z(o_data_bus[157]) );
  AOI22D1BWP30P140LVT U2974 ( .A1(i_data_bus[926]), .A2(n2612), .B1(
        i_data_bus[350]), .B2(n2625), .ZN(n2582) );
  AOI22D1BWP30P140LVT U2975 ( .A1(i_data_bus[318]), .A2(n2604), .B1(
        i_data_bus[158]), .B2(n2600), .ZN(n2581) );
  AOI22D1BWP30P140LVT U2976 ( .A1(i_data_bus[62]), .A2(n2628), .B1(
        i_data_bus[30]), .B2(n2624), .ZN(n2580) );
  AOI22D1BWP30P140LVT U2977 ( .A1(i_data_bus[958]), .A2(n2611), .B1(
        i_data_bus[94]), .B2(n2602), .ZN(n2579) );
  ND4D1BWP30P140LVT U2978 ( .A1(n2582), .A2(n2581), .A3(n2580), .A4(n2579), 
        .ZN(n2598) );
  AOI22D1BWP30P140LVT U2979 ( .A1(i_data_bus[1022]), .A2(n2616), .B1(
        i_data_bus[286]), .B2(n2606), .ZN(n2586) );
  AOI22D1BWP30P140LVT U2980 ( .A1(i_data_bus[990]), .A2(n2626), .B1(
        i_data_bus[382]), .B2(n2613), .ZN(n2585) );
  AOI22D1BWP30P140LVT U2981 ( .A1(i_data_bus[606]), .A2(n2630), .B1(
        i_data_bus[478]), .B2(n2599), .ZN(n2584) );
  AOI22D1BWP30P140LVT U2982 ( .A1(i_data_bus[222]), .A2(n2627), .B1(
        i_data_bus[446]), .B2(n2615), .ZN(n2583) );
  ND4D1BWP30P140LVT U2983 ( .A1(n2586), .A2(n2585), .A3(n2584), .A4(n2583), 
        .ZN(n2597) );
  AOI22D1BWP30P140LVT U2984 ( .A1(i_data_bus[574]), .A2(n2618), .B1(
        i_data_bus[510]), .B2(n2629), .ZN(n2590) );
  AOI22D1BWP30P140LVT U2985 ( .A1(i_data_bus[190]), .A2(n2605), .B1(
        i_data_bus[414]), .B2(n2614), .ZN(n2589) );
  AOI22D1BWP30P140LVT U2986 ( .A1(i_data_bus[542]), .A2(n2601), .B1(
        i_data_bus[126]), .B2(n2623), .ZN(n2588) );
  AOI22D1BWP30P140LVT U2987 ( .A1(i_data_bus[638]), .A2(n2617), .B1(
        i_data_bus[254]), .B2(n2603), .ZN(n2587) );
  ND4D1BWP30P140LVT U2988 ( .A1(n2590), .A2(n2589), .A3(n2588), .A4(n2587), 
        .ZN(n2596) );
  AOI22D1BWP30P140LVT U2989 ( .A1(i_data_bus[862]), .A2(n2638), .B1(
        i_data_bus[702]), .B2(n2637), .ZN(n2594) );
  AOI22D1BWP30P140LVT U2990 ( .A1(i_data_bus[670]), .A2(n1989), .B1(
        i_data_bus[734]), .B2(n2640), .ZN(n2593) );
  AOI22D1BWP30P140LVT U2991 ( .A1(i_data_bus[830]), .A2(n2635), .B1(
        i_data_bus[894]), .B2(n2639), .ZN(n2592) );
  AOI22D1BWP30P140LVT U2992 ( .A1(i_data_bus[798]), .A2(n1986), .B1(
        i_data_bus[766]), .B2(n2636), .ZN(n2591) );
  ND4D1BWP30P140LVT U2993 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), 
        .ZN(n2595) );
  OR4D1BWP30P140LVT U2994 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), 
        .Z(o_data_bus[158]) );
  AOI22D1BWP30P140LVT U2995 ( .A1(i_data_bus[159]), .A2(n2600), .B1(
        i_data_bus[479]), .B2(n2599), .ZN(n2610) );
  AOI22D1BWP30P140LVT U2996 ( .A1(i_data_bus[95]), .A2(n2602), .B1(
        i_data_bus[543]), .B2(n2601), .ZN(n2609) );
  AOI22D1BWP30P140LVT U2997 ( .A1(i_data_bus[319]), .A2(n2604), .B1(
        i_data_bus[255]), .B2(n2603), .ZN(n2608) );
  AOI22D1BWP30P140LVT U2998 ( .A1(i_data_bus[287]), .A2(n2606), .B1(
        i_data_bus[191]), .B2(n2605), .ZN(n2607) );
  ND4D1BWP30P140LVT U2999 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), 
        .ZN(n2648) );
  AOI22D1BWP30P140LVT U3000 ( .A1(i_data_bus[927]), .A2(n2612), .B1(
        i_data_bus[959]), .B2(n2611), .ZN(n2622) );
  AOI22D1BWP30P140LVT U3001 ( .A1(i_data_bus[415]), .A2(n2614), .B1(
        i_data_bus[383]), .B2(n2613), .ZN(n2621) );
  AOI22D1BWP30P140LVT U3002 ( .A1(i_data_bus[1023]), .A2(n2616), .B1(
        i_data_bus[447]), .B2(n2615), .ZN(n2620) );
  AOI22D1BWP30P140LVT U3003 ( .A1(i_data_bus[575]), .A2(n2618), .B1(
        i_data_bus[639]), .B2(n2617), .ZN(n2619) );
  ND4D1BWP30P140LVT U3004 ( .A1(n2622), .A2(n2621), .A3(n2620), .A4(n2619), 
        .ZN(n2647) );
  AOI22D1BWP30P140LVT U3005 ( .A1(i_data_bus[31]), .A2(n2624), .B1(
        i_data_bus[127]), .B2(n2623), .ZN(n2634) );
  AOI22D1BWP30P140LVT U3006 ( .A1(i_data_bus[991]), .A2(n2626), .B1(
        i_data_bus[351]), .B2(n2625), .ZN(n2633) );
  AOI22D1BWP30P140LVT U3007 ( .A1(i_data_bus[63]), .A2(n2628), .B1(
        i_data_bus[223]), .B2(n2627), .ZN(n2632) );
  AOI22D1BWP30P140LVT U3008 ( .A1(i_data_bus[607]), .A2(n2630), .B1(
        i_data_bus[511]), .B2(n2629), .ZN(n2631) );
  ND4D1BWP30P140LVT U3009 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), 
        .ZN(n2646) );
  AOI22D1BWP30P140LVT U3010 ( .A1(i_data_bus[767]), .A2(n2636), .B1(
        i_data_bus[831]), .B2(n2635), .ZN(n2644) );
  AOI22D1BWP30P140LVT U3011 ( .A1(i_data_bus[863]), .A2(n2638), .B1(
        i_data_bus[703]), .B2(n2637), .ZN(n2643) );
  AOI22D1BWP30P140LVT U3012 ( .A1(i_data_bus[799]), .A2(n1986), .B1(
        i_data_bus[671]), .B2(n1989), .ZN(n2642) );
  AOI22D1BWP30P140LVT U3013 ( .A1(i_data_bus[735]), .A2(n2640), .B1(
        i_data_bus[895]), .B2(n2639), .ZN(n2641) );
  ND4D1BWP30P140LVT U3014 ( .A1(n2644), .A2(n2643), .A3(n2642), .A4(n2641), 
        .ZN(n2645) );
  OR4D1BWP30P140LVT U3015 ( .A1(n2648), .A2(n2647), .A3(n2646), .A4(n2645), 
        .Z(o_data_bus[159]) );
  INR3D2BWP30P140LVT U3016 ( .A1(i_cmd[13]), .B1(n5442), .B2(n2656), .ZN(n3305) );
  INVD1BWP30P140LVT U3017 ( .I(i_cmd[5]), .ZN(n2649) );
  AOI22D1BWP30P140LVT U3018 ( .A1(i_data_bus[32]), .A2(n3305), .B1(
        i_data_bus[0]), .B2(n3319), .ZN(n2694) );
  NR3D0P7BWP30P140LVT U3019 ( .A1(n5473), .A2(n2650), .A3(n2668), .ZN(n3309)
         );
  INR3D2BWP30P140LVT U3020 ( .A1(i_cmd[85]), .B1(n4084), .B2(n2667), .ZN(n3306) );
  AOI22D1BWP30P140LVT U3021 ( .A1(i_data_bus[896]), .A2(n3309), .B1(
        i_data_bus[320]), .B2(n3306), .ZN(n2693) );
  INVD1BWP30P140LVT U3022 ( .I(i_cmd[37]), .ZN(n2652) );
  AOI22D1BWP30P140LVT U3023 ( .A1(i_data_bus[128]), .A2(n2935), .B1(
        i_data_bus[224]), .B2(n3328), .ZN(n2692) );
  AOI22D1BWP30P140LVT U3024 ( .A1(i_data_bus[832]), .A2(n3316), .B1(
        i_data_bus[672]), .B2(n2653), .ZN(n2663) );
  INR3D2BWP30P140LVT U3025 ( .A1(i_cmd[29]), .B1(n5446), .B2(n2656), .ZN(n3308) );
  INVD1BWP30P140LVT U3026 ( .I(i_cmd[69]), .ZN(n2654) );
  NR3D0P7BWP30P140LVT U3027 ( .A1(n5497), .A2(n2654), .A3(n2667), .ZN(n2655)
         );
  AOI22D1BWP30P140LVT U3028 ( .A1(i_data_bus[96]), .A2(n3308), .B1(
        i_data_bus[256]), .B2(n3318), .ZN(n2662) );
  INR3D2BWP30P140LVT U3029 ( .A1(i_cmd[21]), .B1(n5451), .B2(n2656), .ZN(n3317) );
  INVD1BWP30P140LVT U3030 ( .I(i_cmd[165]), .ZN(n2657) );
  NR3D0P7BWP30P140LVT U3031 ( .A1(n5455), .A2(n2657), .A3(n2666), .ZN(n2658)
         );
  AOI22D1BWP30P140LVT U3032 ( .A1(i_data_bus[64]), .A2(n3317), .B1(
        i_data_bus[640]), .B2(n3302), .ZN(n2661) );
  AOI22D1BWP30P140LVT U3033 ( .A1(i_data_bus[736]), .A2(n2659), .B1(
        i_data_bus[800]), .B2(n3304), .ZN(n2660) );
  ND4D1BWP30P140LVT U3034 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), 
        .ZN(n2690) );
  NR3D0P7BWP30P140LVT U3035 ( .A1(n5470), .A2(n2664), .A3(n2668), .ZN(n3320)
         );
  INR3D2BWP30P140LVT U3036 ( .A1(i_cmd[93]), .B1(n4074), .B2(n2667), .ZN(n3321) );
  AOI22D1BWP30P140LVT U3037 ( .A1(i_data_bus[992]), .A2(n58), .B1(
        i_data_bus[352]), .B2(n3321), .ZN(n2675) );
  NR3D0P7BWP30P140LVT U3038 ( .A1(n5486), .A2(n2665), .A3(n2668), .ZN(n3311)
         );
  INR3D2BWP30P140LVT U3039 ( .A1(i_cmd[181]), .B1(n5448), .B2(n2666), .ZN(
        n3310) );
  AOI22D1BWP30P140LVT U3040 ( .A1(i_data_bus[928]), .A2(n3311), .B1(
        i_data_bus[704]), .B2(n3310), .ZN(n2674) );
  INR3D2BWP30P140LVT U3041 ( .A1(i_cmd[77]), .B1(n4095), .B2(n2667), .ZN(n3322) );
  AOI22D1BWP30P140LVT U3042 ( .A1(i_data_bus[864]), .A2(n113), .B1(
        i_data_bus[288]), .B2(n3322), .ZN(n2673) );
  INVD1BWP30P140LVT U3043 ( .I(i_cmd[197]), .ZN(n2671) );
  AOI22D1BWP30P140LVT U3044 ( .A1(i_data_bus[960]), .A2(n3301), .B1(
        i_data_bus[768]), .B2(n3307), .ZN(n2672) );
  ND4D1BWP30P140LVT U3045 ( .A1(n2675), .A2(n2674), .A3(n2673), .A4(n2672), 
        .ZN(n2689) );
  INVD1BWP30P140LVT U3046 ( .I(i_data_bus[448]), .ZN(n3372) );
  ND3D1BWP30P140LVT U3047 ( .A1(i_valid[6]), .A2(i_cmd[53]), .A3(n2677), .ZN(
        n3125) );
  MOAI22D1BWP30P140LVT U3048 ( .A1(n3372), .A2(n3246), .B1(i_data_bus[192]), 
        .B2(n2676), .ZN(n2688) );
  ND3D1BWP30P140LVT U3049 ( .A1(i_valid[5]), .A2(i_cmd[45]), .A3(n2677), .ZN(
        n3327) );
  AOI22D1BWP30P140LVT U3050 ( .A1(i_data_bus[416]), .A2(n3303), .B1(
        i_data_bus[160]), .B2(n2678), .ZN(n2686) );
  INR3D0BWP30P140LVT U3051 ( .A1(n2680), .B1(n143), .B2(n5476), .ZN(n2679) );
  AOI22D1BWP30P140LVT U3052 ( .A1(i_data_bus[384]), .A2(n3), .B1(
        i_data_bus[480]), .B2(n3329), .ZN(n2685) );
  INR3D2BWP30P140LVT U3053 ( .A1(i_cmd[157]), .B1(n5478), .B2(n2682), .ZN(
        n3333) );
  AOI22D1BWP30P140LVT U3054 ( .A1(i_data_bus[512]), .A2(n3331), .B1(
        i_data_bus[608]), .B2(n3333), .ZN(n2684) );
  INR3D2BWP30P140LVT U3055 ( .A1(i_cmd[141]), .B1(n5479), .B2(n2682), .ZN(
        n3332) );
  INR3D2BWP30P140LVT U3056 ( .A1(i_cmd[149]), .B1(n5481), .B2(n2682), .ZN(
        n3334) );
  AOI22D1BWP30P140LVT U3057 ( .A1(i_data_bus[544]), .A2(n3332), .B1(
        i_data_bus[576]), .B2(n3334), .ZN(n2683) );
  ND4D1BWP30P140LVT U3058 ( .A1(n2686), .A2(n2685), .A3(n2684), .A4(n2683), 
        .ZN(n2687) );
  NR4D0BWP30P140LVT U3059 ( .A1(n2690), .A2(n2689), .A3(n2688), .A4(n2687), 
        .ZN(n2691) );
  ND4D1BWP30P140LVT U3060 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), 
        .ZN(o_data_bus[160]) );
  AOI22D1BWP30P140LVT U3061 ( .A1(i_data_bus[673]), .A2(n2653), .B1(
        i_data_bus[865]), .B2(n113), .ZN(n2714) );
  AOI22D1BWP30P140LVT U3062 ( .A1(i_data_bus[289]), .A2(n3322), .B1(
        i_data_bus[321]), .B2(n3306), .ZN(n2713) );
  AOI22D1BWP30P140LVT U3063 ( .A1(i_data_bus[161]), .A2(n2678), .B1(
        i_data_bus[193]), .B2(n2676), .ZN(n2712) );
  AOI22D1BWP30P140LVT U3064 ( .A1(i_data_bus[97]), .A2(n3308), .B1(
        i_data_bus[1]), .B2(n3319), .ZN(n2698) );
  AOI22D1BWP30P140LVT U3065 ( .A1(i_data_bus[897]), .A2(n3309), .B1(
        i_data_bus[641]), .B2(n3302), .ZN(n2697) );
  AOI22D1BWP30P140LVT U3066 ( .A1(i_data_bus[33]), .A2(n3305), .B1(
        i_data_bus[65]), .B2(n3317), .ZN(n2696) );
  ND4D1BWP30P140LVT U3067 ( .A1(n2698), .A2(n2697), .A3(n2696), .A4(n2695), 
        .ZN(n2710) );
  AOI22D1BWP30P140LVT U3068 ( .A1(i_data_bus[929]), .A2(n3311), .B1(
        i_data_bus[769]), .B2(n3307), .ZN(n2702) );
  AOI22D1BWP30P140LVT U3069 ( .A1(i_data_bus[993]), .A2(n59), .B1(
        i_data_bus[737]), .B2(n2659), .ZN(n2701) );
  AOI22D1BWP30P140LVT U3070 ( .A1(i_data_bus[705]), .A2(n3310), .B1(
        i_data_bus[353]), .B2(n3321), .ZN(n2700) );
  AOI22D1BWP30P140LVT U3071 ( .A1(i_data_bus[801]), .A2(n3304), .B1(
        i_data_bus[257]), .B2(n3318), .ZN(n2699) );
  ND4D1BWP30P140LVT U3072 ( .A1(n2702), .A2(n2701), .A3(n2700), .A4(n2699), 
        .ZN(n2709) );
  INVD1BWP30P140LVT U3073 ( .I(i_data_bus[481]), .ZN(n5514) );
  MOAI22D1BWP30P140LVT U3074 ( .A1(n5514), .A2(n3267), .B1(i_data_bus[449]), 
        .B2(n3330), .ZN(n2708) );
  AOI22D1BWP30P140LVT U3075 ( .A1(i_data_bus[417]), .A2(n3303), .B1(
        i_data_bus[129]), .B2(n2935), .ZN(n2706) );
  AOI22D1BWP30P140LVT U3076 ( .A1(i_data_bus[385]), .A2(n3), .B1(
        i_data_bus[225]), .B2(n3328), .ZN(n2705) );
  AOI22D1BWP30P140LVT U3077 ( .A1(i_data_bus[577]), .A2(n3334), .B1(
        i_data_bus[609]), .B2(n3333), .ZN(n2704) );
  AOI22D1BWP30P140LVT U3078 ( .A1(i_data_bus[545]), .A2(n3332), .B1(
        i_data_bus[513]), .B2(n3331), .ZN(n2703) );
  ND4D1BWP30P140LVT U3079 ( .A1(n2706), .A2(n2705), .A3(n2704), .A4(n2703), 
        .ZN(n2707) );
  NR4D0BWP30P140LVT U3080 ( .A1(n2710), .A2(n2709), .A3(n2708), .A4(n2707), 
        .ZN(n2711) );
  ND4D1BWP30P140LVT U3081 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), 
        .ZN(o_data_bus[161]) );
  AOI22D1BWP30P140LVT U3082 ( .A1(i_data_bus[962]), .A2(n3301), .B1(
        i_data_bus[258]), .B2(n3318), .ZN(n2734) );
  AOI22D1BWP30P140LVT U3083 ( .A1(i_data_bus[898]), .A2(n3309), .B1(
        i_data_bus[2]), .B2(n3319), .ZN(n2733) );
  AOI22D1BWP30P140LVT U3084 ( .A1(i_data_bus[482]), .A2(n3329), .B1(
        i_data_bus[418]), .B2(n3303), .ZN(n2732) );
  AOI22D1BWP30P140LVT U3085 ( .A1(i_data_bus[994]), .A2(n59), .B1(
        i_data_bus[706]), .B2(n3310), .ZN(n2718) );
  AOI22D1BWP30P140LVT U3086 ( .A1(i_data_bus[98]), .A2(n3308), .B1(
        i_data_bus[674]), .B2(n2653), .ZN(n2717) );
  AOI22D1BWP30P140LVT U3087 ( .A1(i_data_bus[66]), .A2(n3317), .B1(
        i_data_bus[322]), .B2(n3306), .ZN(n2716) );
  AOI22D1BWP30P140LVT U3088 ( .A1(i_data_bus[290]), .A2(n3322), .B1(
        i_data_bus[642]), .B2(n3302), .ZN(n2715) );
  ND4D1BWP30P140LVT U3089 ( .A1(n2718), .A2(n2717), .A3(n2716), .A4(n2715), 
        .ZN(n2730) );
  AOI22D1BWP30P140LVT U3090 ( .A1(i_data_bus[930]), .A2(n3311), .B1(
        i_data_bus[770]), .B2(n3307), .ZN(n2722) );
  AOI22D1BWP30P140LVT U3091 ( .A1(i_data_bus[834]), .A2(n3316), .B1(
        i_data_bus[738]), .B2(n2659), .ZN(n2721) );
  AOI22D1BWP30P140LVT U3092 ( .A1(i_data_bus[802]), .A2(n3304), .B1(
        i_data_bus[354]), .B2(n3321), .ZN(n2720) );
  AOI22D1BWP30P140LVT U3093 ( .A1(i_data_bus[34]), .A2(n3305), .B1(
        i_data_bus[866]), .B2(n113), .ZN(n2719) );
  ND4D1BWP30P140LVT U3094 ( .A1(n2722), .A2(n2721), .A3(n2720), .A4(n2719), 
        .ZN(n2729) );
  INVD1BWP30P140LVT U3095 ( .I(i_data_bus[194]), .ZN(n5536) );
  INVD1BWP30P140LVT U3096 ( .I(i_data_bus[450]), .ZN(n3425) );
  OAI22D1BWP30P140LVT U3097 ( .A1(n5536), .A2(n3125), .B1(n3425), .B2(n3246), 
        .ZN(n2728) );
  AOI22D1BWP30P140LVT U3098 ( .A1(i_data_bus[226]), .A2(n3328), .B1(
        i_data_bus[130]), .B2(n2935), .ZN(n2726) );
  AOI22D1BWP30P140LVT U3099 ( .A1(i_data_bus[162]), .A2(n2678), .B1(
        i_data_bus[386]), .B2(n3), .ZN(n2725) );
  AOI22D1BWP30P140LVT U3100 ( .A1(i_data_bus[546]), .A2(n3332), .B1(
        i_data_bus[610]), .B2(n3333), .ZN(n2724) );
  AOI22D1BWP30P140LVT U3101 ( .A1(i_data_bus[578]), .A2(n3334), .B1(
        i_data_bus[514]), .B2(n3331), .ZN(n2723) );
  ND4D1BWP30P140LVT U3102 ( .A1(n2726), .A2(n2725), .A3(n2724), .A4(n2723), 
        .ZN(n2727) );
  NR4D0BWP30P140LVT U3103 ( .A1(n2730), .A2(n2729), .A3(n2728), .A4(n2727), 
        .ZN(n2731) );
  ND4D1BWP30P140LVT U3104 ( .A1(n2734), .A2(n2733), .A3(n2732), .A4(n2731), 
        .ZN(o_data_bus[162]) );
  AOI22D1BWP30P140LVT U3105 ( .A1(i_data_bus[771]), .A2(n3307), .B1(
        i_data_bus[803]), .B2(n3304), .ZN(n2754) );
  AOI22D1BWP30P140LVT U3106 ( .A1(i_data_bus[867]), .A2(n113), .B1(
        i_data_bus[707]), .B2(n3310), .ZN(n2753) );
  AOI22D1BWP30P140LVT U3107 ( .A1(i_data_bus[387]), .A2(n3), .B1(
        i_data_bus[483]), .B2(n3329), .ZN(n2752) );
  AOI22D1BWP30P140LVT U3108 ( .A1(i_data_bus[355]), .A2(n3321), .B1(
        i_data_bus[291]), .B2(n3322), .ZN(n2738) );
  AOI22D1BWP30P140LVT U3109 ( .A1(i_data_bus[259]), .A2(n3318), .B1(
        i_data_bus[323]), .B2(n3306), .ZN(n2737) );
  AOI22D1BWP30P140LVT U3110 ( .A1(i_data_bus[995]), .A2(n59), .B1(
        i_data_bus[643]), .B2(n3302), .ZN(n2736) );
  ND4D1BWP30P140LVT U3111 ( .A1(n2738), .A2(n2737), .A3(n2736), .A4(n2735), 
        .ZN(n2750) );
  AOI22D1BWP30P140LVT U3112 ( .A1(i_data_bus[67]), .A2(n3317), .B1(
        i_data_bus[675]), .B2(n2653), .ZN(n2742) );
  AOI22D1BWP30P140LVT U3113 ( .A1(i_data_bus[899]), .A2(n3309), .B1(
        i_data_bus[3]), .B2(n3319), .ZN(n2741) );
  AOI22D1BWP30P140LVT U3114 ( .A1(i_data_bus[931]), .A2(n3311), .B1(
        i_data_bus[739]), .B2(n2659), .ZN(n2740) );
  AOI22D1BWP30P140LVT U3115 ( .A1(i_data_bus[35]), .A2(n3305), .B1(
        i_data_bus[963]), .B2(n3301), .ZN(n2739) );
  ND4D1BWP30P140LVT U3116 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), 
        .ZN(n2749) );
  INVD1BWP30P140LVT U3117 ( .I(i_data_bus[131]), .ZN(n5557) );
  INVD1BWP30P140LVT U3118 ( .I(i_data_bus[451]), .ZN(n3446) );
  OAI22D1BWP30P140LVT U3119 ( .A1(n5557), .A2(n3044), .B1(n3446), .B2(n3246), 
        .ZN(n2748) );
  AOI22D1BWP30P140LVT U3120 ( .A1(i_data_bus[163]), .A2(n2678), .B1(
        i_data_bus[195]), .B2(n2676), .ZN(n2746) );
  AOI22D1BWP30P140LVT U3121 ( .A1(i_data_bus[419]), .A2(n3303), .B1(
        i_data_bus[227]), .B2(n3328), .ZN(n2745) );
  AOI22D1BWP30P140LVT U3122 ( .A1(i_data_bus[515]), .A2(n3331), .B1(
        i_data_bus[547]), .B2(n3332), .ZN(n2744) );
  AOI22D1BWP30P140LVT U3123 ( .A1(i_data_bus[579]), .A2(n3334), .B1(
        i_data_bus[611]), .B2(n3333), .ZN(n2743) );
  ND4D1BWP30P140LVT U3124 ( .A1(n2746), .A2(n2745), .A3(n2744), .A4(n2743), 
        .ZN(n2747) );
  NR4D0BWP30P140LVT U3125 ( .A1(n2750), .A2(n2749), .A3(n2748), .A4(n2747), 
        .ZN(n2751) );
  ND4D1BWP30P140LVT U3126 ( .A1(n2754), .A2(n2753), .A3(n2752), .A4(n2751), 
        .ZN(o_data_bus[163]) );
  AOI22D1BWP30P140LVT U3127 ( .A1(i_data_bus[4]), .A2(n3319), .B1(
        i_data_bus[740]), .B2(n2659), .ZN(n2774) );
  AOI22D1BWP30P140LVT U3128 ( .A1(i_data_bus[964]), .A2(n3301), .B1(
        i_data_bus[932]), .B2(n3311), .ZN(n2773) );
  AOI22D1BWP30P140LVT U3129 ( .A1(i_data_bus[132]), .A2(n2935), .B1(
        i_data_bus[420]), .B2(n3303), .ZN(n2772) );
  AOI22D1BWP30P140LVT U3130 ( .A1(i_data_bus[996]), .A2(n58), .B1(
        i_data_bus[324]), .B2(n3306), .ZN(n2758) );
  AOI22D1BWP30P140LVT U3131 ( .A1(i_data_bus[68]), .A2(n3317), .B1(
        i_data_bus[644]), .B2(n3302), .ZN(n2757) );
  AOI22D1BWP30P140LVT U3132 ( .A1(i_data_bus[356]), .A2(n3321), .B1(
        i_data_bus[260]), .B2(n3318), .ZN(n2755) );
  ND4D1BWP30P140LVT U3133 ( .A1(n2758), .A2(n2757), .A3(n2756), .A4(n2755), 
        .ZN(n2770) );
  AOI22D1BWP30P140LVT U3134 ( .A1(i_data_bus[772]), .A2(n3307), .B1(
        i_data_bus[804]), .B2(n3304), .ZN(n2762) );
  AOI22D1BWP30P140LVT U3135 ( .A1(i_data_bus[900]), .A2(n3309), .B1(
        i_data_bus[36]), .B2(n3305), .ZN(n2761) );
  AOI22D1BWP30P140LVT U3136 ( .A1(i_data_bus[100]), .A2(n3308), .B1(
        i_data_bus[868]), .B2(n113), .ZN(n2760) );
  AOI22D1BWP30P140LVT U3137 ( .A1(i_data_bus[708]), .A2(n3310), .B1(
        i_data_bus[292]), .B2(n3322), .ZN(n2759) );
  ND4D1BWP30P140LVT U3138 ( .A1(n2762), .A2(n2761), .A3(n2760), .A4(n2759), 
        .ZN(n2769) );
  INVD1BWP30P140LVT U3139 ( .I(i_data_bus[452]), .ZN(n5579) );
  INVD1BWP30P140LVT U3140 ( .I(i_data_bus[388]), .ZN(n3464) );
  OAI22D1BWP30P140LVT U3141 ( .A1(n5579), .A2(n3246), .B1(n3464), .B2(n3288), 
        .ZN(n2768) );
  AOI22D1BWP30P140LVT U3142 ( .A1(i_data_bus[228]), .A2(n3328), .B1(
        i_data_bus[164]), .B2(n2678), .ZN(n2766) );
  AOI22D1BWP30P140LVT U3143 ( .A1(i_data_bus[196]), .A2(n2676), .B1(
        i_data_bus[484]), .B2(n3329), .ZN(n2765) );
  AOI22D1BWP30P140LVT U3144 ( .A1(i_data_bus[548]), .A2(n3332), .B1(
        i_data_bus[612]), .B2(n3333), .ZN(n2764) );
  AOI22D1BWP30P140LVT U3145 ( .A1(i_data_bus[516]), .A2(n3331), .B1(
        i_data_bus[580]), .B2(n3334), .ZN(n2763) );
  ND4D1BWP30P140LVT U3146 ( .A1(n2766), .A2(n2765), .A3(n2764), .A4(n2763), 
        .ZN(n2767) );
  NR4D0BWP30P140LVT U3147 ( .A1(n2770), .A2(n2769), .A3(n2768), .A4(n2767), 
        .ZN(n2771) );
  ND4D1BWP30P140LVT U3148 ( .A1(n2774), .A2(n2773), .A3(n2772), .A4(n2771), 
        .ZN(o_data_bus[164]) );
  AOI22D1BWP30P140LVT U3149 ( .A1(i_data_bus[901]), .A2(n3309), .B1(
        i_data_bus[869]), .B2(n113), .ZN(n2794) );
  AOI22D1BWP30P140LVT U3150 ( .A1(i_data_bus[997]), .A2(n59), .B1(
        i_data_bus[805]), .B2(n3304), .ZN(n2793) );
  AOI22D1BWP30P140LVT U3151 ( .A1(i_data_bus[165]), .A2(n2678), .B1(
        i_data_bus[485]), .B2(n3329), .ZN(n2792) );
  AOI22D1BWP30P140LVT U3152 ( .A1(i_data_bus[197]), .A2(n2676), .B1(
        i_data_bus[133]), .B2(n2935), .ZN(n2790) );
  AOI22D1BWP30P140LVT U3153 ( .A1(i_data_bus[933]), .A2(n3311), .B1(
        i_data_bus[69]), .B2(n3317), .ZN(n2777) );
  AOI22D1BWP30P140LVT U3154 ( .A1(i_data_bus[773]), .A2(n3307), .B1(
        i_data_bus[709]), .B2(n3310), .ZN(n2776) );
  AOI22D1BWP30P140LVT U3155 ( .A1(i_data_bus[965]), .A2(n3301), .B1(
        i_data_bus[293]), .B2(n3322), .ZN(n2775) );
  ND4D1BWP30P140LVT U3156 ( .A1(n2778), .A2(n2777), .A3(n2776), .A4(n2775), 
        .ZN(n2789) );
  AOI22D1BWP30P140LVT U3157 ( .A1(i_data_bus[5]), .A2(n3319), .B1(
        i_data_bus[261]), .B2(n3318), .ZN(n2782) );
  AOI22D1BWP30P140LVT U3158 ( .A1(i_data_bus[645]), .A2(n3302), .B1(
        i_data_bus[741]), .B2(n2659), .ZN(n2781) );
  AOI22D1BWP30P140LVT U3159 ( .A1(i_data_bus[101]), .A2(n3308), .B1(
        i_data_bus[357]), .B2(n3321), .ZN(n2780) );
  AOI22D1BWP30P140LVT U3160 ( .A1(i_data_bus[37]), .A2(n3305), .B1(
        i_data_bus[325]), .B2(n3306), .ZN(n2779) );
  ND4D1BWP30P140LVT U3161 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), 
        .ZN(n2788) );
  AOI22D1BWP30P140LVT U3162 ( .A1(i_data_bus[421]), .A2(n3303), .B1(
        i_data_bus[389]), .B2(n3), .ZN(n2786) );
  AOI22D1BWP30P140LVT U3163 ( .A1(i_data_bus[453]), .A2(n3330), .B1(
        i_data_bus[229]), .B2(n3328), .ZN(n2785) );
  AOI22D1BWP30P140LVT U3164 ( .A1(i_data_bus[517]), .A2(n3331), .B1(
        i_data_bus[549]), .B2(n3332), .ZN(n2784) );
  AOI22D1BWP30P140LVT U3165 ( .A1(i_data_bus[581]), .A2(n3334), .B1(
        i_data_bus[613]), .B2(n3333), .ZN(n2783) );
  ND4D1BWP30P140LVT U3166 ( .A1(n2786), .A2(n2785), .A3(n2784), .A4(n2783), 
        .ZN(n2787) );
  INR4D0BWP30P140LVT U3167 ( .A1(n2790), .B1(n2789), .B2(n2788), .B3(n2787), 
        .ZN(n2791) );
  ND4D1BWP30P140LVT U3168 ( .A1(n2794), .A2(n2793), .A3(n2792), .A4(n2791), 
        .ZN(o_data_bus[165]) );
  AOI22D1BWP30P140LVT U3169 ( .A1(i_data_bus[6]), .A2(n3319), .B1(
        i_data_bus[838]), .B2(n3316), .ZN(n2814) );
  AOI22D1BWP30P140LVT U3170 ( .A1(i_data_bus[998]), .A2(n58), .B1(
        i_data_bus[678]), .B2(n2653), .ZN(n2813) );
  AOI22D1BWP30P140LVT U3171 ( .A1(i_data_bus[230]), .A2(n3328), .B1(
        i_data_bus[422]), .B2(n3303), .ZN(n2812) );
  AOI22D1BWP30P140LVT U3172 ( .A1(i_data_bus[742]), .A2(n2659), .B1(
        i_data_bus[774]), .B2(n3307), .ZN(n2798) );
  AOI22D1BWP30P140LVT U3173 ( .A1(i_data_bus[966]), .A2(n3301), .B1(
        i_data_bus[262]), .B2(n3318), .ZN(n2797) );
  AOI22D1BWP30P140LVT U3174 ( .A1(i_data_bus[102]), .A2(n3308), .B1(
        i_data_bus[806]), .B2(n3304), .ZN(n2796) );
  AOI22D1BWP30P140LVT U3175 ( .A1(i_data_bus[710]), .A2(n3310), .B1(
        i_data_bus[294]), .B2(n3322), .ZN(n2795) );
  ND4D1BWP30P140LVT U3176 ( .A1(n2798), .A2(n2797), .A3(n2796), .A4(n2795), 
        .ZN(n2810) );
  AOI22D1BWP30P140LVT U3177 ( .A1(i_data_bus[902]), .A2(n3309), .B1(
        i_data_bus[358]), .B2(n3321), .ZN(n2802) );
  AOI22D1BWP30P140LVT U3178 ( .A1(i_data_bus[934]), .A2(n3311), .B1(
        i_data_bus[870]), .B2(n113), .ZN(n2801) );
  AOI22D1BWP30P140LVT U3179 ( .A1(i_data_bus[38]), .A2(n3305), .B1(
        i_data_bus[70]), .B2(n3317), .ZN(n2800) );
  AOI22D1BWP30P140LVT U3180 ( .A1(i_data_bus[646]), .A2(n3302), .B1(
        i_data_bus[326]), .B2(n3306), .ZN(n2799) );
  ND4D1BWP30P140LVT U3181 ( .A1(n2802), .A2(n2801), .A3(n2800), .A4(n2799), 
        .ZN(n2809) );
  INVD1BWP30P140LVT U3182 ( .I(i_data_bus[454]), .ZN(n5621) );
  MOAI22D1BWP30P140LVT U3183 ( .A1(n5621), .A2(n3246), .B1(i_data_bus[198]), 
        .B2(n2676), .ZN(n2808) );
  AOI22D1BWP30P140LVT U3184 ( .A1(i_data_bus[486]), .A2(n3329), .B1(
        i_data_bus[390]), .B2(n3), .ZN(n2806) );
  AOI22D1BWP30P140LVT U3185 ( .A1(i_data_bus[166]), .A2(n2678), .B1(
        i_data_bus[134]), .B2(n2935), .ZN(n2805) );
  AOI22D1BWP30P140LVT U3186 ( .A1(i_data_bus[582]), .A2(n3334), .B1(
        i_data_bus[518]), .B2(n3331), .ZN(n2804) );
  AOI22D1BWP30P140LVT U3187 ( .A1(i_data_bus[614]), .A2(n3333), .B1(
        i_data_bus[550]), .B2(n3332), .ZN(n2803) );
  ND4D1BWP30P140LVT U3188 ( .A1(n2806), .A2(n2805), .A3(n2804), .A4(n2803), 
        .ZN(n2807) );
  NR4D0BWP30P140LVT U3189 ( .A1(n2810), .A2(n2809), .A3(n2808), .A4(n2807), 
        .ZN(n2811) );
  ND4D1BWP30P140LVT U3190 ( .A1(n2814), .A2(n2813), .A3(n2812), .A4(n2811), 
        .ZN(o_data_bus[166]) );
  AOI22D1BWP30P140LVT U3191 ( .A1(i_data_bus[775]), .A2(n3307), .B1(
        i_data_bus[295]), .B2(n3322), .ZN(n2834) );
  AOI22D1BWP30P140LVT U3192 ( .A1(i_data_bus[967]), .A2(n3301), .B1(
        i_data_bus[935]), .B2(n3311), .ZN(n2833) );
  AOI22D1BWP30P140LVT U3193 ( .A1(i_data_bus[391]), .A2(n3), .B1(
        i_data_bus[135]), .B2(n2935), .ZN(n2832) );
  AOI22D1BWP30P140LVT U3194 ( .A1(i_data_bus[871]), .A2(n113), .B1(
        i_data_bus[679]), .B2(n2653), .ZN(n2818) );
  AOI22D1BWP30P140LVT U3195 ( .A1(i_data_bus[359]), .A2(n3321), .B1(
        i_data_bus[327]), .B2(n3306), .ZN(n2817) );
  AOI22D1BWP30P140LVT U3196 ( .A1(i_data_bus[263]), .A2(n3318), .B1(
        i_data_bus[807]), .B2(n3304), .ZN(n2816) );
  AOI22D1BWP30P140LVT U3197 ( .A1(i_data_bus[7]), .A2(n3319), .B1(
        i_data_bus[71]), .B2(n3317), .ZN(n2815) );
  ND4D1BWP30P140LVT U3198 ( .A1(n2818), .A2(n2817), .A3(n2816), .A4(n2815), 
        .ZN(n2830) );
  AOI22D1BWP30P140LVT U3199 ( .A1(i_data_bus[839]), .A2(n3316), .B1(
        i_data_bus[647]), .B2(n3302), .ZN(n2822) );
  AOI22D1BWP30P140LVT U3200 ( .A1(i_data_bus[903]), .A2(n3309), .B1(
        i_data_bus[743]), .B2(n2659), .ZN(n2821) );
  AOI22D1BWP30P140LVT U3201 ( .A1(i_data_bus[103]), .A2(n3308), .B1(
        i_data_bus[999]), .B2(n3320), .ZN(n2820) );
  AOI22D1BWP30P140LVT U3202 ( .A1(i_data_bus[39]), .A2(n3305), .B1(
        i_data_bus[711]), .B2(n3310), .ZN(n2819) );
  ND4D1BWP30P140LVT U3203 ( .A1(n2822), .A2(n2821), .A3(n2820), .A4(n2819), 
        .ZN(n2829) );
  INVD1BWP30P140LVT U3204 ( .I(i_data_bus[487]), .ZN(n3525) );
  INVD1BWP30P140LVT U3205 ( .I(i_data_bus[199]), .ZN(n5642) );
  OAI22D1BWP30P140LVT U3206 ( .A1(n3525), .A2(n3267), .B1(n5642), .B2(n3125), 
        .ZN(n2828) );
  AOI22D1BWP30P140LVT U3207 ( .A1(i_data_bus[167]), .A2(n2678), .B1(
        i_data_bus[231]), .B2(n3328), .ZN(n2826) );
  AOI22D1BWP30P140LVT U3208 ( .A1(i_data_bus[455]), .A2(n3330), .B1(
        i_data_bus[423]), .B2(n3303), .ZN(n2825) );
  AOI22D1BWP30P140LVT U3209 ( .A1(i_data_bus[615]), .A2(n3333), .B1(
        i_data_bus[551]), .B2(n3332), .ZN(n2824) );
  AOI22D1BWP30P140LVT U3210 ( .A1(i_data_bus[519]), .A2(n3331), .B1(
        i_data_bus[583]), .B2(n3334), .ZN(n2823) );
  ND4D1BWP30P140LVT U3211 ( .A1(n2826), .A2(n2825), .A3(n2824), .A4(n2823), 
        .ZN(n2827) );
  NR4D0BWP30P140LVT U3212 ( .A1(n2830), .A2(n2829), .A3(n2828), .A4(n2827), 
        .ZN(n2831) );
  ND4D1BWP30P140LVT U3213 ( .A1(n2834), .A2(n2833), .A3(n2832), .A4(n2831), 
        .ZN(o_data_bus[167]) );
  AOI22D1BWP30P140LVT U3214 ( .A1(i_data_bus[936]), .A2(n7), .B1(
        i_data_bus[808]), .B2(n3304), .ZN(n2854) );
  AOI22D1BWP30P140LVT U3215 ( .A1(i_data_bus[904]), .A2(n3309), .B1(
        i_data_bus[40]), .B2(n3305), .ZN(n2853) );
  AOI22D1BWP30P140LVT U3216 ( .A1(i_data_bus[456]), .A2(n3330), .B1(
        i_data_bus[488]), .B2(n3329), .ZN(n2852) );
  AOI22D1BWP30P140LVT U3217 ( .A1(i_data_bus[200]), .A2(n2676), .B1(
        i_data_bus[136]), .B2(n2935), .ZN(n2850) );
  AOI22D1BWP30P140LVT U3218 ( .A1(i_data_bus[104]), .A2(n3308), .B1(
        i_data_bus[1000]), .B2(n3320), .ZN(n2838) );
  AOI22D1BWP30P140LVT U3219 ( .A1(i_data_bus[72]), .A2(n3317), .B1(
        i_data_bus[712]), .B2(n3310), .ZN(n2837) );
  AOI22D1BWP30P140LVT U3220 ( .A1(i_data_bus[840]), .A2(n3316), .B1(
        i_data_bus[648]), .B2(n3302), .ZN(n2836) );
  AOI22D1BWP30P140LVT U3221 ( .A1(i_data_bus[968]), .A2(n3301), .B1(
        i_data_bus[328]), .B2(n3306), .ZN(n2835) );
  ND4D1BWP30P140LVT U3222 ( .A1(n2838), .A2(n2837), .A3(n2836), .A4(n2835), 
        .ZN(n2849) );
  AOI22D1BWP30P140LVT U3223 ( .A1(i_data_bus[8]), .A2(n3319), .B1(
        i_data_bus[776]), .B2(n3307), .ZN(n2842) );
  AOI22D1BWP30P140LVT U3224 ( .A1(i_data_bus[744]), .A2(n2659), .B1(
        i_data_bus[680]), .B2(n2653), .ZN(n2841) );
  AOI22D1BWP30P140LVT U3225 ( .A1(i_data_bus[264]), .A2(n3318), .B1(
        i_data_bus[872]), .B2(n113), .ZN(n2840) );
  AOI22D1BWP30P140LVT U3226 ( .A1(i_data_bus[296]), .A2(n3322), .B1(
        i_data_bus[360]), .B2(n3321), .ZN(n2839) );
  ND4D1BWP30P140LVT U3227 ( .A1(n2842), .A2(n2841), .A3(n2840), .A4(n2839), 
        .ZN(n2848) );
  AOI22D1BWP30P140LVT U3228 ( .A1(i_data_bus[424]), .A2(n3303), .B1(
        i_data_bus[392]), .B2(n3), .ZN(n2846) );
  AOI22D1BWP30P140LVT U3229 ( .A1(i_data_bus[168]), .A2(n2678), .B1(
        i_data_bus[232]), .B2(n3328), .ZN(n2845) );
  AOI22D1BWP30P140LVT U3230 ( .A1(i_data_bus[616]), .A2(n3333), .B1(
        i_data_bus[552]), .B2(n3332), .ZN(n2844) );
  AOI22D1BWP30P140LVT U3231 ( .A1(i_data_bus[584]), .A2(n3334), .B1(
        i_data_bus[520]), .B2(n3331), .ZN(n2843) );
  ND4D1BWP30P140LVT U3232 ( .A1(n2846), .A2(n2845), .A3(n2844), .A4(n2843), 
        .ZN(n2847) );
  INR4D0BWP30P140LVT U3233 ( .A1(n2850), .B1(n2849), .B2(n2848), .B3(n2847), 
        .ZN(n2851) );
  ND4D1BWP30P140LVT U3234 ( .A1(n2854), .A2(n2853), .A3(n2852), .A4(n2851), 
        .ZN(o_data_bus[168]) );
  AOI22D1BWP30P140LVT U3235 ( .A1(i_data_bus[105]), .A2(n3308), .B1(
        i_data_bus[41]), .B2(n3305), .ZN(n2874) );
  AOI22D1BWP30P140LVT U3236 ( .A1(i_data_bus[969]), .A2(n3301), .B1(
        i_data_bus[713]), .B2(n3310), .ZN(n2873) );
  AOI22D1BWP30P140LVT U3237 ( .A1(i_data_bus[233]), .A2(n3328), .B1(
        i_data_bus[457]), .B2(n3330), .ZN(n2872) );
  AOI22D1BWP30P140LVT U3238 ( .A1(i_data_bus[873]), .A2(n113), .B1(
        i_data_bus[649]), .B2(n3302), .ZN(n2858) );
  AOI22D1BWP30P140LVT U3239 ( .A1(i_data_bus[1001]), .A2(n59), .B1(
        i_data_bus[361]), .B2(n3321), .ZN(n2857) );
  AOI22D1BWP30P140LVT U3240 ( .A1(i_data_bus[745]), .A2(n2659), .B1(
        i_data_bus[297]), .B2(n3322), .ZN(n2856) );
  AOI22D1BWP30P140LVT U3241 ( .A1(i_data_bus[681]), .A2(n2653), .B1(
        i_data_bus[809]), .B2(n3304), .ZN(n2855) );
  ND4D1BWP30P140LVT U3242 ( .A1(n2858), .A2(n2857), .A3(n2856), .A4(n2855), 
        .ZN(n2870) );
  AOI22D1BWP30P140LVT U3243 ( .A1(i_data_bus[9]), .A2(n3319), .B1(
        i_data_bus[329]), .B2(n3306), .ZN(n2862) );
  AOI22D1BWP30P140LVT U3244 ( .A1(i_data_bus[905]), .A2(n3309), .B1(
        i_data_bus[73]), .B2(n3317), .ZN(n2861) );
  AOI22D1BWP30P140LVT U3245 ( .A1(i_data_bus[937]), .A2(n3311), .B1(
        i_data_bus[265]), .B2(n3318), .ZN(n2860) );
  ND4D1BWP30P140LVT U3246 ( .A1(n2862), .A2(n2861), .A3(n2860), .A4(n2859), 
        .ZN(n2869) );
  INVD1BWP30P140LVT U3247 ( .I(i_data_bus[489]), .ZN(n4953) );
  INVD1BWP30P140LVT U3248 ( .I(i_data_bus[393]), .ZN(n3570) );
  OAI22D1BWP30P140LVT U3249 ( .A1(n4953), .A2(n3267), .B1(n3570), .B2(n3288), 
        .ZN(n2868) );
  AOI22D1BWP30P140LVT U3250 ( .A1(i_data_bus[201]), .A2(n2676), .B1(
        i_data_bus[425]), .B2(n3303), .ZN(n2866) );
  AOI22D1BWP30P140LVT U3251 ( .A1(i_data_bus[169]), .A2(n2678), .B1(
        i_data_bus[137]), .B2(n2935), .ZN(n2865) );
  AOI22D1BWP30P140LVT U3252 ( .A1(i_data_bus[521]), .A2(n3331), .B1(
        i_data_bus[617]), .B2(n3333), .ZN(n2864) );
  AOI22D1BWP30P140LVT U3253 ( .A1(i_data_bus[585]), .A2(n3334), .B1(
        i_data_bus[553]), .B2(n3332), .ZN(n2863) );
  ND4D1BWP30P140LVT U3254 ( .A1(n2866), .A2(n2865), .A3(n2864), .A4(n2863), 
        .ZN(n2867) );
  NR4D0BWP30P140LVT U3255 ( .A1(n2870), .A2(n2869), .A3(n2868), .A4(n2867), 
        .ZN(n2871) );
  ND4D1BWP30P140LVT U3256 ( .A1(n2874), .A2(n2873), .A3(n2872), .A4(n2871), 
        .ZN(o_data_bus[169]) );
  AOI22D1BWP30P140LVT U3257 ( .A1(i_data_bus[874]), .A2(n113), .B1(
        i_data_bus[714]), .B2(n3310), .ZN(n2894) );
  AOI22D1BWP30P140LVT U3258 ( .A1(i_data_bus[362]), .A2(n3321), .B1(
        i_data_bus[810]), .B2(n3304), .ZN(n2893) );
  AOI22D1BWP30P140LVT U3259 ( .A1(i_data_bus[490]), .A2(n3329), .B1(
        i_data_bus[138]), .B2(n2935), .ZN(n2892) );
  AOI22D1BWP30P140LVT U3260 ( .A1(i_data_bus[106]), .A2(n3308), .B1(
        i_data_bus[74]), .B2(n3317), .ZN(n2878) );
  AOI22D1BWP30P140LVT U3261 ( .A1(i_data_bus[970]), .A2(n3301), .B1(
        i_data_bus[266]), .B2(n3318), .ZN(n2877) );
  AOI22D1BWP30P140LVT U3262 ( .A1(i_data_bus[1002]), .A2(n59), .B1(
        i_data_bus[42]), .B2(n3305), .ZN(n2875) );
  ND4D1BWP30P140LVT U3263 ( .A1(n2878), .A2(n2877), .A3(n2876), .A4(n2875), 
        .ZN(n2890) );
  AOI22D1BWP30P140LVT U3264 ( .A1(i_data_bus[938]), .A2(n3311), .B1(
        i_data_bus[330]), .B2(n3306), .ZN(n2882) );
  AOI22D1BWP30P140LVT U3265 ( .A1(i_data_bus[650]), .A2(n3302), .B1(
        i_data_bus[298]), .B2(n3322), .ZN(n2881) );
  AOI22D1BWP30P140LVT U3266 ( .A1(i_data_bus[10]), .A2(n3319), .B1(
        i_data_bus[746]), .B2(n2659), .ZN(n2880) );
  AOI22D1BWP30P140LVT U3267 ( .A1(i_data_bus[906]), .A2(n3309), .B1(
        i_data_bus[682]), .B2(n2653), .ZN(n2879) );
  ND4D1BWP30P140LVT U3268 ( .A1(n2882), .A2(n2881), .A3(n2880), .A4(n2879), 
        .ZN(n2889) );
  INVD1BWP30P140LVT U3269 ( .I(i_data_bus[394]), .ZN(n5705) );
  MOAI22D1BWP30P140LVT U3270 ( .A1(n5705), .A2(n3288), .B1(i_data_bus[202]), 
        .B2(n2676), .ZN(n2888) );
  AOI22D1BWP30P140LVT U3271 ( .A1(i_data_bus[170]), .A2(n2678), .B1(
        i_data_bus[426]), .B2(n3303), .ZN(n2886) );
  AOI22D1BWP30P140LVT U3272 ( .A1(i_data_bus[234]), .A2(n3328), .B1(
        i_data_bus[458]), .B2(n3330), .ZN(n2885) );
  AOI22D1BWP30P140LVT U3273 ( .A1(i_data_bus[554]), .A2(n3332), .B1(
        i_data_bus[522]), .B2(n3331), .ZN(n2884) );
  AOI22D1BWP30P140LVT U3274 ( .A1(i_data_bus[618]), .A2(n3333), .B1(
        i_data_bus[586]), .B2(n3334), .ZN(n2883) );
  ND4D1BWP30P140LVT U3275 ( .A1(n2886), .A2(n2885), .A3(n2884), .A4(n2883), 
        .ZN(n2887) );
  NR4D0BWP30P140LVT U3276 ( .A1(n2890), .A2(n2889), .A3(n2888), .A4(n2887), 
        .ZN(n2891) );
  ND4D1BWP30P140LVT U3277 ( .A1(n2894), .A2(n2893), .A3(n2892), .A4(n2891), 
        .ZN(o_data_bus[170]) );
  AOI22D1BWP30P140LVT U3278 ( .A1(i_data_bus[75]), .A2(n3317), .B1(
        i_data_bus[651]), .B2(n3302), .ZN(n2914) );
  AOI22D1BWP30P140LVT U3279 ( .A1(i_data_bus[747]), .A2(n2659), .B1(
        i_data_bus[299]), .B2(n3322), .ZN(n2913) );
  AOI22D1BWP30P140LVT U3280 ( .A1(i_data_bus[203]), .A2(n2676), .B1(
        i_data_bus[139]), .B2(n2935), .ZN(n2912) );
  AOI22D1BWP30P140LVT U3281 ( .A1(i_data_bus[43]), .A2(n3305), .B1(
        i_data_bus[779]), .B2(n3307), .ZN(n2898) );
  AOI22D1BWP30P140LVT U3282 ( .A1(i_data_bus[907]), .A2(n3309), .B1(
        i_data_bus[363]), .B2(n3321), .ZN(n2897) );
  AOI22D1BWP30P140LVT U3283 ( .A1(i_data_bus[107]), .A2(n3308), .B1(
        i_data_bus[683]), .B2(n2653), .ZN(n2896) );
  AOI22D1BWP30P140LVT U3284 ( .A1(i_data_bus[939]), .A2(n3311), .B1(
        i_data_bus[11]), .B2(n3319), .ZN(n2895) );
  ND4D1BWP30P140LVT U3285 ( .A1(n2898), .A2(n2897), .A3(n2896), .A4(n2895), 
        .ZN(n2910) );
  AOI22D1BWP30P140LVT U3286 ( .A1(i_data_bus[875]), .A2(n113), .B1(
        i_data_bus[715]), .B2(n3310), .ZN(n2902) );
  AOI22D1BWP30P140LVT U3287 ( .A1(i_data_bus[811]), .A2(n3304), .B1(
        i_data_bus[331]), .B2(n3306), .ZN(n2900) );
  AOI22D1BWP30P140LVT U3288 ( .A1(i_data_bus[1003]), .A2(n3320), .B1(
        i_data_bus[267]), .B2(n3318), .ZN(n2899) );
  ND4D1BWP30P140LVT U3289 ( .A1(n2902), .A2(n2901), .A3(n2900), .A4(n2899), 
        .ZN(n2909) );
  INVD1BWP30P140LVT U3290 ( .I(i_data_bus[459]), .ZN(n5729) );
  MOAI22D1BWP30P140LVT U3291 ( .A1(n5729), .A2(n3246), .B1(i_data_bus[171]), 
        .B2(n2678), .ZN(n2908) );
  AOI22D1BWP30P140LVT U3292 ( .A1(i_data_bus[395]), .A2(n3), .B1(
        i_data_bus[235]), .B2(n3328), .ZN(n2906) );
  AOI22D1BWP30P140LVT U3293 ( .A1(i_data_bus[491]), .A2(n3329), .B1(
        i_data_bus[427]), .B2(n3303), .ZN(n2905) );
  AOI22D1BWP30P140LVT U3294 ( .A1(i_data_bus[619]), .A2(n3333), .B1(
        i_data_bus[587]), .B2(n3334), .ZN(n2904) );
  AOI22D1BWP30P140LVT U3295 ( .A1(i_data_bus[523]), .A2(n3331), .B1(
        i_data_bus[555]), .B2(n3332), .ZN(n2903) );
  ND4D1BWP30P140LVT U3296 ( .A1(n2906), .A2(n2905), .A3(n2904), .A4(n2903), 
        .ZN(n2907) );
  NR4D0BWP30P140LVT U3297 ( .A1(n2910), .A2(n2909), .A3(n2908), .A4(n2907), 
        .ZN(n2911) );
  ND4D1BWP30P140LVT U3298 ( .A1(n2914), .A2(n2913), .A3(n2912), .A4(n2911), 
        .ZN(o_data_bus[171]) );
  AOI22D1BWP30P140LVT U3299 ( .A1(i_data_bus[876]), .A2(n113), .B1(
        i_data_bus[332]), .B2(n3306), .ZN(n2934) );
  AOI22D1BWP30P140LVT U3300 ( .A1(i_data_bus[12]), .A2(n3319), .B1(
        i_data_bus[972]), .B2(n3301), .ZN(n2933) );
  AOI22D1BWP30P140LVT U3301 ( .A1(i_data_bus[460]), .A2(n3330), .B1(
        i_data_bus[396]), .B2(n3), .ZN(n2932) );
  AOI22D1BWP30P140LVT U3302 ( .A1(i_data_bus[908]), .A2(n3309), .B1(
        i_data_bus[108]), .B2(n3308), .ZN(n2918) );
  AOI22D1BWP30P140LVT U3303 ( .A1(i_data_bus[364]), .A2(n3321), .B1(
        i_data_bus[652]), .B2(n3302), .ZN(n2916) );
  AOI22D1BWP30P140LVT U3304 ( .A1(i_data_bus[780]), .A2(n3307), .B1(
        i_data_bus[812]), .B2(n3304), .ZN(n2915) );
  ND4D1BWP30P140LVT U3305 ( .A1(n2918), .A2(n2917), .A3(n2916), .A4(n2915), 
        .ZN(n2930) );
  AOI22D1BWP30P140LVT U3306 ( .A1(i_data_bus[44]), .A2(n3305), .B1(
        i_data_bus[1004]), .B2(n3320), .ZN(n2922) );
  AOI22D1BWP30P140LVT U3307 ( .A1(i_data_bus[940]), .A2(n3311), .B1(
        i_data_bus[300]), .B2(n3322), .ZN(n2921) );
  AOI22D1BWP30P140LVT U3308 ( .A1(i_data_bus[716]), .A2(n3310), .B1(
        i_data_bus[748]), .B2(n2659), .ZN(n2920) );
  AOI22D1BWP30P140LVT U3309 ( .A1(i_data_bus[684]), .A2(n2653), .B1(
        i_data_bus[268]), .B2(n3318), .ZN(n2919) );
  ND4D1BWP30P140LVT U3310 ( .A1(n2922), .A2(n2921), .A3(n2920), .A4(n2919), 
        .ZN(n2929) );
  INVD1BWP30P140LVT U3311 ( .I(i_data_bus[492]), .ZN(n5014) );
  INVD1BWP30P140LVT U3312 ( .I(i_data_bus[172]), .ZN(n5750) );
  OAI22D1BWP30P140LVT U3313 ( .A1(n5014), .A2(n3267), .B1(n5750), .B2(n3327), 
        .ZN(n2928) );
  AOI22D1BWP30P140LVT U3314 ( .A1(i_data_bus[204]), .A2(n2676), .B1(
        i_data_bus[236]), .B2(n3328), .ZN(n2926) );
  AOI22D1BWP30P140LVT U3315 ( .A1(i_data_bus[428]), .A2(n3303), .B1(
        i_data_bus[140]), .B2(n2935), .ZN(n2925) );
  AOI22D1BWP30P140LVT U3316 ( .A1(i_data_bus[620]), .A2(n3333), .B1(
        i_data_bus[524]), .B2(n3331), .ZN(n2924) );
  AOI22D1BWP30P140LVT U3317 ( .A1(i_data_bus[556]), .A2(n3332), .B1(
        i_data_bus[588]), .B2(n3334), .ZN(n2923) );
  ND4D1BWP30P140LVT U3318 ( .A1(n2926), .A2(n2925), .A3(n2924), .A4(n2923), 
        .ZN(n2927) );
  NR4D0BWP30P140LVT U3319 ( .A1(n2930), .A2(n2929), .A3(n2928), .A4(n2927), 
        .ZN(n2931) );
  ND4D1BWP30P140LVT U3320 ( .A1(n2934), .A2(n2933), .A3(n2932), .A4(n2931), 
        .ZN(o_data_bus[172]) );
  AOI22D1BWP30P140LVT U3321 ( .A1(i_data_bus[77]), .A2(n3317), .B1(
        i_data_bus[813]), .B2(n3304), .ZN(n2955) );
  AOI22D1BWP30P140LVT U3322 ( .A1(i_data_bus[365]), .A2(n3321), .B1(
        i_data_bus[877]), .B2(n113), .ZN(n2954) );
  AOI22D1BWP30P140LVT U3323 ( .A1(i_data_bus[141]), .A2(n2935), .B1(
        i_data_bus[461]), .B2(n3330), .ZN(n2953) );
  AOI22D1BWP30P140LVT U3324 ( .A1(i_data_bus[749]), .A2(n2659), .B1(
        i_data_bus[717]), .B2(n3310), .ZN(n2939) );
  AOI22D1BWP30P140LVT U3325 ( .A1(i_data_bus[1005]), .A2(n58), .B1(
        i_data_bus[653]), .B2(n3302), .ZN(n2938) );
  AOI22D1BWP30P140LVT U3326 ( .A1(i_data_bus[909]), .A2(n3309), .B1(
        i_data_bus[301]), .B2(n3322), .ZN(n2937) );
  AOI22D1BWP30P140LVT U3327 ( .A1(i_data_bus[973]), .A2(n3301), .B1(
        i_data_bus[109]), .B2(n3308), .ZN(n2936) );
  ND4D1BWP30P140LVT U3328 ( .A1(n2939), .A2(n2938), .A3(n2937), .A4(n2936), 
        .ZN(n2951) );
  AOI22D1BWP30P140LVT U3329 ( .A1(i_data_bus[45]), .A2(n3305), .B1(
        i_data_bus[685]), .B2(n2653), .ZN(n2942) );
  AOI22D1BWP30P140LVT U3330 ( .A1(i_data_bus[941]), .A2(n3311), .B1(
        i_data_bus[781]), .B2(n3307), .ZN(n2941) );
  AOI22D1BWP30P140LVT U3331 ( .A1(i_data_bus[13]), .A2(n3319), .B1(
        i_data_bus[333]), .B2(n3306), .ZN(n2940) );
  ND4D1BWP30P140LVT U3332 ( .A1(n2943), .A2(n2942), .A3(n2941), .A4(n2940), 
        .ZN(n2950) );
  INVD1BWP30P140LVT U3333 ( .I(i_data_bus[493]), .ZN(n5036) );
  INVD1BWP30P140LVT U3334 ( .I(i_data_bus[173]), .ZN(n5771) );
  OAI22D1BWP30P140LVT U3335 ( .A1(n5036), .A2(n3267), .B1(n5771), .B2(n3327), 
        .ZN(n2949) );
  AOI22D1BWP30P140LVT U3336 ( .A1(i_data_bus[237]), .A2(n3328), .B1(
        i_data_bus[397]), .B2(n3), .ZN(n2947) );
  AOI22D1BWP30P140LVT U3337 ( .A1(i_data_bus[429]), .A2(n3303), .B1(
        i_data_bus[205]), .B2(n2676), .ZN(n2946) );
  AOI22D1BWP30P140LVT U3338 ( .A1(i_data_bus[525]), .A2(n3331), .B1(
        i_data_bus[557]), .B2(n3332), .ZN(n2945) );
  AOI22D1BWP30P140LVT U3339 ( .A1(i_data_bus[621]), .A2(n3333), .B1(
        i_data_bus[589]), .B2(n3334), .ZN(n2944) );
  ND4D1BWP30P140LVT U3340 ( .A1(n2947), .A2(n2946), .A3(n2945), .A4(n2944), 
        .ZN(n2948) );
  NR4D0BWP30P140LVT U3341 ( .A1(n2951), .A2(n2950), .A3(n2949), .A4(n2948), 
        .ZN(n2952) );
  ND4D1BWP30P140LVT U3342 ( .A1(n2955), .A2(n2954), .A3(n2953), .A4(n2952), 
        .ZN(o_data_bus[173]) );
  AOI22D1BWP30P140LVT U3343 ( .A1(i_data_bus[110]), .A2(n3308), .B1(
        i_data_bus[686]), .B2(n2653), .ZN(n2975) );
  AOI22D1BWP30P140LVT U3344 ( .A1(i_data_bus[302]), .A2(n3322), .B1(
        i_data_bus[718]), .B2(n3310), .ZN(n2974) );
  AOI22D1BWP30P140LVT U3345 ( .A1(i_data_bus[430]), .A2(n3303), .B1(
        i_data_bus[494]), .B2(n3329), .ZN(n2973) );
  AOI22D1BWP30P140LVT U3346 ( .A1(i_data_bus[942]), .A2(n3311), .B1(
        i_data_bus[782]), .B2(n3307), .ZN(n2959) );
  AOI22D1BWP30P140LVT U3347 ( .A1(i_data_bus[910]), .A2(n3309), .B1(
        i_data_bus[878]), .B2(n113), .ZN(n2958) );
  AOI22D1BWP30P140LVT U3348 ( .A1(i_data_bus[1006]), .A2(n58), .B1(
        i_data_bus[46]), .B2(n3305), .ZN(n2956) );
  ND4D1BWP30P140LVT U3349 ( .A1(n2959), .A2(n2958), .A3(n2957), .A4(n2956), 
        .ZN(n2971) );
  AOI22D1BWP30P140LVT U3350 ( .A1(i_data_bus[974]), .A2(n3301), .B1(
        i_data_bus[270]), .B2(n3318), .ZN(n2963) );
  AOI22D1BWP30P140LVT U3351 ( .A1(i_data_bus[14]), .A2(n3319), .B1(
        i_data_bus[750]), .B2(n2659), .ZN(n2962) );
  AOI22D1BWP30P140LVT U3352 ( .A1(i_data_bus[78]), .A2(n3317), .B1(
        i_data_bus[366]), .B2(n3321), .ZN(n2961) );
  AOI22D1BWP30P140LVT U3353 ( .A1(i_data_bus[334]), .A2(n3306), .B1(
        i_data_bus[654]), .B2(n3302), .ZN(n2960) );
  ND4D1BWP30P140LVT U3354 ( .A1(n2963), .A2(n2962), .A3(n2961), .A4(n2960), 
        .ZN(n2970) );
  INVD1BWP30P140LVT U3355 ( .I(i_data_bus[398]), .ZN(n3671) );
  MOAI22D1BWP30P140LVT U3356 ( .A1(n3671), .A2(n3288), .B1(i_data_bus[462]), 
        .B2(n3330), .ZN(n2969) );
  AOI22D1BWP30P140LVT U3357 ( .A1(i_data_bus[174]), .A2(n2678), .B1(
        i_data_bus[238]), .B2(n3328), .ZN(n2967) );
  AOI22D1BWP30P140LVT U3358 ( .A1(i_data_bus[206]), .A2(n2676), .B1(
        i_data_bus[142]), .B2(n2935), .ZN(n2966) );
  AOI22D1BWP30P140LVT U3359 ( .A1(i_data_bus[590]), .A2(n3334), .B1(
        i_data_bus[526]), .B2(n3331), .ZN(n2965) );
  AOI22D1BWP30P140LVT U3360 ( .A1(i_data_bus[558]), .A2(n3332), .B1(
        i_data_bus[622]), .B2(n3333), .ZN(n2964) );
  ND4D1BWP30P140LVT U3361 ( .A1(n2967), .A2(n2966), .A3(n2965), .A4(n2964), 
        .ZN(n2968) );
  NR4D0BWP30P140LVT U3362 ( .A1(n2971), .A2(n2970), .A3(n2969), .A4(n2968), 
        .ZN(n2972) );
  ND4D1BWP30P140LVT U3363 ( .A1(n2975), .A2(n2974), .A3(n2973), .A4(n2972), 
        .ZN(o_data_bus[174]) );
  AOI22D1BWP30P140LVT U3364 ( .A1(i_data_bus[847]), .A2(n3316), .B1(
        i_data_bus[303]), .B2(n3322), .ZN(n2995) );
  AOI22D1BWP30P140LVT U3365 ( .A1(i_data_bus[111]), .A2(n3308), .B1(
        i_data_bus[335]), .B2(n3306), .ZN(n2994) );
  AOI22D1BWP30P140LVT U3366 ( .A1(i_data_bus[239]), .A2(n3328), .B1(
        i_data_bus[495]), .B2(n3329), .ZN(n2993) );
  AOI22D1BWP30P140LVT U3367 ( .A1(i_data_bus[271]), .A2(n3318), .B1(
        i_data_bus[815]), .B2(n3304), .ZN(n2979) );
  AOI22D1BWP30P140LVT U3368 ( .A1(i_data_bus[15]), .A2(n3319), .B1(
        i_data_bus[783]), .B2(n3307), .ZN(n2978) );
  AOI22D1BWP30P140LVT U3369 ( .A1(i_data_bus[911]), .A2(n3309), .B1(
        i_data_bus[879]), .B2(n113), .ZN(n2977) );
  AOI22D1BWP30P140LVT U3370 ( .A1(i_data_bus[719]), .A2(n3310), .B1(
        i_data_bus[655]), .B2(n3302), .ZN(n2976) );
  ND4D1BWP30P140LVT U3371 ( .A1(n2979), .A2(n2978), .A3(n2977), .A4(n2976), 
        .ZN(n2991) );
  AOI22D1BWP30P140LVT U3372 ( .A1(i_data_bus[975]), .A2(n3301), .B1(
        i_data_bus[367]), .B2(n3321), .ZN(n2983) );
  AOI22D1BWP30P140LVT U3373 ( .A1(i_data_bus[943]), .A2(n3311), .B1(
        i_data_bus[687]), .B2(n2653), .ZN(n2982) );
  AOI22D1BWP30P140LVT U3374 ( .A1(i_data_bus[1007]), .A2(n59), .B1(
        i_data_bus[751]), .B2(n2659), .ZN(n2981) );
  AOI22D1BWP30P140LVT U3375 ( .A1(i_data_bus[79]), .A2(n3317), .B1(
        i_data_bus[47]), .B2(n3305), .ZN(n2980) );
  ND4D1BWP30P140LVT U3376 ( .A1(n2983), .A2(n2982), .A3(n2981), .A4(n2980), 
        .ZN(n2990) );
  INVD1BWP30P140LVT U3377 ( .I(i_data_bus[463]), .ZN(n3688) );
  MOAI22D1BWP30P140LVT U3378 ( .A1(n3688), .A2(n3246), .B1(i_data_bus[143]), 
        .B2(n2935), .ZN(n2989) );
  AOI22D1BWP30P140LVT U3379 ( .A1(i_data_bus[431]), .A2(n3303), .B1(
        i_data_bus[399]), .B2(n3), .ZN(n2987) );
  AOI22D1BWP30P140LVT U3380 ( .A1(i_data_bus[207]), .A2(n2676), .B1(
        i_data_bus[175]), .B2(n2678), .ZN(n2986) );
  AOI22D1BWP30P140LVT U3381 ( .A1(i_data_bus[559]), .A2(n3332), .B1(
        i_data_bus[527]), .B2(n3331), .ZN(n2985) );
  AOI22D1BWP30P140LVT U3382 ( .A1(i_data_bus[591]), .A2(n3334), .B1(
        i_data_bus[623]), .B2(n3333), .ZN(n2984) );
  ND4D1BWP30P140LVT U3383 ( .A1(n2987), .A2(n2986), .A3(n2985), .A4(n2984), 
        .ZN(n2988) );
  NR4D0BWP30P140LVT U3384 ( .A1(n2991), .A2(n2990), .A3(n2989), .A4(n2988), 
        .ZN(n2992) );
  ND4D1BWP30P140LVT U3385 ( .A1(n2995), .A2(n2994), .A3(n2993), .A4(n2992), 
        .ZN(o_data_bus[175]) );
  AOI22D1BWP30P140LVT U3386 ( .A1(i_data_bus[112]), .A2(n3308), .B1(
        i_data_bus[752]), .B2(n2659), .ZN(n3015) );
  AOI22D1BWP30P140LVT U3387 ( .A1(i_data_bus[16]), .A2(n3319), .B1(
        i_data_bus[1008]), .B2(n58), .ZN(n3014) );
  AOI22D1BWP30P140LVT U3388 ( .A1(i_data_bus[432]), .A2(n3303), .B1(
        i_data_bus[240]), .B2(n3328), .ZN(n3013) );
  AOI22D1BWP30P140LVT U3389 ( .A1(i_data_bus[944]), .A2(n3311), .B1(
        i_data_bus[272]), .B2(n3318), .ZN(n2999) );
  AOI22D1BWP30P140LVT U3390 ( .A1(i_data_bus[80]), .A2(n3317), .B1(
        i_data_bus[688]), .B2(n2653), .ZN(n2998) );
  AOI22D1BWP30P140LVT U3391 ( .A1(i_data_bus[656]), .A2(n3302), .B1(
        i_data_bus[816]), .B2(n3304), .ZN(n2997) );
  AOI22D1BWP30P140LVT U3392 ( .A1(i_data_bus[976]), .A2(n3301), .B1(
        i_data_bus[304]), .B2(n3322), .ZN(n2996) );
  ND4D1BWP30P140LVT U3393 ( .A1(n2999), .A2(n2998), .A3(n2997), .A4(n2996), 
        .ZN(n3011) );
  AOI22D1BWP30P140LVT U3394 ( .A1(i_data_bus[336]), .A2(n3306), .B1(
        i_data_bus[880]), .B2(n113), .ZN(n3003) );
  AOI22D1BWP30P140LVT U3395 ( .A1(i_data_bus[912]), .A2(n3309), .B1(
        i_data_bus[368]), .B2(n3321), .ZN(n3002) );
  AOI22D1BWP30P140LVT U3396 ( .A1(i_data_bus[48]), .A2(n3305), .B1(
        i_data_bus[720]), .B2(n3310), .ZN(n3000) );
  ND4D1BWP30P140LVT U3397 ( .A1(n3003), .A2(n3002), .A3(n3001), .A4(n3000), 
        .ZN(n3010) );
  INVD1BWP30P140LVT U3398 ( .I(i_data_bus[496]), .ZN(n3709) );
  MOAI22D1BWP30P140LVT U3399 ( .A1(n3709), .A2(n3267), .B1(i_data_bus[176]), 
        .B2(n2678), .ZN(n3009) );
  AOI22D1BWP30P140LVT U3400 ( .A1(i_data_bus[144]), .A2(n2935), .B1(
        i_data_bus[400]), .B2(n3), .ZN(n3007) );
  AOI22D1BWP30P140LVT U3401 ( .A1(i_data_bus[208]), .A2(n2676), .B1(
        i_data_bus[464]), .B2(n3330), .ZN(n3006) );
  AOI22D1BWP30P140LVT U3402 ( .A1(i_data_bus[560]), .A2(n3332), .B1(
        i_data_bus[528]), .B2(n3331), .ZN(n3005) );
  AOI22D1BWP30P140LVT U3403 ( .A1(i_data_bus[624]), .A2(n3333), .B1(
        i_data_bus[592]), .B2(n3334), .ZN(n3004) );
  ND4D1BWP30P140LVT U3404 ( .A1(n3007), .A2(n3006), .A3(n3005), .A4(n3004), 
        .ZN(n3008) );
  NR4D0BWP30P140LVT U3405 ( .A1(n3011), .A2(n3010), .A3(n3009), .A4(n3008), 
        .ZN(n3012) );
  ND4D1BWP30P140LVT U3406 ( .A1(n3015), .A2(n3014), .A3(n3013), .A4(n3012), 
        .ZN(o_data_bus[176]) );
  AOI22D1BWP30P140LVT U3407 ( .A1(i_data_bus[337]), .A2(n3306), .B1(
        i_data_bus[273]), .B2(n3318), .ZN(n3035) );
  AOI22D1BWP30P140LVT U3408 ( .A1(i_data_bus[945]), .A2(n3311), .B1(
        i_data_bus[113]), .B2(n3308), .ZN(n3034) );
  AOI22D1BWP30P140LVT U3409 ( .A1(i_data_bus[433]), .A2(n3303), .B1(
        i_data_bus[497]), .B2(n3329), .ZN(n3033) );
  AOI22D1BWP30P140LVT U3410 ( .A1(i_data_bus[209]), .A2(n2676), .B1(
        i_data_bus[177]), .B2(n2678), .ZN(n3031) );
  AOI22D1BWP30P140LVT U3411 ( .A1(i_data_bus[1009]), .A2(n3320), .B1(
        i_data_bus[817]), .B2(n3304), .ZN(n3018) );
  AOI22D1BWP30P140LVT U3412 ( .A1(i_data_bus[17]), .A2(n3319), .B1(
        i_data_bus[305]), .B2(n3322), .ZN(n3017) );
  AOI22D1BWP30P140LVT U3413 ( .A1(i_data_bus[689]), .A2(n2653), .B1(
        i_data_bus[753]), .B2(n2659), .ZN(n3016) );
  ND4D1BWP30P140LVT U3414 ( .A1(n3019), .A2(n3018), .A3(n3017), .A4(n3016), 
        .ZN(n3030) );
  AOI22D1BWP30P140LVT U3415 ( .A1(i_data_bus[977]), .A2(n3301), .B1(
        i_data_bus[721]), .B2(n3310), .ZN(n3023) );
  AOI22D1BWP30P140LVT U3416 ( .A1(i_data_bus[81]), .A2(n3317), .B1(
        i_data_bus[657]), .B2(n3302), .ZN(n3022) );
  AOI22D1BWP30P140LVT U3417 ( .A1(i_data_bus[913]), .A2(n3309), .B1(
        i_data_bus[881]), .B2(n113), .ZN(n3021) );
  AOI22D1BWP30P140LVT U3418 ( .A1(i_data_bus[785]), .A2(n3307), .B1(
        i_data_bus[369]), .B2(n3321), .ZN(n3020) );
  ND4D1BWP30P140LVT U3419 ( .A1(n3023), .A2(n3022), .A3(n3021), .A4(n3020), 
        .ZN(n3029) );
  AOI22D1BWP30P140LVT U3420 ( .A1(i_data_bus[145]), .A2(n2935), .B1(
        i_data_bus[241]), .B2(n3328), .ZN(n3027) );
  AOI22D1BWP30P140LVT U3421 ( .A1(i_data_bus[401]), .A2(n3), .B1(
        i_data_bus[465]), .B2(n3330), .ZN(n3026) );
  AOI22D1BWP30P140LVT U3422 ( .A1(i_data_bus[593]), .A2(n3334), .B1(
        i_data_bus[561]), .B2(n3332), .ZN(n3025) );
  AOI22D1BWP30P140LVT U3423 ( .A1(i_data_bus[625]), .A2(n3333), .B1(
        i_data_bus[529]), .B2(n3331), .ZN(n3024) );
  ND4D1BWP30P140LVT U3424 ( .A1(n3027), .A2(n3026), .A3(n3025), .A4(n3024), 
        .ZN(n3028) );
  INR4D0BWP30P140LVT U3425 ( .A1(n3031), .B1(n3030), .B2(n3029), .B3(n3028), 
        .ZN(n3032) );
  ND4D1BWP30P140LVT U3426 ( .A1(n3035), .A2(n3034), .A3(n3033), .A4(n3032), 
        .ZN(o_data_bus[177]) );
  AOI22D1BWP30P140LVT U3427 ( .A1(i_data_bus[1010]), .A2(n3320), .B1(
        i_data_bus[722]), .B2(n3310), .ZN(n3056) );
  AOI22D1BWP30P140LVT U3428 ( .A1(i_data_bus[818]), .A2(n3304), .B1(
        i_data_bus[338]), .B2(n3306), .ZN(n3055) );
  AOI22D1BWP30P140LVT U3429 ( .A1(i_data_bus[210]), .A2(n2676), .B1(
        i_data_bus[498]), .B2(n3329), .ZN(n3054) );
  AOI22D1BWP30P140LVT U3430 ( .A1(i_data_bus[946]), .A2(n3311), .B1(
        i_data_bus[370]), .B2(n3321), .ZN(n3039) );
  AOI22D1BWP30P140LVT U3431 ( .A1(i_data_bus[50]), .A2(n3305), .B1(
        i_data_bus[914]), .B2(n3309), .ZN(n3038) );
  AOI22D1BWP30P140LVT U3432 ( .A1(i_data_bus[882]), .A2(n113), .B1(
        i_data_bus[658]), .B2(n3302), .ZN(n3037) );
  AOI22D1BWP30P140LVT U3433 ( .A1(i_data_bus[274]), .A2(n3318), .B1(
        i_data_bus[754]), .B2(n2659), .ZN(n3036) );
  ND4D1BWP30P140LVT U3434 ( .A1(n3039), .A2(n3038), .A3(n3037), .A4(n3036), 
        .ZN(n3052) );
  AOI22D1BWP30P140LVT U3435 ( .A1(i_data_bus[978]), .A2(n3301), .B1(
        i_data_bus[690]), .B2(n2653), .ZN(n3042) );
  AOI22D1BWP30P140LVT U3436 ( .A1(i_data_bus[114]), .A2(n3308), .B1(
        i_data_bus[82]), .B2(n3317), .ZN(n3041) );
  AOI22D1BWP30P140LVT U3437 ( .A1(i_data_bus[18]), .A2(n3319), .B1(
        i_data_bus[850]), .B2(n3316), .ZN(n3040) );
  INVD1BWP30P140LVT U3438 ( .I(i_data_bus[146]), .ZN(n5877) );
  MOAI22D1BWP30P140LVT U3439 ( .A1(n5877), .A2(n3044), .B1(i_data_bus[178]), 
        .B2(n2678), .ZN(n3050) );
  AOI22D1BWP30P140LVT U3440 ( .A1(i_data_bus[402]), .A2(n3), .B1(
        i_data_bus[242]), .B2(n3328), .ZN(n3048) );
  AOI22D1BWP30P140LVT U3441 ( .A1(i_data_bus[466]), .A2(n3330), .B1(
        i_data_bus[434]), .B2(n3303), .ZN(n3047) );
  AOI22D1BWP30P140LVT U3442 ( .A1(i_data_bus[594]), .A2(n3334), .B1(
        i_data_bus[530]), .B2(n3331), .ZN(n3046) );
  AOI22D1BWP30P140LVT U3443 ( .A1(i_data_bus[626]), .A2(n3333), .B1(
        i_data_bus[562]), .B2(n3332), .ZN(n3045) );
  ND4D1BWP30P140LVT U3444 ( .A1(n3048), .A2(n3047), .A3(n3046), .A4(n3045), 
        .ZN(n3049) );
  NR4D0BWP30P140LVT U3445 ( .A1(n3051), .A2(n3052), .A3(n3050), .A4(n3049), 
        .ZN(n3053) );
  AOI22D1BWP30P140LVT U3446 ( .A1(i_data_bus[339]), .A2(n3306), .B1(
        i_data_bus[851]), .B2(n3316), .ZN(n3076) );
  AOI22D1BWP30P140LVT U3447 ( .A1(i_data_bus[83]), .A2(n3317), .B1(
        i_data_bus[659]), .B2(n3302), .ZN(n3075) );
  AOI22D1BWP30P140LVT U3448 ( .A1(i_data_bus[211]), .A2(n2676), .B1(
        i_data_bus[467]), .B2(n3330), .ZN(n3074) );
  AOI22D1BWP30P140LVT U3449 ( .A1(i_data_bus[179]), .A2(n2678), .B1(
        i_data_bus[147]), .B2(n2935), .ZN(n3072) );
  AOI22D1BWP30P140LVT U3450 ( .A1(i_data_bus[115]), .A2(n3308), .B1(
        i_data_bus[275]), .B2(n3318), .ZN(n3060) );
  AOI22D1BWP30P140LVT U3451 ( .A1(i_data_bus[307]), .A2(n3322), .B1(
        i_data_bus[819]), .B2(n3304), .ZN(n3059) );
  AOI22D1BWP30P140LVT U3452 ( .A1(i_data_bus[947]), .A2(n3311), .B1(
        i_data_bus[787]), .B2(n3307), .ZN(n3058) );
  AOI22D1BWP30P140LVT U3453 ( .A1(i_data_bus[979]), .A2(n3301), .B1(
        i_data_bus[883]), .B2(n113), .ZN(n3057) );
  ND4D1BWP30P140LVT U3454 ( .A1(n3060), .A2(n3059), .A3(n3058), .A4(n3057), 
        .ZN(n3071) );
  AOI22D1BWP30P140LVT U3455 ( .A1(i_data_bus[19]), .A2(n3319), .B1(
        i_data_bus[691]), .B2(n2653), .ZN(n3064) );
  AOI22D1BWP30P140LVT U3456 ( .A1(i_data_bus[915]), .A2(n3309), .B1(
        i_data_bus[755]), .B2(n2659), .ZN(n3063) );
  AOI22D1BWP30P140LVT U3457 ( .A1(i_data_bus[51]), .A2(n3305), .B1(
        i_data_bus[723]), .B2(n3310), .ZN(n3062) );
  AOI22D1BWP30P140LVT U3458 ( .A1(i_data_bus[1011]), .A2(n3320), .B1(
        i_data_bus[371]), .B2(n3321), .ZN(n3061) );
  ND4D1BWP30P140LVT U3459 ( .A1(n3064), .A2(n3063), .A3(n3062), .A4(n3061), 
        .ZN(n3070) );
  AOI22D1BWP30P140LVT U3460 ( .A1(i_data_bus[243]), .A2(n3328), .B1(
        i_data_bus[435]), .B2(n3303), .ZN(n3068) );
  AOI22D1BWP30P140LVT U3461 ( .A1(i_data_bus[403]), .A2(n3), .B1(
        i_data_bus[499]), .B2(n3329), .ZN(n3067) );
  AOI22D1BWP30P140LVT U3462 ( .A1(i_data_bus[531]), .A2(n3331), .B1(
        i_data_bus[595]), .B2(n3334), .ZN(n3066) );
  AOI22D1BWP30P140LVT U3463 ( .A1(i_data_bus[563]), .A2(n3332), .B1(
        i_data_bus[627]), .B2(n3333), .ZN(n3065) );
  ND4D1BWP30P140LVT U3464 ( .A1(n3068), .A2(n3067), .A3(n3066), .A4(n3065), 
        .ZN(n3069) );
  INR4D0BWP30P140LVT U3465 ( .A1(n3072), .B1(n3071), .B2(n3070), .B3(n3069), 
        .ZN(n3073) );
  ND4D1BWP30P140LVT U3466 ( .A1(n3076), .A2(n3075), .A3(n3074), .A4(n3073), 
        .ZN(o_data_bus[179]) );
  AOI22D1BWP30P140LVT U3467 ( .A1(i_data_bus[948]), .A2(n7), .B1(
        i_data_bus[84]), .B2(n3317), .ZN(n3096) );
  AOI22D1BWP30P140LVT U3468 ( .A1(i_data_bus[1012]), .A2(n59), .B1(
        i_data_bus[884]), .B2(n113), .ZN(n3095) );
  AOI22D1BWP30P140LVT U3469 ( .A1(i_data_bus[244]), .A2(n3328), .B1(
        i_data_bus[436]), .B2(n3303), .ZN(n3094) );
  AOI22D1BWP30P140LVT U3470 ( .A1(i_data_bus[276]), .A2(n3318), .B1(
        i_data_bus[660]), .B2(n3302), .ZN(n3080) );
  AOI22D1BWP30P140LVT U3471 ( .A1(i_data_bus[52]), .A2(n3305), .B1(
        i_data_bus[692]), .B2(n2653), .ZN(n3079) );
  AOI22D1BWP30P140LVT U3472 ( .A1(i_data_bus[980]), .A2(n3301), .B1(
        i_data_bus[116]), .B2(n3308), .ZN(n3078) );
  AOI22D1BWP30P140LVT U3473 ( .A1(i_data_bus[916]), .A2(n3309), .B1(
        i_data_bus[724]), .B2(n3310), .ZN(n3077) );
  ND4D1BWP30P140LVT U3474 ( .A1(n3080), .A2(n3079), .A3(n3078), .A4(n3077), 
        .ZN(n3092) );
  AOI22D1BWP30P140LVT U3475 ( .A1(i_data_bus[340]), .A2(n3306), .B1(
        i_data_bus[820]), .B2(n3304), .ZN(n3084) );
  AOI22D1BWP30P140LVT U3476 ( .A1(i_data_bus[20]), .A2(n3319), .B1(
        i_data_bus[756]), .B2(n2659), .ZN(n3083) );
  AOI22D1BWP30P140LVT U3477 ( .A1(i_data_bus[852]), .A2(n3316), .B1(
        i_data_bus[372]), .B2(n3321), .ZN(n3082) );
  AOI22D1BWP30P140LVT U3478 ( .A1(i_data_bus[788]), .A2(n3307), .B1(
        i_data_bus[308]), .B2(n3322), .ZN(n3081) );
  ND4D1BWP30P140LVT U3479 ( .A1(n3082), .A2(n3083), .A3(n3084), .A4(n3081), 
        .ZN(n3091) );
  INVD1BWP30P140LVT U3480 ( .I(i_data_bus[468]), .ZN(n3790) );
  MOAI22D1BWP30P140LVT U3481 ( .A1(n3790), .A2(n3246), .B1(i_data_bus[212]), 
        .B2(n2676), .ZN(n3090) );
  AOI22D1BWP30P140LVT U3482 ( .A1(i_data_bus[404]), .A2(n3), .B1(
        i_data_bus[148]), .B2(n2935), .ZN(n3088) );
  AOI22D1BWP30P140LVT U3483 ( .A1(i_data_bus[180]), .A2(n2678), .B1(
        i_data_bus[500]), .B2(n3329), .ZN(n3087) );
  AOI22D1BWP30P140LVT U3484 ( .A1(i_data_bus[532]), .A2(n3331), .B1(
        i_data_bus[628]), .B2(n3333), .ZN(n3086) );
  AOI22D1BWP30P140LVT U3485 ( .A1(i_data_bus[596]), .A2(n3334), .B1(
        i_data_bus[564]), .B2(n3332), .ZN(n3085) );
  ND4D1BWP30P140LVT U3486 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), 
        .ZN(n3089) );
  NR4D0BWP30P140LVT U3487 ( .A1(n3092), .A2(n3091), .A3(n3090), .A4(n3089), 
        .ZN(n3093) );
  ND4D1BWP30P140LVT U3488 ( .A1(n3096), .A2(n3095), .A3(n3094), .A4(n3093), 
        .ZN(o_data_bus[180]) );
  AOI22D1BWP30P140LVT U3489 ( .A1(i_data_bus[981]), .A2(n3301), .B1(
        i_data_bus[885]), .B2(n113), .ZN(n3116) );
  AOI22D1BWP30P140LVT U3490 ( .A1(i_data_bus[85]), .A2(n3317), .B1(
        i_data_bus[1013]), .B2(n59), .ZN(n3115) );
  AOI22D1BWP30P140LVT U3491 ( .A1(i_data_bus[181]), .A2(n2678), .B1(
        i_data_bus[469]), .B2(n3330), .ZN(n3114) );
  AOI22D1BWP30P140LVT U3492 ( .A1(i_data_bus[341]), .A2(n3306), .B1(
        i_data_bus[725]), .B2(n3310), .ZN(n3100) );
  AOI22D1BWP30P140LVT U3493 ( .A1(i_data_bus[21]), .A2(n3319), .B1(
        i_data_bus[661]), .B2(n3302), .ZN(n3099) );
  AOI22D1BWP30P140LVT U3494 ( .A1(i_data_bus[949]), .A2(n3311), .B1(
        i_data_bus[693]), .B2(n2653), .ZN(n3098) );
  AOI22D1BWP30P140LVT U3495 ( .A1(i_data_bus[53]), .A2(n3305), .B1(
        i_data_bus[117]), .B2(n3308), .ZN(n3097) );
  ND4D1BWP30P140LVT U3496 ( .A1(n3100), .A2(n3099), .A3(n3098), .A4(n3097), 
        .ZN(n3112) );
  AOI22D1BWP30P140LVT U3497 ( .A1(i_data_bus[917]), .A2(n3309), .B1(
        i_data_bus[789]), .B2(n3307), .ZN(n3104) );
  AOI22D1BWP30P140LVT U3498 ( .A1(i_data_bus[277]), .A2(n3318), .B1(
        i_data_bus[373]), .B2(n3321), .ZN(n3103) );
  AOI22D1BWP30P140LVT U3499 ( .A1(i_data_bus[757]), .A2(n2659), .B1(
        i_data_bus[821]), .B2(n3304), .ZN(n3102) );
  AOI22D1BWP30P140LVT U3500 ( .A1(i_data_bus[853]), .A2(n3316), .B1(
        i_data_bus[309]), .B2(n3322), .ZN(n3101) );
  ND4D1BWP30P140LVT U3501 ( .A1(n3101), .A2(n3103), .A3(n3102), .A4(n3104), 
        .ZN(n3111) );
  INVD1BWP30P140LVT U3502 ( .I(i_data_bus[405]), .ZN(n3811) );
  MOAI22D1BWP30P140LVT U3503 ( .A1(n3811), .A2(n3288), .B1(i_data_bus[149]), 
        .B2(n2935), .ZN(n3110) );
  AOI22D1BWP30P140LVT U3504 ( .A1(i_data_bus[437]), .A2(n3303), .B1(
        i_data_bus[245]), .B2(n3328), .ZN(n3108) );
  AOI22D1BWP30P140LVT U3505 ( .A1(i_data_bus[501]), .A2(n3329), .B1(
        i_data_bus[213]), .B2(n2676), .ZN(n3107) );
  AOI22D1BWP30P140LVT U3506 ( .A1(i_data_bus[597]), .A2(n3334), .B1(
        i_data_bus[533]), .B2(n3331), .ZN(n3106) );
  AOI22D1BWP30P140LVT U3507 ( .A1(i_data_bus[629]), .A2(n3333), .B1(
        i_data_bus[565]), .B2(n3332), .ZN(n3105) );
  ND4D1BWP30P140LVT U3508 ( .A1(n3108), .A2(n3107), .A3(n3106), .A4(n3105), 
        .ZN(n3109) );
  NR4D0BWP30P140LVT U3509 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), 
        .ZN(n3113) );
  ND4D1BWP30P140LVT U3510 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), 
        .ZN(o_data_bus[181]) );
  AOI22D1BWP30P140LVT U3511 ( .A1(i_data_bus[1014]), .A2(n58), .B1(
        i_data_bus[918]), .B2(n3309), .ZN(n3137) );
  AOI22D1BWP30P140LVT U3512 ( .A1(i_data_bus[86]), .A2(n3317), .B1(
        i_data_bus[726]), .B2(n3310), .ZN(n3136) );
  AOI22D1BWP30P140LVT U3513 ( .A1(i_data_bus[246]), .A2(n3328), .B1(
        i_data_bus[502]), .B2(n3329), .ZN(n3135) );
  AOI22D1BWP30P140LVT U3514 ( .A1(i_data_bus[982]), .A2(n3301), .B1(
        i_data_bus[662]), .B2(n3302), .ZN(n3120) );
  AOI22D1BWP30P140LVT U3515 ( .A1(i_data_bus[118]), .A2(n3308), .B1(
        i_data_bus[310]), .B2(n3322), .ZN(n3119) );
  AOI22D1BWP30P140LVT U3516 ( .A1(i_data_bus[886]), .A2(n113), .B1(
        i_data_bus[342]), .B2(n3306), .ZN(n3118) );
  AOI22D1BWP30P140LVT U3517 ( .A1(i_data_bus[22]), .A2(n3319), .B1(
        i_data_bus[822]), .B2(n3304), .ZN(n3117) );
  ND4D1BWP30P140LVT U3518 ( .A1(n3120), .A2(n3119), .A3(n3118), .A4(n3117), 
        .ZN(n3133) );
  AOI22D1BWP30P140LVT U3519 ( .A1(i_data_bus[374]), .A2(n3321), .B1(
        i_data_bus[278]), .B2(n3318), .ZN(n3124) );
  AOI22D1BWP30P140LVT U3520 ( .A1(i_data_bus[950]), .A2(n3311), .B1(
        i_data_bus[758]), .B2(n2659), .ZN(n3122) );
  AOI22D1BWP30P140LVT U3521 ( .A1(i_data_bus[54]), .A2(n3305), .B1(
        i_data_bus[790]), .B2(n3307), .ZN(n3121) );
  ND4D1BWP30P140LVT U3522 ( .A1(n3124), .A2(n3123), .A3(n3122), .A4(n3121), 
        .ZN(n3132) );
  INVD1BWP30P140LVT U3523 ( .I(i_data_bus[470]), .ZN(n5222) );
  INVD1BWP30P140LVT U3524 ( .I(i_data_bus[214]), .ZN(n5964) );
  OAI22D1BWP30P140LVT U3525 ( .A1(n5222), .A2(n3246), .B1(n5964), .B2(n3125), 
        .ZN(n3131) );
  AOI22D1BWP30P140LVT U3526 ( .A1(i_data_bus[182]), .A2(n2678), .B1(
        i_data_bus[150]), .B2(n2935), .ZN(n3129) );
  AOI22D1BWP30P140LVT U3527 ( .A1(i_data_bus[438]), .A2(n3303), .B1(
        i_data_bus[406]), .B2(n3), .ZN(n3128) );
  AOI22D1BWP30P140LVT U3528 ( .A1(i_data_bus[534]), .A2(n3331), .B1(
        i_data_bus[630]), .B2(n3333), .ZN(n3127) );
  AOI22D1BWP30P140LVT U3529 ( .A1(i_data_bus[566]), .A2(n3332), .B1(
        i_data_bus[598]), .B2(n3334), .ZN(n3126) );
  ND4D1BWP30P140LVT U3530 ( .A1(n3129), .A2(n3128), .A3(n3127), .A4(n3126), 
        .ZN(n3130) );
  NR4D0BWP30P140LVT U3531 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), 
        .ZN(n3134) );
  ND4D1BWP30P140LVT U3532 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), 
        .ZN(o_data_bus[182]) );
  AOI22D1BWP30P140LVT U3533 ( .A1(i_data_bus[1015]), .A2(n59), .B1(
        i_data_bus[87]), .B2(n3317), .ZN(n3157) );
  AOI22D1BWP30P140LVT U3534 ( .A1(i_data_bus[919]), .A2(n3309), .B1(
        i_data_bus[279]), .B2(n3318), .ZN(n3156) );
  AOI22D1BWP30P140LVT U3535 ( .A1(i_data_bus[247]), .A2(n3328), .B1(
        i_data_bus[439]), .B2(n3303), .ZN(n3155) );
  AOI22D1BWP30P140LVT U3536 ( .A1(i_data_bus[695]), .A2(n2653), .B1(
        i_data_bus[663]), .B2(n3302), .ZN(n3141) );
  AOI22D1BWP30P140LVT U3537 ( .A1(i_data_bus[311]), .A2(n3322), .B1(
        i_data_bus[375]), .B2(n3321), .ZN(n3140) );
  AOI22D1BWP30P140LVT U3538 ( .A1(i_data_bus[983]), .A2(n3301), .B1(
        i_data_bus[823]), .B2(n3304), .ZN(n3139) );
  AOI22D1BWP30P140LVT U3539 ( .A1(i_data_bus[55]), .A2(n3305), .B1(
        i_data_bus[887]), .B2(n113), .ZN(n3138) );
  ND4D1BWP30P140LVT U3540 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), 
        .ZN(n3153) );
  AOI22D1BWP30P140LVT U3541 ( .A1(i_data_bus[23]), .A2(n3319), .B1(
        i_data_bus[791]), .B2(n3307), .ZN(n3145) );
  AOI22D1BWP30P140LVT U3542 ( .A1(i_data_bus[119]), .A2(n3308), .B1(
        i_data_bus[727]), .B2(n3310), .ZN(n3144) );
  AOI22D1BWP30P140LVT U3543 ( .A1(i_data_bus[951]), .A2(n3311), .B1(
        i_data_bus[343]), .B2(n3306), .ZN(n3143) );
  ND4D1BWP30P140LVT U3544 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), 
        .ZN(n3152) );
  INVD1BWP30P140LVT U3545 ( .I(i_data_bus[471]), .ZN(n5243) );
  MOAI22D1BWP30P140LVT U3546 ( .A1(n5243), .A2(n3246), .B1(i_data_bus[183]), 
        .B2(n2678), .ZN(n3151) );
  AOI22D1BWP30P140LVT U3547 ( .A1(i_data_bus[151]), .A2(n2935), .B1(
        i_data_bus[407]), .B2(n3), .ZN(n3149) );
  AOI22D1BWP30P140LVT U3548 ( .A1(i_data_bus[215]), .A2(n2676), .B1(
        i_data_bus[503]), .B2(n3329), .ZN(n3148) );
  AOI22D1BWP30P140LVT U3549 ( .A1(i_data_bus[631]), .A2(n3333), .B1(
        i_data_bus[567]), .B2(n3332), .ZN(n3147) );
  AOI22D1BWP30P140LVT U3550 ( .A1(i_data_bus[599]), .A2(n3334), .B1(
        i_data_bus[535]), .B2(n3331), .ZN(n3146) );
  ND4D1BWP30P140LVT U3551 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), 
        .ZN(n3150) );
  NR4D0BWP30P140LVT U3552 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), 
        .ZN(n3154) );
  ND4D1BWP30P140LVT U3553 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), 
        .ZN(o_data_bus[183]) );
  AOI22D1BWP30P140LVT U3554 ( .A1(i_data_bus[984]), .A2(n3301), .B1(
        i_data_bus[120]), .B2(n3308), .ZN(n3177) );
  AOI22D1BWP30P140LVT U3555 ( .A1(i_data_bus[280]), .A2(n3318), .B1(
        i_data_bus[792]), .B2(n3307), .ZN(n3176) );
  AOI22D1BWP30P140LVT U3556 ( .A1(i_data_bus[248]), .A2(n3328), .B1(
        i_data_bus[472]), .B2(n3330), .ZN(n3175) );
  AOI22D1BWP30P140LVT U3557 ( .A1(i_data_bus[696]), .A2(n2653), .B1(
        i_data_bus[824]), .B2(n3304), .ZN(n3161) );
  AOI22D1BWP30P140LVT U3558 ( .A1(i_data_bus[24]), .A2(n3319), .B1(
        i_data_bus[760]), .B2(n2659), .ZN(n3160) );
  AOI22D1BWP30P140LVT U3559 ( .A1(i_data_bus[344]), .A2(n3306), .B1(
        i_data_bus[312]), .B2(n3322), .ZN(n3159) );
  ND4D1BWP30P140LVT U3560 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), 
        .ZN(n3173) );
  AOI22D1BWP30P140LVT U3561 ( .A1(i_data_bus[376]), .A2(n3321), .B1(
        i_data_bus[888]), .B2(n113), .ZN(n3165) );
  AOI22D1BWP30P140LVT U3562 ( .A1(i_data_bus[88]), .A2(n3317), .B1(
        i_data_bus[952]), .B2(n3311), .ZN(n3164) );
  AOI22D1BWP30P140LVT U3563 ( .A1(i_data_bus[56]), .A2(n3305), .B1(
        i_data_bus[728]), .B2(n3310), .ZN(n3163) );
  AOI22D1BWP30P140LVT U3564 ( .A1(i_data_bus[920]), .A2(n3309), .B1(
        i_data_bus[664]), .B2(n3302), .ZN(n3162) );
  ND4D1BWP30P140LVT U3565 ( .A1(n3165), .A2(n3164), .A3(n3163), .A4(n3162), 
        .ZN(n3172) );
  INVD1BWP30P140LVT U3566 ( .I(i_data_bus[504]), .ZN(n3877) );
  MOAI22D1BWP30P140LVT U3567 ( .A1(n3877), .A2(n3267), .B1(i_data_bus[408]), 
        .B2(n3), .ZN(n3171) );
  AOI22D1BWP30P140LVT U3568 ( .A1(i_data_bus[152]), .A2(n2935), .B1(
        i_data_bus[216]), .B2(n2676), .ZN(n3169) );
  AOI22D1BWP30P140LVT U3569 ( .A1(i_data_bus[440]), .A2(n3303), .B1(
        i_data_bus[184]), .B2(n2678), .ZN(n3168) );
  AOI22D1BWP30P140LVT U3570 ( .A1(i_data_bus[600]), .A2(n3334), .B1(
        i_data_bus[536]), .B2(n3331), .ZN(n3167) );
  AOI22D1BWP30P140LVT U3571 ( .A1(i_data_bus[632]), .A2(n3333), .B1(
        i_data_bus[568]), .B2(n3332), .ZN(n3166) );
  ND4D1BWP30P140LVT U3572 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), 
        .ZN(n3170) );
  NR4D0BWP30P140LVT U3573 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), 
        .ZN(n3174) );
  ND4D1BWP30P140LVT U3574 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), 
        .ZN(o_data_bus[184]) );
  AOI22D1BWP30P140LVT U3575 ( .A1(i_data_bus[953]), .A2(n7), .B1(
        i_data_bus[729]), .B2(n3310), .ZN(n3197) );
  AOI22D1BWP30P140LVT U3576 ( .A1(i_data_bus[121]), .A2(n3308), .B1(
        i_data_bus[889]), .B2(n113), .ZN(n3196) );
  AOI22D1BWP30P140LVT U3577 ( .A1(i_data_bus[153]), .A2(n2935), .B1(
        i_data_bus[217]), .B2(n2676), .ZN(n3195) );
  AOI22D1BWP30P140LVT U3578 ( .A1(i_data_bus[665]), .A2(n3302), .B1(
        i_data_bus[377]), .B2(n3321), .ZN(n3181) );
  AOI22D1BWP30P140LVT U3579 ( .A1(i_data_bus[825]), .A2(n3304), .B1(
        i_data_bus[697]), .B2(n2653), .ZN(n3180) );
  AOI22D1BWP30P140LVT U3580 ( .A1(i_data_bus[921]), .A2(n3309), .B1(
        i_data_bus[793]), .B2(n3307), .ZN(n3178) );
  ND4D1BWP30P140LVT U3581 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), 
        .ZN(n3193) );
  AOI22D1BWP30P140LVT U3582 ( .A1(i_data_bus[1017]), .A2(n59), .B1(
        i_data_bus[985]), .B2(n3301), .ZN(n3185) );
  AOI22D1BWP30P140LVT U3583 ( .A1(i_data_bus[89]), .A2(n3317), .B1(
        i_data_bus[281]), .B2(n3318), .ZN(n3184) );
  AOI22D1BWP30P140LVT U3584 ( .A1(i_data_bus[25]), .A2(n3319), .B1(
        i_data_bus[345]), .B2(n3306), .ZN(n3183) );
  AOI22D1BWP30P140LVT U3585 ( .A1(i_data_bus[57]), .A2(n3305), .B1(
        i_data_bus[761]), .B2(n2659), .ZN(n3182) );
  ND4D1BWP30P140LVT U3586 ( .A1(n3185), .A2(n3184), .A3(n3183), .A4(n3182), 
        .ZN(n3192) );
  INVD1BWP30P140LVT U3587 ( .I(i_data_bus[409]), .ZN(n6029) );
  INVD1BWP30P140LVT U3588 ( .I(i_data_bus[505]), .ZN(n5286) );
  OAI22D1BWP30P140LVT U3589 ( .A1(n6029), .A2(n3288), .B1(n5286), .B2(n3267), 
        .ZN(n3191) );
  AOI22D1BWP30P140LVT U3590 ( .A1(i_data_bus[473]), .A2(n3330), .B1(
        i_data_bus[249]), .B2(n3328), .ZN(n3189) );
  AOI22D1BWP30P140LVT U3591 ( .A1(i_data_bus[185]), .A2(n2678), .B1(
        i_data_bus[441]), .B2(n3303), .ZN(n3188) );
  AOI22D1BWP30P140LVT U3592 ( .A1(i_data_bus[569]), .A2(n3332), .B1(
        i_data_bus[633]), .B2(n3333), .ZN(n3187) );
  AOI22D1BWP30P140LVT U3593 ( .A1(i_data_bus[601]), .A2(n3334), .B1(
        i_data_bus[537]), .B2(n3331), .ZN(n3186) );
  ND4D1BWP30P140LVT U3594 ( .A1(n3189), .A2(n3188), .A3(n3187), .A4(n3186), 
        .ZN(n3190) );
  NR4D0BWP30P140LVT U3595 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), 
        .ZN(n3194) );
  ND4D1BWP30P140LVT U3596 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), 
        .ZN(o_data_bus[185]) );
  AOI22D1BWP30P140LVT U3597 ( .A1(i_data_bus[922]), .A2(n3309), .B1(
        i_data_bus[378]), .B2(n3321), .ZN(n3217) );
  AOI22D1BWP30P140LVT U3598 ( .A1(i_data_bus[954]), .A2(n3311), .B1(
        i_data_bus[986]), .B2(n3301), .ZN(n3216) );
  AOI22D1BWP30P140LVT U3599 ( .A1(i_data_bus[250]), .A2(n3328), .B1(
        i_data_bus[474]), .B2(n3330), .ZN(n3215) );
  AOI22D1BWP30P140LVT U3600 ( .A1(i_data_bus[858]), .A2(n3316), .B1(
        i_data_bus[346]), .B2(n3306), .ZN(n3201) );
  AOI22D1BWP30P140LVT U3601 ( .A1(i_data_bus[58]), .A2(n3305), .B1(
        i_data_bus[826]), .B2(n3304), .ZN(n3200) );
  AOI22D1BWP30P140LVT U3602 ( .A1(i_data_bus[90]), .A2(n3317), .B1(
        i_data_bus[762]), .B2(n2659), .ZN(n3199) );
  AOI22D1BWP30P140LVT U3603 ( .A1(i_data_bus[1018]), .A2(n59), .B1(
        i_data_bus[666]), .B2(n3302), .ZN(n3198) );
  ND4D1BWP30P140LVT U3604 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), 
        .ZN(n3213) );
  AOI22D1BWP30P140LVT U3605 ( .A1(i_data_bus[122]), .A2(n3308), .B1(
        i_data_bus[314]), .B2(n3322), .ZN(n3205) );
  AOI22D1BWP30P140LVT U3606 ( .A1(i_data_bus[890]), .A2(n113), .B1(
        i_data_bus[730]), .B2(n3310), .ZN(n3204) );
  AOI22D1BWP30P140LVT U3607 ( .A1(i_data_bus[282]), .A2(n3318), .B1(
        i_data_bus[794]), .B2(n3307), .ZN(n3203) );
  AOI22D1BWP30P140LVT U3608 ( .A1(i_data_bus[26]), .A2(n3319), .B1(
        i_data_bus[698]), .B2(n2653), .ZN(n3202) );
  ND4D1BWP30P140LVT U3609 ( .A1(n3205), .A2(n3204), .A3(n3203), .A4(n3202), 
        .ZN(n3212) );
  INVD1BWP30P140LVT U3610 ( .I(i_data_bus[410]), .ZN(n5307) );
  MOAI22D1BWP30P140LVT U3611 ( .A1(n5307), .A2(n3288), .B1(i_data_bus[186]), 
        .B2(n2678), .ZN(n3211) );
  AOI22D1BWP30P140LVT U3612 ( .A1(i_data_bus[442]), .A2(n3303), .B1(
        i_data_bus[154]), .B2(n2935), .ZN(n3209) );
  AOI22D1BWP30P140LVT U3613 ( .A1(i_data_bus[218]), .A2(n2676), .B1(
        i_data_bus[506]), .B2(n3329), .ZN(n3208) );
  AOI22D1BWP30P140LVT U3614 ( .A1(i_data_bus[634]), .A2(n3333), .B1(
        i_data_bus[570]), .B2(n3332), .ZN(n3207) );
  AOI22D1BWP30P140LVT U3615 ( .A1(i_data_bus[602]), .A2(n3334), .B1(
        i_data_bus[538]), .B2(n3331), .ZN(n3206) );
  ND4D1BWP30P140LVT U3616 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), 
        .ZN(n3210) );
  NR4D0BWP30P140LVT U3617 ( .A1(n3213), .A2(n3212), .A3(n3211), .A4(n3210), 
        .ZN(n3214) );
  ND4D1BWP30P140LVT U3618 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), 
        .ZN(o_data_bus[186]) );
  AOI22D1BWP30P140LVT U3619 ( .A1(i_data_bus[731]), .A2(n3310), .B1(
        i_data_bus[827]), .B2(n3304), .ZN(n3237) );
  AOI22D1BWP30P140LVT U3620 ( .A1(i_data_bus[91]), .A2(n3317), .B1(
        i_data_bus[347]), .B2(n3306), .ZN(n3236) );
  AOI22D1BWP30P140LVT U3621 ( .A1(i_data_bus[507]), .A2(n3329), .B1(
        i_data_bus[251]), .B2(n3328), .ZN(n3235) );
  AOI22D1BWP30P140LVT U3622 ( .A1(i_data_bus[315]), .A2(n3322), .B1(
        i_data_bus[795]), .B2(n3307), .ZN(n3221) );
  AOI22D1BWP30P140LVT U3623 ( .A1(i_data_bus[987]), .A2(n3301), .B1(
        i_data_bus[1019]), .B2(n59), .ZN(n3220) );
  AOI22D1BWP30P140LVT U3624 ( .A1(i_data_bus[667]), .A2(n3302), .B1(
        i_data_bus[699]), .B2(n2653), .ZN(n3219) );
  ND4D1BWP30P140LVT U3625 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), 
        .ZN(n3233) );
  AOI22D1BWP30P140LVT U3626 ( .A1(i_data_bus[123]), .A2(n3308), .B1(
        i_data_bus[283]), .B2(n3318), .ZN(n3225) );
  AOI22D1BWP30P140LVT U3627 ( .A1(i_data_bus[923]), .A2(n3309), .B1(
        i_data_bus[59]), .B2(n3305), .ZN(n3224) );
  AOI22D1BWP30P140LVT U3628 ( .A1(i_data_bus[955]), .A2(n3311), .B1(
        i_data_bus[891]), .B2(n113), .ZN(n3223) );
  AOI22D1BWP30P140LVT U3629 ( .A1(i_data_bus[27]), .A2(n3319), .B1(
        i_data_bus[763]), .B2(n2659), .ZN(n3222) );
  ND4D1BWP30P140LVT U3630 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), 
        .ZN(n3232) );
  INVD1BWP30P140LVT U3631 ( .I(i_data_bus[187]), .ZN(n6071) );
  MOAI22D1BWP30P140LVT U3632 ( .A1(n6071), .A2(n3327), .B1(i_data_bus[219]), 
        .B2(n2676), .ZN(n3231) );
  AOI22D1BWP30P140LVT U3633 ( .A1(i_data_bus[411]), .A2(n3), .B1(
        i_data_bus[443]), .B2(n3303), .ZN(n3229) );
  AOI22D1BWP30P140LVT U3634 ( .A1(i_data_bus[539]), .A2(n3331), .B1(
        i_data_bus[635]), .B2(n3333), .ZN(n3227) );
  AOI22D1BWP30P140LVT U3635 ( .A1(i_data_bus[571]), .A2(n3332), .B1(
        i_data_bus[603]), .B2(n3334), .ZN(n3226) );
  ND4D1BWP30P140LVT U3636 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), 
        .ZN(n3230) );
  NR4D0BWP30P140LVT U3637 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), 
        .ZN(n3234) );
  ND4D1BWP30P140LVT U3638 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3234), 
        .ZN(o_data_bus[187]) );
  AOI22D1BWP30P140LVT U3639 ( .A1(i_data_bus[60]), .A2(n3305), .B1(
        i_data_bus[860]), .B2(n3316), .ZN(n3258) );
  AOI22D1BWP30P140LVT U3640 ( .A1(i_data_bus[924]), .A2(n3309), .B1(
        i_data_bus[348]), .B2(n3306), .ZN(n3257) );
  AOI22D1BWP30P140LVT U3641 ( .A1(i_data_bus[252]), .A2(n3328), .B1(
        i_data_bus[188]), .B2(n2678), .ZN(n3256) );
  AOI22D1BWP30P140LVT U3642 ( .A1(i_data_bus[92]), .A2(n3317), .B1(
        i_data_bus[700]), .B2(n2653), .ZN(n3241) );
  AOI22D1BWP30P140LVT U3643 ( .A1(i_data_bus[988]), .A2(n3301), .B1(
        i_data_bus[668]), .B2(n3302), .ZN(n3240) );
  AOI22D1BWP30P140LVT U3644 ( .A1(i_data_bus[1020]), .A2(n58), .B1(
        i_data_bus[892]), .B2(n113), .ZN(n3239) );
  AOI22D1BWP30P140LVT U3645 ( .A1(i_data_bus[956]), .A2(n3311), .B1(
        i_data_bus[732]), .B2(n3310), .ZN(n3238) );
  ND4D1BWP30P140LVT U3646 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), 
        .ZN(n3254) );
  AOI22D1BWP30P140LVT U3647 ( .A1(i_data_bus[28]), .A2(n3319), .B1(
        i_data_bus[828]), .B2(n3304), .ZN(n3245) );
  AOI22D1BWP30P140LVT U3648 ( .A1(i_data_bus[124]), .A2(n3308), .B1(
        i_data_bus[764]), .B2(n2659), .ZN(n3244) );
  AOI22D1BWP30P140LVT U3649 ( .A1(i_data_bus[284]), .A2(n3318), .B1(
        i_data_bus[316]), .B2(n3322), .ZN(n3243) );
  AOI22D1BWP30P140LVT U3650 ( .A1(i_data_bus[380]), .A2(n3321), .B1(
        i_data_bus[796]), .B2(n3307), .ZN(n3242) );
  ND4D1BWP30P140LVT U3651 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), 
        .ZN(n3253) );
  INVD1BWP30P140LVT U3652 ( .I(i_data_bus[476]), .ZN(n3960) );
  MOAI22D1BWP30P140LVT U3653 ( .A1(n3960), .A2(n3246), .B1(i_data_bus[156]), 
        .B2(n2935), .ZN(n3252) );
  AOI22D1BWP30P140LVT U3654 ( .A1(i_data_bus[508]), .A2(n3329), .B1(
        i_data_bus[412]), .B2(n3), .ZN(n3250) );
  AOI22D1BWP30P140LVT U3655 ( .A1(i_data_bus[444]), .A2(n3303), .B1(
        i_data_bus[220]), .B2(n2676), .ZN(n3249) );
  AOI22D1BWP30P140LVT U3656 ( .A1(i_data_bus[604]), .A2(n3334), .B1(
        i_data_bus[572]), .B2(n3332), .ZN(n3248) );
  AOI22D1BWP30P140LVT U3657 ( .A1(i_data_bus[540]), .A2(n3331), .B1(
        i_data_bus[636]), .B2(n3333), .ZN(n3247) );
  ND4D1BWP30P140LVT U3658 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), 
        .ZN(n3251) );
  NR4D0BWP30P140LVT U3659 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), 
        .ZN(n3255) );
  ND4D1BWP30P140LVT U3660 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), 
        .ZN(o_data_bus[188]) );
  AOI22D1BWP30P140LVT U3661 ( .A1(i_data_bus[1021]), .A2(n58), .B1(
        i_data_bus[861]), .B2(n3316), .ZN(n3279) );
  AOI22D1BWP30P140LVT U3662 ( .A1(i_data_bus[957]), .A2(n7), .B1(
        i_data_bus[797]), .B2(n3307), .ZN(n3278) );
  AOI22D1BWP30P140LVT U3663 ( .A1(i_data_bus[477]), .A2(n3330), .B1(
        i_data_bus[221]), .B2(n2676), .ZN(n3277) );
  AOI22D1BWP30P140LVT U3664 ( .A1(i_data_bus[125]), .A2(n3308), .B1(
        i_data_bus[893]), .B2(n113), .ZN(n3262) );
  AOI22D1BWP30P140LVT U3665 ( .A1(i_data_bus[29]), .A2(n3319), .B1(
        i_data_bus[317]), .B2(n3322), .ZN(n3261) );
  AOI22D1BWP30P140LVT U3666 ( .A1(i_data_bus[989]), .A2(n3301), .B1(
        i_data_bus[381]), .B2(n3321), .ZN(n3260) );
  AOI22D1BWP30P140LVT U3667 ( .A1(i_data_bus[701]), .A2(n2653), .B1(
        i_data_bus[733]), .B2(n3310), .ZN(n3259) );
  ND4D1BWP30P140LVT U3668 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), 
        .ZN(n3275) );
  AOI22D1BWP30P140LVT U3669 ( .A1(i_data_bus[61]), .A2(n3305), .B1(
        i_data_bus[669]), .B2(n3302), .ZN(n3266) );
  AOI22D1BWP30P140LVT U3670 ( .A1(i_data_bus[925]), .A2(n3309), .B1(
        i_data_bus[349]), .B2(n3306), .ZN(n3265) );
  AOI22D1BWP30P140LVT U3671 ( .A1(i_data_bus[93]), .A2(n3317), .B1(
        i_data_bus[829]), .B2(n3304), .ZN(n3264) );
  AOI22D1BWP30P140LVT U3672 ( .A1(i_data_bus[765]), .A2(n2659), .B1(
        i_data_bus[285]), .B2(n3318), .ZN(n3263) );
  ND4D1BWP30P140LVT U3673 ( .A1(n3266), .A2(n3265), .A3(n3264), .A4(n3263), 
        .ZN(n3274) );
  INVD1BWP30P140LVT U3674 ( .I(i_data_bus[509]), .ZN(n3985) );
  MOAI22D1BWP30P140LVT U3675 ( .A1(n3985), .A2(n3267), .B1(i_data_bus[413]), 
        .B2(n3), .ZN(n3273) );
  AOI22D1BWP30P140LVT U3676 ( .A1(i_data_bus[445]), .A2(n3303), .B1(
        i_data_bus[189]), .B2(n2678), .ZN(n3271) );
  AOI22D1BWP30P140LVT U3677 ( .A1(i_data_bus[157]), .A2(n2935), .B1(
        i_data_bus[253]), .B2(n3328), .ZN(n3270) );
  AOI22D1BWP30P140LVT U3678 ( .A1(i_data_bus[573]), .A2(n3332), .B1(
        i_data_bus[541]), .B2(n3331), .ZN(n3269) );
  AOI22D1BWP30P140LVT U3679 ( .A1(i_data_bus[637]), .A2(n3333), .B1(
        i_data_bus[605]), .B2(n3334), .ZN(n3268) );
  ND4D1BWP30P140LVT U3680 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), 
        .ZN(n3272) );
  NR4D0BWP30P140LVT U3681 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), 
        .ZN(n3276) );
  ND4D1BWP30P140LVT U3682 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), 
        .ZN(o_data_bus[189]) );
  AOI22D1BWP30P140LVT U3683 ( .A1(i_data_bus[926]), .A2(n3309), .B1(
        i_data_bus[62]), .B2(n3305), .ZN(n3300) );
  AOI22D1BWP30P140LVT U3684 ( .A1(i_data_bus[30]), .A2(n3319), .B1(
        i_data_bus[734]), .B2(n3310), .ZN(n3299) );
  AOI22D1BWP30P140LVT U3685 ( .A1(i_data_bus[222]), .A2(n2676), .B1(
        i_data_bus[158]), .B2(n2935), .ZN(n3298) );
  AOI22D1BWP30P140LVT U3686 ( .A1(i_data_bus[798]), .A2(n3307), .B1(
        i_data_bus[766]), .B2(n2659), .ZN(n3283) );
  AOI22D1BWP30P140LVT U3687 ( .A1(i_data_bus[990]), .A2(n3301), .B1(
        i_data_bus[702]), .B2(n2653), .ZN(n3282) );
  AOI22D1BWP30P140LVT U3688 ( .A1(i_data_bus[670]), .A2(n3302), .B1(
        i_data_bus[894]), .B2(n113), .ZN(n3281) );
  AOI22D1BWP30P140LVT U3689 ( .A1(i_data_bus[862]), .A2(n3316), .B1(
        i_data_bus[382]), .B2(n3321), .ZN(n3280) );
  ND4D1BWP30P140LVT U3690 ( .A1(n3280), .A2(n3282), .A3(n3281), .A4(n3283), 
        .ZN(n3296) );
  AOI22D1BWP30P140LVT U3691 ( .A1(i_data_bus[958]), .A2(n3311), .B1(
        i_data_bus[830]), .B2(n3304), .ZN(n3287) );
  AOI22D1BWP30P140LVT U3692 ( .A1(i_data_bus[126]), .A2(n3308), .B1(
        i_data_bus[318]), .B2(n3322), .ZN(n3286) );
  AOI22D1BWP30P140LVT U3693 ( .A1(i_data_bus[1022]), .A2(n59), .B1(
        i_data_bus[286]), .B2(n3318), .ZN(n3285) );
  AOI22D1BWP30P140LVT U3694 ( .A1(i_data_bus[94]), .A2(n3317), .B1(
        i_data_bus[350]), .B2(n3306), .ZN(n3284) );
  ND4D1BWP30P140LVT U3695 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), 
        .ZN(n3295) );
  INVD1BWP30P140LVT U3696 ( .I(i_data_bus[414]), .ZN(n6138) );
  MOAI22D1BWP30P140LVT U3697 ( .A1(n6138), .A2(n3288), .B1(i_data_bus[510]), 
        .B2(n3329), .ZN(n3294) );
  AOI22D1BWP30P140LVT U3698 ( .A1(i_data_bus[446]), .A2(n3303), .B1(
        i_data_bus[254]), .B2(n3328), .ZN(n3292) );
  AOI22D1BWP30P140LVT U3699 ( .A1(i_data_bus[190]), .A2(n2678), .B1(
        i_data_bus[478]), .B2(n3330), .ZN(n3291) );
  AOI22D1BWP30P140LVT U3700 ( .A1(i_data_bus[606]), .A2(n3334), .B1(
        i_data_bus[638]), .B2(n3333), .ZN(n3290) );
  AOI22D1BWP30P140LVT U3701 ( .A1(i_data_bus[542]), .A2(n3331), .B1(
        i_data_bus[574]), .B2(n3332), .ZN(n3289) );
  ND4D1BWP30P140LVT U3702 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), 
        .ZN(n3293) );
  NR4D0BWP30P140LVT U3703 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), 
        .ZN(n3297) );
  ND4D1BWP30P140LVT U3704 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), 
        .ZN(o_data_bus[190]) );
  AOI22D1BWP30P140LVT U3705 ( .A1(i_data_bus[991]), .A2(n3301), .B1(
        i_data_bus[703]), .B2(n2653), .ZN(n3346) );
  AOI22D1BWP30P140LVT U3706 ( .A1(i_data_bus[671]), .A2(n3302), .B1(
        i_data_bus[767]), .B2(n2659), .ZN(n3345) );
  AOI22D1BWP30P140LVT U3707 ( .A1(i_data_bus[447]), .A2(n3303), .B1(
        i_data_bus[159]), .B2(n2935), .ZN(n3344) );
  AOI22D1BWP30P140LVT U3708 ( .A1(i_data_bus[63]), .A2(n3305), .B1(
        i_data_bus[831]), .B2(n3304), .ZN(n3315) );
  AOI22D1BWP30P140LVT U3709 ( .A1(i_data_bus[799]), .A2(n3307), .B1(
        i_data_bus[351]), .B2(n3306), .ZN(n3314) );
  AOI22D1BWP30P140LVT U3710 ( .A1(i_data_bus[927]), .A2(n3309), .B1(
        i_data_bus[127]), .B2(n3308), .ZN(n3313) );
  AOI22D1BWP30P140LVT U3711 ( .A1(i_data_bus[959]), .A2(n3311), .B1(
        i_data_bus[735]), .B2(n3310), .ZN(n3312) );
  ND4D1BWP30P140LVT U3712 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), 
        .ZN(n3342) );
  AOI22D1BWP30P140LVT U3713 ( .A1(i_data_bus[31]), .A2(n3319), .B1(
        i_data_bus[287]), .B2(n3318), .ZN(n3325) );
  AOI22D1BWP30P140LVT U3714 ( .A1(i_data_bus[1023]), .A2(n59), .B1(
        i_data_bus[895]), .B2(n113), .ZN(n3324) );
  AOI22D1BWP30P140LVT U3715 ( .A1(i_data_bus[319]), .A2(n3322), .B1(
        i_data_bus[383]), .B2(n3321), .ZN(n3323) );
  ND4D1BWP30P140LVT U3716 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), 
        .ZN(n3341) );
  INVD1BWP30P140LVT U3717 ( .I(i_data_bus[191]), .ZN(n6176) );
  MOAI22D1BWP30P140LVT U3718 ( .A1(n6176), .A2(n3327), .B1(i_data_bus[223]), 
        .B2(n2676), .ZN(n3340) );
  AOI22D1BWP30P140LVT U3719 ( .A1(i_data_bus[511]), .A2(n3329), .B1(
        i_data_bus[255]), .B2(n3328), .ZN(n3338) );
  AOI22D1BWP30P140LVT U3720 ( .A1(i_data_bus[415]), .A2(n3), .B1(
        i_data_bus[479]), .B2(n3330), .ZN(n3337) );
  AOI22D1BWP30P140LVT U3721 ( .A1(i_data_bus[575]), .A2(n3332), .B1(
        i_data_bus[543]), .B2(n3331), .ZN(n3336) );
  AOI22D1BWP30P140LVT U3722 ( .A1(i_data_bus[607]), .A2(n3334), .B1(
        i_data_bus[639]), .B2(n3333), .ZN(n3335) );
  ND4D1BWP30P140LVT U3723 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), 
        .ZN(n3339) );
  NR4D0BWP30P140LVT U3724 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), 
        .ZN(n3343) );
  ND4D1BWP30P140LVT U3725 ( .A1(n3346), .A2(n3345), .A3(n3344), .A4(n3343), 
        .ZN(o_data_bus[191]) );
  ND3D1BWP30P140LVT U3726 ( .A1(i_valid[9]), .A2(i_cmd[74]), .A3(n3371), .ZN(
        n3878) );
  ND3D1BWP30P140LVT U3727 ( .A1(i_valid[10]), .A2(i_cmd[82]), .A3(n3371), .ZN(
        n3961) );
  AOI22D1BWP30P140LVT U3728 ( .A1(i_data_bus[288]), .A2(n3347), .B1(
        i_data_bus[320]), .B2(n3348), .ZN(n3396) );
  ND3D1BWP30P140LVT U3729 ( .A1(i_valid[11]), .A2(i_cmd[90]), .A3(n3371), .ZN(
        n3983) );
  INVD2BWP30P140LVT U3730 ( .I(n3983), .ZN(n4033) );
  AOI22D1BWP30P140LVT U3731 ( .A1(i_data_bus[384]), .A2(n4022), .B1(
        i_data_bus[352]), .B2(n4033), .ZN(n3395) );
  AOI22D1BWP30P140LVT U3732 ( .A1(i_data_bus[832]), .A2(n4036), .B1(
        i_data_bus[864]), .B2(n4039), .ZN(n3359) );
  INVD1BWP30P140LVT U3733 ( .I(i_cmd[162]), .ZN(n3349) );
  NR3D0P7BWP30P140LVT U3734 ( .A1(n5455), .A2(n3349), .A3(n3361), .ZN(n3350)
         );
  AOI22D1BWP30P140LVT U3735 ( .A1(i_data_bus[0]), .A2(n4038), .B1(
        i_data_bus[640]), .B2(n4040), .ZN(n3358) );
  AOI22D1BWP30P140LVT U3736 ( .A1(i_data_bus[192]), .A2(n3351), .B1(
        i_data_bus[224]), .B2(n3352), .ZN(n3357) );
  INVD1BWP30P140LVT U3737 ( .I(i_cmd[34]), .ZN(n3354) );
  AOI22D1BWP30P140LVT U3738 ( .A1(i_data_bus[736]), .A2(n3353), .B1(
        i_data_bus[128]), .B2(n3355), .ZN(n3356) );
  INR3D2BWP30P140LVT U3739 ( .A1(i_cmd[170]), .B1(n5463), .B2(n3361), .ZN(
        n4035) );
  AOI22D1BWP30P140LVT U3740 ( .A1(i_data_bus[704]), .A2(n3360), .B1(
        i_data_bus[672]), .B2(n4035), .ZN(n3369) );
  AOI22D1BWP30P140LVT U3741 ( .A1(i_data_bus[32]), .A2(n4025), .B1(
        i_data_bus[800]), .B2(n4024), .ZN(n3367) );
  INVD1BWP30P140LVT U3742 ( .I(i_cmd[194]), .ZN(n3364) );
  INR3D2BWP30P140LVT U3743 ( .A1(i_cmd[42]), .B1(n5487), .B2(n3365), .ZN(n4037) );
  AOI22D1BWP30P140LVT U3744 ( .A1(i_data_bus[768]), .A2(n4027), .B1(
        i_data_bus[160]), .B2(n4037), .ZN(n3366) );
  ND4D1BWP30P140LVT U3745 ( .A1(n3368), .A2(n3369), .A3(n3367), .A4(n3366), 
        .ZN(n3392) );
  ND3D1BWP30P140LVT U3746 ( .A1(i_valid[14]), .A2(i_cmd[114]), .A3(n3373), 
        .ZN(n4046) );
  INVD1BWP30P140LVT U3747 ( .I(i_data_bus[256]), .ZN(n4766) );
  ND3D1BWP30P140LVT U3748 ( .A1(i_valid[8]), .A2(i_cmd[66]), .A3(n3371), .ZN(
        n3982) );
  OAI22D1BWP30P140LVT U3749 ( .A1(n3372), .A2(n4046), .B1(n4766), .B2(n3982), 
        .ZN(n3391) );
  INVD1BWP30P140LVT U3750 ( .I(i_data_bus[480]), .ZN(n5469) );
  ND3D1BWP30P140LVT U3751 ( .A1(i_valid[15]), .A2(i_cmd[122]), .A3(n3373), 
        .ZN(n3984) );
  ND3D1BWP30P140LVT U3752 ( .A1(i_valid[13]), .A2(i_cmd[106]), .A3(n3373), 
        .ZN(n3856) );
  MOAI22D1BWP30P140LVT U3753 ( .A1(n5469), .A2(n3984), .B1(i_data_bus[416]), 
        .B2(n4021), .ZN(n3390) );
  INR3D2BWP30P140LVT U3754 ( .A1(i_cmd[138]), .B1(n5479), .B2(n3384), .ZN(
        n4047) );
  AOI22D1BWP30P140LVT U3755 ( .A1(i_data_bus[544]), .A2(n4047), .B1(
        i_data_bus[960]), .B2(n4048), .ZN(n3388) );
  NR3D0P7BWP30P140LVT U3756 ( .A1(n5486), .A2(n3375), .A3(n3381), .ZN(n3376)
         );
  AOI22D1BWP30P140LVT U3757 ( .A1(i_data_bus[928]), .A2(n4051), .B1(
        i_data_bus[896]), .B2(n3378), .ZN(n3387) );
  INVD1BWP30P140LVT U3758 ( .I(n3379), .ZN(n3380) );
  INR3D2BWP30P140LVT U3759 ( .A1(i_cmd[154]), .B1(n5478), .B2(n3384), .ZN(
        n4049) );
  AOI22D1BWP30P140LVT U3760 ( .A1(i_data_bus[512]), .A2(n4052), .B1(
        i_data_bus[608]), .B2(n4049), .ZN(n3386) );
  INR3D2BWP30P140LVT U3761 ( .A1(i_cmd[146]), .B1(n5481), .B2(n3384), .ZN(
        n4050) );
  AOI22D1BWP30P140LVT U3762 ( .A1(i_data_bus[992]), .A2(n3383), .B1(
        i_data_bus[576]), .B2(n4050), .ZN(n3385) );
  ND4D1BWP30P140LVT U3763 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), 
        .ZN(n3389) );
  NR4D0BWP30P140LVT U3764 ( .A1(n3392), .A2(n3391), .A3(n3390), .A4(n3389), 
        .ZN(n3393) );
  ND4D1BWP30P140LVT U3765 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), 
        .ZN(o_data_bus[64]) );
  AOI22D1BWP30P140LVT U3766 ( .A1(i_data_bus[449]), .A2(n4006), .B1(
        i_data_bus[417]), .B2(n4021), .ZN(n3416) );
  AOI22D1BWP30P140LVT U3767 ( .A1(i_data_bus[353]), .A2(n4033), .B1(
        i_data_bus[321]), .B2(n3348), .ZN(n3415) );
  AOI22D1BWP30P140LVT U3768 ( .A1(i_data_bus[97]), .A2(n4026), .B1(
        i_data_bus[705]), .B2(n3360), .ZN(n3400) );
  AOI22D1BWP30P140LVT U3769 ( .A1(i_data_bus[129]), .A2(n3355), .B1(
        i_data_bus[833]), .B2(n4036), .ZN(n3399) );
  AOI22D1BWP30P140LVT U3770 ( .A1(i_data_bus[161]), .A2(n4037), .B1(
        i_data_bus[225]), .B2(n3352), .ZN(n3398) );
  AOI22D1BWP30P140LVT U3771 ( .A1(i_data_bus[65]), .A2(n4028), .B1(
        i_data_bus[801]), .B2(n4024), .ZN(n3397) );
  AOI22D1BWP30P140LVT U3772 ( .A1(i_data_bus[769]), .A2(n4027), .B1(
        i_data_bus[673]), .B2(n4035), .ZN(n3404) );
  AOI22D1BWP30P140LVT U3773 ( .A1(i_data_bus[737]), .A2(n3353), .B1(
        i_data_bus[193]), .B2(n3351), .ZN(n3403) );
  AOI22D1BWP30P140LVT U3774 ( .A1(i_data_bus[1]), .A2(n4038), .B1(
        i_data_bus[865]), .B2(n4039), .ZN(n3402) );
  AOI22D1BWP30P140LVT U3775 ( .A1(i_data_bus[33]), .A2(n4025), .B1(
        i_data_bus[641]), .B2(n4040), .ZN(n3401) );
  ND4D1BWP30P140LVT U3776 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), 
        .ZN(n3412) );
  INVD1BWP30P140LVT U3777 ( .I(i_data_bus[257]), .ZN(n4787) );
  MOAI22D1BWP30P140LVT U3778 ( .A1(n4787), .A2(n3982), .B1(i_data_bus[289]), 
        .B2(n3347), .ZN(n3411) );
  MOAI22D1BWP30P140LVT U3779 ( .A1(n5514), .A2(n3984), .B1(i_data_bus[385]), 
        .B2(n4022), .ZN(n3410) );
  AOI22D1BWP30P140LVT U3780 ( .A1(i_data_bus[577]), .A2(n4050), .B1(
        i_data_bus[993]), .B2(n3383), .ZN(n3408) );
  AOI22D1BWP30P140LVT U3781 ( .A1(i_data_bus[897]), .A2(n3378), .B1(
        i_data_bus[513]), .B2(n4052), .ZN(n3407) );
  AOI22D1BWP30P140LVT U3782 ( .A1(i_data_bus[961]), .A2(n4048), .B1(
        i_data_bus[609]), .B2(n4049), .ZN(n3406) );
  AOI22D1BWP30P140LVT U3783 ( .A1(i_data_bus[545]), .A2(n4047), .B1(
        i_data_bus[929]), .B2(n4051), .ZN(n3405) );
  ND4D1BWP30P140LVT U3784 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), 
        .ZN(n3409) );
  NR4D0BWP30P140LVT U3785 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), 
        .ZN(n3413) );
  ND4D1BWP30P140LVT U3786 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), 
        .ZN(o_data_bus[65]) );
  AOI22D1BWP30P140LVT U3787 ( .A1(i_data_bus[386]), .A2(n4022), .B1(
        i_data_bus[354]), .B2(n4033), .ZN(n3437) );
  AOI22D1BWP30P140LVT U3788 ( .A1(i_data_bus[290]), .A2(n3347), .B1(
        i_data_bus[418]), .B2(n4021), .ZN(n3436) );
  AOI22D1BWP30P140LVT U3789 ( .A1(i_data_bus[162]), .A2(n4037), .B1(
        i_data_bus[130]), .B2(n3355), .ZN(n3420) );
  AOI22D1BWP30P140LVT U3790 ( .A1(i_data_bus[738]), .A2(n3353), .B1(
        i_data_bus[706]), .B2(n3360), .ZN(n3419) );
  AOI22D1BWP30P140LVT U3791 ( .A1(i_data_bus[34]), .A2(n4025), .B1(
        i_data_bus[194]), .B2(n3351), .ZN(n3418) );
  AOI22D1BWP30P140LVT U3792 ( .A1(i_data_bus[866]), .A2(n4039), .B1(
        i_data_bus[834]), .B2(n4036), .ZN(n3417) );
  AOI22D1BWP30P140LVT U3793 ( .A1(i_data_bus[98]), .A2(n4026), .B1(
        i_data_bus[226]), .B2(n3352), .ZN(n3424) );
  AOI22D1BWP30P140LVT U3794 ( .A1(i_data_bus[2]), .A2(n4038), .B1(
        i_data_bus[642]), .B2(n4040), .ZN(n3423) );
  AOI22D1BWP30P140LVT U3795 ( .A1(i_data_bus[802]), .A2(n4024), .B1(
        i_data_bus[770]), .B2(n4027), .ZN(n3422) );
  AOI22D1BWP30P140LVT U3796 ( .A1(i_data_bus[66]), .A2(n4028), .B1(
        i_data_bus[674]), .B2(n4035), .ZN(n3421) );
  ND4D1BWP30P140LVT U3797 ( .A1(n3424), .A2(n3423), .A3(n3422), .A4(n3421), 
        .ZN(n3433) );
  INVD1BWP30P140LVT U3798 ( .I(i_data_bus[322]), .ZN(n4808) );
  OAI22D1BWP30P140LVT U3799 ( .A1(n3425), .A2(n4046), .B1(n4808), .B2(n3961), 
        .ZN(n3432) );
  INVD1BWP30P140LVT U3800 ( .I(i_data_bus[258]), .ZN(n5535) );
  MOAI22D1BWP30P140LVT U3801 ( .A1(n5535), .A2(n3982), .B1(i_data_bus[482]), 
        .B2(n4020), .ZN(n3431) );
  AOI22D1BWP30P140LVT U3802 ( .A1(i_data_bus[578]), .A2(n4050), .B1(
        i_data_bus[610]), .B2(n4049), .ZN(n3429) );
  AOI22D1BWP30P140LVT U3803 ( .A1(i_data_bus[546]), .A2(n4047), .B1(
        i_data_bus[898]), .B2(n3378), .ZN(n3428) );
  AOI22D1BWP30P140LVT U3804 ( .A1(i_data_bus[962]), .A2(n4048), .B1(
        i_data_bus[514]), .B2(n4052), .ZN(n3427) );
  AOI22D1BWP30P140LVT U3805 ( .A1(i_data_bus[994]), .A2(n3383), .B1(
        i_data_bus[930]), .B2(n4051), .ZN(n3426) );
  ND4D1BWP30P140LVT U3806 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), 
        .ZN(n3430) );
  NR4D0BWP30P140LVT U3807 ( .A1(n3433), .A2(n3432), .A3(n3431), .A4(n3430), 
        .ZN(n3434) );
  ND4D1BWP30P140LVT U3808 ( .A1(n3437), .A2(n3436), .A3(n3435), .A4(n3434), 
        .ZN(o_data_bus[66]) );
  AOI22D1BWP30P140LVT U3809 ( .A1(i_data_bus[323]), .A2(n3348), .B1(
        i_data_bus[291]), .B2(n3347), .ZN(n3459) );
  AOI22D1BWP30P140LVT U3810 ( .A1(i_data_bus[387]), .A2(n4022), .B1(
        i_data_bus[483]), .B2(n4020), .ZN(n3458) );
  AOI22D1BWP30P140LVT U3811 ( .A1(i_data_bus[227]), .A2(n3352), .B1(
        i_data_bus[195]), .B2(n3351), .ZN(n3441) );
  AOI22D1BWP30P140LVT U3812 ( .A1(i_data_bus[643]), .A2(n4040), .B1(
        i_data_bus[867]), .B2(n4039), .ZN(n3440) );
  AOI22D1BWP30P140LVT U3813 ( .A1(i_data_bus[35]), .A2(n4025), .B1(
        i_data_bus[835]), .B2(n4036), .ZN(n3439) );
  AOI22D1BWP30P140LVT U3814 ( .A1(i_data_bus[3]), .A2(n4038), .B1(
        i_data_bus[99]), .B2(n4026), .ZN(n3438) );
  AOI22D1BWP30P140LVT U3815 ( .A1(i_data_bus[163]), .A2(n4037), .B1(
        i_data_bus[803]), .B2(n4024), .ZN(n3445) );
  AOI22D1BWP30P140LVT U3816 ( .A1(i_data_bus[131]), .A2(n3355), .B1(
        i_data_bus[675]), .B2(n4035), .ZN(n3444) );
  AOI22D1BWP30P140LVT U3817 ( .A1(i_data_bus[771]), .A2(n4027), .B1(
        i_data_bus[739]), .B2(n3353), .ZN(n3443) );
  AOI22D1BWP30P140LVT U3818 ( .A1(i_data_bus[67]), .A2(n4028), .B1(
        i_data_bus[707]), .B2(n3360), .ZN(n3442) );
  ND4D1BWP30P140LVT U3819 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), 
        .ZN(n3455) );
  MOAI22D1BWP30P140LVT U3820 ( .A1(n3446), .A2(n4046), .B1(i_data_bus[355]), 
        .B2(n4033), .ZN(n3454) );
  INVD1BWP30P140LVT U3821 ( .I(i_data_bus[419]), .ZN(n5558) );
  BUFFD2BWP30P140LVT U3822 ( .I(n3447), .Z(n4023) );
  MOAI22D1BWP30P140LVT U3823 ( .A1(n5558), .A2(n3856), .B1(i_data_bus[259]), 
        .B2(n4023), .ZN(n3453) );
  AOI22D1BWP30P140LVT U3824 ( .A1(i_data_bus[515]), .A2(n4052), .B1(
        i_data_bus[995]), .B2(n3383), .ZN(n3451) );
  AOI22D1BWP30P140LVT U3825 ( .A1(i_data_bus[899]), .A2(n3378), .B1(
        i_data_bus[611]), .B2(n4049), .ZN(n3450) );
  AOI22D1BWP30P140LVT U3826 ( .A1(i_data_bus[963]), .A2(n4048), .B1(
        i_data_bus[931]), .B2(n4051), .ZN(n3449) );
  AOI22D1BWP30P140LVT U3827 ( .A1(i_data_bus[579]), .A2(n4050), .B1(
        i_data_bus[547]), .B2(n4047), .ZN(n3448) );
  ND4D1BWP30P140LVT U3828 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), 
        .ZN(n3452) );
  NR4D0BWP30P140LVT U3829 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), 
        .ZN(n3456) );
  ND4D1BWP30P140LVT U3830 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), 
        .ZN(o_data_bus[67]) );
  AOI22D1BWP30P140LVT U3831 ( .A1(i_data_bus[420]), .A2(n4021), .B1(
        i_data_bus[292]), .B2(n3347), .ZN(n3480) );
  AOI22D1BWP30P140LVT U3832 ( .A1(i_data_bus[356]), .A2(n4033), .B1(
        i_data_bus[260]), .B2(n4023), .ZN(n3479) );
  AOI22D1BWP30P140LVT U3833 ( .A1(i_data_bus[612]), .A2(n4049), .B1(
        i_data_bus[900]), .B2(n3378), .ZN(n3463) );
  AOI22D1BWP30P140LVT U3834 ( .A1(i_data_bus[548]), .A2(n4047), .B1(
        i_data_bus[932]), .B2(n4051), .ZN(n3462) );
  AOI22D1BWP30P140LVT U3835 ( .A1(i_data_bus[964]), .A2(n4048), .B1(
        i_data_bus[580]), .B2(n4050), .ZN(n3461) );
  AOI22D1BWP30P140LVT U3836 ( .A1(i_data_bus[516]), .A2(n4052), .B1(
        i_data_bus[996]), .B2(n3383), .ZN(n3460) );
  MOAI22D1BWP30P140LVT U3837 ( .A1(n3464), .A2(n4007), .B1(i_data_bus[484]), 
        .B2(n4020), .ZN(n3476) );
  INVD1BWP30P140LVT U3838 ( .I(i_data_bus[324]), .ZN(n4849) );
  OAI22D1BWP30P140LVT U3839 ( .A1(n5579), .A2(n4046), .B1(n4849), .B2(n3961), 
        .ZN(n3475) );
  AOI22D1BWP30P140LVT U3840 ( .A1(i_data_bus[228]), .A2(n3352), .B1(
        i_data_bus[868]), .B2(n4039), .ZN(n3468) );
  AOI22D1BWP30P140LVT U3841 ( .A1(i_data_bus[708]), .A2(n3360), .B1(
        i_data_bus[644]), .B2(n4040), .ZN(n3467) );
  AOI22D1BWP30P140LVT U3842 ( .A1(i_data_bus[4]), .A2(n4038), .B1(
        i_data_bus[740]), .B2(n3353), .ZN(n3466) );
  AOI22D1BWP30P140LVT U3843 ( .A1(i_data_bus[132]), .A2(n3355), .B1(
        i_data_bus[804]), .B2(n4024), .ZN(n3465) );
  ND4D1BWP30P140LVT U3844 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), 
        .ZN(n3474) );
  AOI22D1BWP30P140LVT U3845 ( .A1(i_data_bus[100]), .A2(n4026), .B1(
        i_data_bus[68]), .B2(n4028), .ZN(n3472) );
  AOI22D1BWP30P140LVT U3846 ( .A1(i_data_bus[196]), .A2(n3351), .B1(
        i_data_bus[772]), .B2(n4027), .ZN(n3471) );
  AOI22D1BWP30P140LVT U3847 ( .A1(i_data_bus[36]), .A2(n4025), .B1(
        i_data_bus[836]), .B2(n4036), .ZN(n3470) );
  AOI22D1BWP30P140LVT U3848 ( .A1(i_data_bus[676]), .A2(n4035), .B1(
        i_data_bus[164]), .B2(n4037), .ZN(n3469) );
  ND4D1BWP30P140LVT U3849 ( .A1(n3472), .A2(n3471), .A3(n3470), .A4(n3469), 
        .ZN(n3473) );
  NR4D0BWP30P140LVT U3850 ( .A1(n3473), .A2(n3475), .A3(n3474), .A4(n3476), 
        .ZN(n3477) );
  ND4D1BWP30P140LVT U3851 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), 
        .ZN(o_data_bus[68]) );
  AOI22D1BWP30P140LVT U3852 ( .A1(i_data_bus[421]), .A2(n4021), .B1(
        i_data_bus[261]), .B2(n4023), .ZN(n3500) );
  AOI22D1BWP30P140LVT U3853 ( .A1(i_data_bus[453]), .A2(n4006), .B1(
        i_data_bus[325]), .B2(n3348), .ZN(n3499) );
  AOI22D1BWP30P140LVT U3854 ( .A1(i_data_bus[677]), .A2(n4035), .B1(
        i_data_bus[741]), .B2(n3353), .ZN(n3484) );
  AOI22D1BWP30P140LVT U3855 ( .A1(i_data_bus[37]), .A2(n4025), .B1(
        i_data_bus[709]), .B2(n3360), .ZN(n3483) );
  AOI22D1BWP30P140LVT U3856 ( .A1(i_data_bus[645]), .A2(n4040), .B1(
        i_data_bus[805]), .B2(n4024), .ZN(n3482) );
  AOI22D1BWP30P140LVT U3857 ( .A1(i_data_bus[101]), .A2(n4026), .B1(
        i_data_bus[69]), .B2(n4028), .ZN(n3481) );
  AOI22D1BWP30P140LVT U3858 ( .A1(i_data_bus[357]), .A2(n4033), .B1(
        i_data_bus[389]), .B2(n4022), .ZN(n3496) );
  AOI22D1BWP30P140LVT U3859 ( .A1(i_data_bus[773]), .A2(n4027), .B1(
        i_data_bus[837]), .B2(n4036), .ZN(n3488) );
  AOI22D1BWP30P140LVT U3860 ( .A1(i_data_bus[197]), .A2(n3351), .B1(
        i_data_bus[869]), .B2(n4039), .ZN(n3487) );
  AOI22D1BWP30P140LVT U3861 ( .A1(i_data_bus[165]), .A2(n4037), .B1(
        i_data_bus[229]), .B2(n3352), .ZN(n3486) );
  AOI22D1BWP30P140LVT U3862 ( .A1(i_data_bus[5]), .A2(n4038), .B1(
        i_data_bus[133]), .B2(n3355), .ZN(n3485) );
  ND4D1BWP30P140LVT U3863 ( .A1(n3488), .A2(n3487), .A3(n3486), .A4(n3485), 
        .ZN(n3495) );
  INVD1BWP30P140LVT U3864 ( .I(i_data_bus[293]), .ZN(n5600) );
  MOAI22D1BWP30P140LVT U3865 ( .A1(n5600), .A2(n3878), .B1(i_data_bus[485]), 
        .B2(n4020), .ZN(n3494) );
  AOI22D1BWP30P140LVT U3866 ( .A1(i_data_bus[581]), .A2(n4050), .B1(
        i_data_bus[933]), .B2(n4051), .ZN(n3492) );
  AOI22D1BWP30P140LVT U3867 ( .A1(i_data_bus[901]), .A2(n3378), .B1(
        i_data_bus[549]), .B2(n4047), .ZN(n3491) );
  AOI22D1BWP30P140LVT U3868 ( .A1(i_data_bus[517]), .A2(n4052), .B1(
        i_data_bus[965]), .B2(n4048), .ZN(n3490) );
  AOI22D1BWP30P140LVT U3869 ( .A1(i_data_bus[613]), .A2(n4049), .B1(
        i_data_bus[997]), .B2(n3383), .ZN(n3489) );
  ND4D1BWP30P140LVT U3870 ( .A1(n3492), .A2(n3491), .A3(n3490), .A4(n3489), 
        .ZN(n3493) );
  INR4D0BWP30P140LVT U3871 ( .A1(n3496), .B1(n3495), .B2(n3494), .B3(n3493), 
        .ZN(n3497) );
  ND4D1BWP30P140LVT U3872 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), 
        .ZN(o_data_bus[69]) );
  AOI22D1BWP30P140LVT U3873 ( .A1(i_data_bus[358]), .A2(n4033), .B1(
        i_data_bus[262]), .B2(n4023), .ZN(n3520) );
  AOI22D1BWP30P140LVT U3874 ( .A1(i_data_bus[294]), .A2(n3347), .B1(
        i_data_bus[326]), .B2(n3348), .ZN(n3519) );
  AOI22D1BWP30P140LVT U3875 ( .A1(i_data_bus[582]), .A2(n4050), .B1(
        i_data_bus[998]), .B2(n3383), .ZN(n3504) );
  AOI22D1BWP30P140LVT U3876 ( .A1(i_data_bus[614]), .A2(n4049), .B1(
        i_data_bus[934]), .B2(n4051), .ZN(n3503) );
  AOI22D1BWP30P140LVT U3877 ( .A1(i_data_bus[966]), .A2(n4048), .B1(
        i_data_bus[518]), .B2(n4052), .ZN(n3502) );
  AOI22D1BWP30P140LVT U3878 ( .A1(i_data_bus[550]), .A2(n4047), .B1(
        i_data_bus[902]), .B2(n3378), .ZN(n3501) );
  AOI22D1BWP30P140LVT U3879 ( .A1(i_data_bus[486]), .A2(n4020), .B1(
        i_data_bus[422]), .B2(n4021), .ZN(n3516) );
  INVD1BWP30P140LVT U3880 ( .I(i_data_bus[390]), .ZN(n4890) );
  OAI22D1BWP30P140LVT U3881 ( .A1(n4890), .A2(n4007), .B1(n5621), .B2(n4046), 
        .ZN(n3515) );
  AOI22D1BWP30P140LVT U3882 ( .A1(i_data_bus[38]), .A2(n4025), .B1(
        i_data_bus[806]), .B2(n4024), .ZN(n3508) );
  AOI22D1BWP30P140LVT U3883 ( .A1(i_data_bus[198]), .A2(n3351), .B1(
        i_data_bus[678]), .B2(n4035), .ZN(n3507) );
  AOI22D1BWP30P140LVT U3884 ( .A1(i_data_bus[646]), .A2(n4040), .B1(
        i_data_bus[774]), .B2(n4027), .ZN(n3506) );
  AOI22D1BWP30P140LVT U3885 ( .A1(i_data_bus[6]), .A2(n4038), .B1(
        i_data_bus[230]), .B2(n3352), .ZN(n3505) );
  ND4D1BWP30P140LVT U3886 ( .A1(n3508), .A2(n3507), .A3(n3506), .A4(n3505), 
        .ZN(n3514) );
  AOI22D1BWP30P140LVT U3887 ( .A1(i_data_bus[742]), .A2(n3353), .B1(
        i_data_bus[710]), .B2(n3360), .ZN(n3512) );
  AOI22D1BWP30P140LVT U3888 ( .A1(i_data_bus[70]), .A2(n4028), .B1(
        i_data_bus[870]), .B2(n4039), .ZN(n3511) );
  AOI22D1BWP30P140LVT U3889 ( .A1(i_data_bus[102]), .A2(n4026), .B1(
        i_data_bus[134]), .B2(n3355), .ZN(n3510) );
  AOI22D1BWP30P140LVT U3890 ( .A1(i_data_bus[838]), .A2(n4036), .B1(
        i_data_bus[166]), .B2(n4037), .ZN(n3509) );
  ND4D1BWP30P140LVT U3891 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), 
        .ZN(n3513) );
  INR4D0BWP30P140LVT U3892 ( .A1(n3516), .B1(n3515), .B2(n3514), .B3(n3513), 
        .ZN(n3517) );
  ND4D1BWP30P140LVT U3893 ( .A1(n3520), .A2(n3519), .A3(n3518), .A4(n3517), 
        .ZN(o_data_bus[70]) );
  AOI22D1BWP30P140LVT U3894 ( .A1(i_data_bus[455]), .A2(n4006), .B1(
        i_data_bus[423]), .B2(n4021), .ZN(n3541) );
  AOI22D1BWP30P140LVT U3895 ( .A1(i_data_bus[263]), .A2(n4023), .B1(
        i_data_bus[391]), .B2(n4022), .ZN(n3540) );
  AOI22D1BWP30P140LVT U3896 ( .A1(i_data_bus[903]), .A2(n3378), .B1(
        i_data_bus[967]), .B2(n4048), .ZN(n3524) );
  AOI22D1BWP30P140LVT U3897 ( .A1(i_data_bus[519]), .A2(n4052), .B1(
        i_data_bus[551]), .B2(n4047), .ZN(n3523) );
  AOI22D1BWP30P140LVT U3898 ( .A1(i_data_bus[615]), .A2(n4049), .B1(
        i_data_bus[583]), .B2(n4050), .ZN(n3522) );
  AOI22D1BWP30P140LVT U3899 ( .A1(i_data_bus[999]), .A2(n3383), .B1(
        i_data_bus[935]), .B2(n4051), .ZN(n3521) );
  INVD1BWP30P140LVT U3900 ( .I(i_data_bus[359]), .ZN(n4912) );
  MOAI22D1BWP30P140LVT U3901 ( .A1(n4912), .A2(n3983), .B1(i_data_bus[295]), 
        .B2(n3347), .ZN(n3537) );
  MOAI22D1BWP30P140LVT U3902 ( .A1(n3525), .A2(n3984), .B1(i_data_bus[327]), 
        .B2(n3348), .ZN(n3536) );
  AOI22D1BWP30P140LVT U3903 ( .A1(i_data_bus[743]), .A2(n3353), .B1(
        i_data_bus[167]), .B2(n4037), .ZN(n3529) );
  AOI22D1BWP30P140LVT U3904 ( .A1(i_data_bus[679]), .A2(n4035), .B1(
        i_data_bus[647]), .B2(n4040), .ZN(n3528) );
  AOI22D1BWP30P140LVT U3905 ( .A1(i_data_bus[71]), .A2(n4028), .B1(
        i_data_bus[231]), .B2(n3352), .ZN(n3527) );
  AOI22D1BWP30P140LVT U3906 ( .A1(i_data_bus[39]), .A2(n4025), .B1(
        i_data_bus[7]), .B2(n4038), .ZN(n3526) );
  ND4D1BWP30P140LVT U3907 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), 
        .ZN(n3535) );
  AOI22D1BWP30P140LVT U3908 ( .A1(i_data_bus[839]), .A2(n4036), .B1(
        i_data_bus[775]), .B2(n4027), .ZN(n3533) );
  AOI22D1BWP30P140LVT U3909 ( .A1(i_data_bus[135]), .A2(n3355), .B1(
        i_data_bus[199]), .B2(n3351), .ZN(n3532) );
  AOI22D1BWP30P140LVT U3910 ( .A1(i_data_bus[871]), .A2(n4039), .B1(
        i_data_bus[711]), .B2(n3360), .ZN(n3531) );
  AOI22D1BWP30P140LVT U3911 ( .A1(i_data_bus[103]), .A2(n4026), .B1(
        i_data_bus[807]), .B2(n4024), .ZN(n3530) );
  ND4D1BWP30P140LVT U3912 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), 
        .ZN(n3534) );
  NR4D0BWP30P140LVT U3913 ( .A1(n3537), .A2(n3536), .A3(n3535), .A4(n3534), 
        .ZN(n3538) );
  ND4D1BWP30P140LVT U3914 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), 
        .ZN(o_data_bus[71]) );
  AOI22D1BWP30P140LVT U3915 ( .A1(i_data_bus[488]), .A2(n4020), .B1(
        i_data_bus[360]), .B2(n4033), .ZN(n3561) );
  AOI22D1BWP30P140LVT U3916 ( .A1(i_data_bus[264]), .A2(n4023), .B1(
        i_data_bus[424]), .B2(n4021), .ZN(n3560) );
  AOI22D1BWP30P140LVT U3917 ( .A1(i_data_bus[840]), .A2(n4036), .B1(
        i_data_bus[776]), .B2(n4027), .ZN(n3545) );
  AOI22D1BWP30P140LVT U3918 ( .A1(i_data_bus[72]), .A2(n4028), .B1(
        i_data_bus[744]), .B2(n3353), .ZN(n3544) );
  AOI22D1BWP30P140LVT U3919 ( .A1(i_data_bus[808]), .A2(n4024), .B1(
        i_data_bus[648]), .B2(n4040), .ZN(n3543) );
  AOI22D1BWP30P140LVT U3920 ( .A1(i_data_bus[680]), .A2(n4035), .B1(
        i_data_bus[136]), .B2(n3355), .ZN(n3542) );
  AOI22D1BWP30P140LVT U3921 ( .A1(i_data_bus[456]), .A2(n4006), .B1(
        i_data_bus[328]), .B2(n3348), .ZN(n3557) );
  AOI22D1BWP30P140LVT U3922 ( .A1(i_data_bus[872]), .A2(n4039), .B1(
        i_data_bus[232]), .B2(n3352), .ZN(n3549) );
  AOI22D1BWP30P140LVT U3923 ( .A1(i_data_bus[8]), .A2(n4038), .B1(
        i_data_bus[200]), .B2(n3351), .ZN(n3548) );
  AOI22D1BWP30P140LVT U3924 ( .A1(i_data_bus[40]), .A2(n4025), .B1(
        i_data_bus[712]), .B2(n3360), .ZN(n3547) );
  AOI22D1BWP30P140LVT U3925 ( .A1(i_data_bus[104]), .A2(n4026), .B1(
        i_data_bus[168]), .B2(n4037), .ZN(n3546) );
  ND4D1BWP30P140LVT U3926 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), 
        .ZN(n3556) );
  INVD1BWP30P140LVT U3927 ( .I(i_data_bus[296]), .ZN(n5663) );
  MOAI22D1BWP30P140LVT U3928 ( .A1(n5663), .A2(n3878), .B1(i_data_bus[392]), 
        .B2(n4022), .ZN(n3555) );
  AOI22D1BWP30P140LVT U3929 ( .A1(i_data_bus[1000]), .A2(n3383), .B1(
        i_data_bus[584]), .B2(n4050), .ZN(n3553) );
  AOI22D1BWP30P140LVT U3930 ( .A1(i_data_bus[616]), .A2(n4049), .B1(
        i_data_bus[520]), .B2(n4052), .ZN(n3552) );
  AOI22D1BWP30P140LVT U3931 ( .A1(i_data_bus[968]), .A2(n4048), .B1(
        i_data_bus[936]), .B2(n4051), .ZN(n3551) );
  AOI22D1BWP30P140LVT U3932 ( .A1(i_data_bus[552]), .A2(n4047), .B1(
        i_data_bus[904]), .B2(n3378), .ZN(n3550) );
  ND4D1BWP30P140LVT U3933 ( .A1(n3553), .A2(n3552), .A3(n3551), .A4(n3550), 
        .ZN(n3554) );
  INR4D0BWP30P140LVT U3934 ( .A1(n3557), .B1(n3556), .B2(n3555), .B3(n3554), 
        .ZN(n3558) );
  ND4D1BWP30P140LVT U3935 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), 
        .ZN(o_data_bus[72]) );
  AOI22D1BWP30P140LVT U3936 ( .A1(i_data_bus[489]), .A2(n4020), .B1(
        i_data_bus[329]), .B2(n3348), .ZN(n3582) );
  AOI22D1BWP30P140LVT U3937 ( .A1(i_data_bus[265]), .A2(n4023), .B1(
        i_data_bus[457]), .B2(n4006), .ZN(n3581) );
  AOI22D1BWP30P140LVT U3938 ( .A1(i_data_bus[41]), .A2(n4025), .B1(
        i_data_bus[745]), .B2(n3353), .ZN(n3565) );
  AOI22D1BWP30P140LVT U3939 ( .A1(i_data_bus[73]), .A2(n4028), .B1(
        i_data_bus[841]), .B2(n4036), .ZN(n3564) );
  AOI22D1BWP30P140LVT U3940 ( .A1(i_data_bus[873]), .A2(n4039), .B1(
        i_data_bus[809]), .B2(n4024), .ZN(n3563) );
  AOI22D1BWP30P140LVT U3941 ( .A1(i_data_bus[681]), .A2(n4035), .B1(
        i_data_bus[777]), .B2(n4027), .ZN(n3562) );
  AOI22D1BWP30P140LVT U3942 ( .A1(i_data_bus[425]), .A2(n4021), .B1(
        i_data_bus[361]), .B2(n4033), .ZN(n3578) );
  AOI22D1BWP30P140LVT U3943 ( .A1(i_data_bus[201]), .A2(n3351), .B1(
        i_data_bus[233]), .B2(n3352), .ZN(n3569) );
  AOI22D1BWP30P140LVT U3944 ( .A1(i_data_bus[169]), .A2(n4037), .B1(
        i_data_bus[649]), .B2(n4040), .ZN(n3568) );
  AOI22D1BWP30P140LVT U3945 ( .A1(i_data_bus[9]), .A2(n4038), .B1(
        i_data_bus[137]), .B2(n3355), .ZN(n3567) );
  AOI22D1BWP30P140LVT U3946 ( .A1(i_data_bus[105]), .A2(n4026), .B1(
        i_data_bus[713]), .B2(n3360), .ZN(n3566) );
  ND4D1BWP30P140LVT U3947 ( .A1(n3569), .A2(n3568), .A3(n3567), .A4(n3566), 
        .ZN(n3577) );
  INVD1BWP30P140LVT U3948 ( .I(i_data_bus[297]), .ZN(n5684) );
  OAI22D1BWP30P140LVT U3949 ( .A1(n5684), .A2(n3878), .B1(n3570), .B2(n4007), 
        .ZN(n3576) );
  AOI22D1BWP30P140LVT U3950 ( .A1(i_data_bus[585]), .A2(n4050), .B1(
        i_data_bus[617]), .B2(n4049), .ZN(n3574) );
  AOI22D1BWP30P140LVT U3951 ( .A1(i_data_bus[521]), .A2(n4052), .B1(
        i_data_bus[969]), .B2(n4048), .ZN(n3573) );
  AOI22D1BWP30P140LVT U3952 ( .A1(i_data_bus[1001]), .A2(n3383), .B1(
        i_data_bus[937]), .B2(n4051), .ZN(n3572) );
  AOI22D1BWP30P140LVT U3953 ( .A1(i_data_bus[905]), .A2(n3378), .B1(
        i_data_bus[553]), .B2(n4047), .ZN(n3571) );
  ND4D1BWP30P140LVT U3954 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), 
        .ZN(n3575) );
  INR4D0BWP30P140LVT U3955 ( .A1(n3578), .B1(n3577), .B2(n3576), .B3(n3575), 
        .ZN(n3579) );
  ND4D1BWP30P140LVT U3956 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), 
        .ZN(o_data_bus[73]) );
  AOI22D1BWP30P140LVT U3957 ( .A1(i_data_bus[298]), .A2(n3347), .B1(
        i_data_bus[426]), .B2(n4021), .ZN(n3602) );
  AOI22D1BWP30P140LVT U3958 ( .A1(i_data_bus[458]), .A2(n4006), .B1(
        i_data_bus[266]), .B2(n4023), .ZN(n3601) );
  AOI22D1BWP30P140LVT U3959 ( .A1(i_data_bus[234]), .A2(n3352), .B1(
        i_data_bus[874]), .B2(n4039), .ZN(n3586) );
  AOI22D1BWP30P140LVT U3960 ( .A1(i_data_bus[106]), .A2(n4026), .B1(
        i_data_bus[170]), .B2(n4037), .ZN(n3585) );
  AOI22D1BWP30P140LVT U3961 ( .A1(i_data_bus[714]), .A2(n3360), .B1(
        i_data_bus[682]), .B2(n4035), .ZN(n3583) );
  AOI22D1BWP30P140LVT U3962 ( .A1(i_data_bus[650]), .A2(n4040), .B1(
        i_data_bus[746]), .B2(n3353), .ZN(n3590) );
  AOI22D1BWP30P140LVT U3963 ( .A1(i_data_bus[10]), .A2(n4038), .B1(
        i_data_bus[778]), .B2(n4027), .ZN(n3589) );
  AOI22D1BWP30P140LVT U3964 ( .A1(i_data_bus[202]), .A2(n3351), .B1(
        i_data_bus[810]), .B2(n4024), .ZN(n3588) );
  AOI22D1BWP30P140LVT U3965 ( .A1(i_data_bus[842]), .A2(n4036), .B1(
        i_data_bus[138]), .B2(n3355), .ZN(n3587) );
  ND4D1BWP30P140LVT U3966 ( .A1(n3590), .A2(n3589), .A3(n3588), .A4(n3587), 
        .ZN(n3598) );
  INVD1BWP30P140LVT U3967 ( .I(i_data_bus[490]), .ZN(n5706) );
  MOAI22D1BWP30P140LVT U3968 ( .A1(n5706), .A2(n3984), .B1(i_data_bus[362]), 
        .B2(n4033), .ZN(n3597) );
  MOAI22D1BWP30P140LVT U3969 ( .A1(n5705), .A2(n4007), .B1(i_data_bus[330]), 
        .B2(n3348), .ZN(n3596) );
  AOI22D1BWP30P140LVT U3970 ( .A1(i_data_bus[970]), .A2(n4048), .B1(
        i_data_bus[522]), .B2(n4052), .ZN(n3594) );
  AOI22D1BWP30P140LVT U3971 ( .A1(i_data_bus[618]), .A2(n4049), .B1(
        i_data_bus[938]), .B2(n4051), .ZN(n3593) );
  AOI22D1BWP30P140LVT U3972 ( .A1(i_data_bus[554]), .A2(n4047), .B1(
        i_data_bus[586]), .B2(n4050), .ZN(n3592) );
  AOI22D1BWP30P140LVT U3973 ( .A1(i_data_bus[1002]), .A2(n3383), .B1(
        i_data_bus[906]), .B2(n3378), .ZN(n3591) );
  ND4D1BWP30P140LVT U3974 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), 
        .ZN(n3595) );
  NR4D0BWP30P140LVT U3975 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), 
        .ZN(n3599) );
  ND4D1BWP30P140LVT U3976 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), 
        .ZN(o_data_bus[74]) );
  AOI22D1BWP30P140LVT U3977 ( .A1(i_data_bus[491]), .A2(n4020), .B1(
        i_data_bus[427]), .B2(n4021), .ZN(n3622) );
  AOI22D1BWP30P140LVT U3978 ( .A1(i_data_bus[363]), .A2(n4033), .B1(
        i_data_bus[299]), .B2(n3347), .ZN(n3621) );
  AOI22D1BWP30P140LVT U3979 ( .A1(i_data_bus[139]), .A2(n3355), .B1(
        i_data_bus[683]), .B2(n4035), .ZN(n3606) );
  AOI22D1BWP30P140LVT U3980 ( .A1(i_data_bus[75]), .A2(n4028), .B1(
        i_data_bus[171]), .B2(n4037), .ZN(n3605) );
  AOI22D1BWP30P140LVT U3981 ( .A1(i_data_bus[747]), .A2(n3353), .B1(
        i_data_bus[779]), .B2(n4027), .ZN(n3604) );
  AOI22D1BWP30P140LVT U3982 ( .A1(i_data_bus[11]), .A2(n4038), .B1(
        i_data_bus[107]), .B2(n4026), .ZN(n3603) );
  AOI22D1BWP30P140LVT U3983 ( .A1(i_data_bus[395]), .A2(n4022), .B1(
        i_data_bus[267]), .B2(n4023), .ZN(n3618) );
  AOI22D1BWP30P140LVT U3984 ( .A1(i_data_bus[651]), .A2(n4040), .B1(
        i_data_bus[715]), .B2(n3360), .ZN(n3610) );
  AOI22D1BWP30P140LVT U3985 ( .A1(i_data_bus[203]), .A2(n3351), .B1(
        i_data_bus[875]), .B2(n4039), .ZN(n3609) );
  AOI22D1BWP30P140LVT U3986 ( .A1(i_data_bus[43]), .A2(n4025), .B1(
        i_data_bus[811]), .B2(n4024), .ZN(n3608) );
  AOI22D1BWP30P140LVT U3987 ( .A1(i_data_bus[843]), .A2(n4036), .B1(
        i_data_bus[235]), .B2(n3352), .ZN(n3607) );
  ND4D1BWP30P140LVT U3988 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), 
        .ZN(n3617) );
  INVD1BWP30P140LVT U3989 ( .I(i_data_bus[331]), .ZN(n5727) );
  OAI22D1BWP30P140LVT U3990 ( .A1(n5729), .A2(n4046), .B1(n5727), .B2(n3961), 
        .ZN(n3616) );
  AOI22D1BWP30P140LVT U3991 ( .A1(i_data_bus[907]), .A2(n3378), .B1(
        i_data_bus[619]), .B2(n4049), .ZN(n3614) );
  AOI22D1BWP30P140LVT U3992 ( .A1(i_data_bus[523]), .A2(n4052), .B1(
        i_data_bus[555]), .B2(n4047), .ZN(n3613) );
  AOI22D1BWP30P140LVT U3993 ( .A1(i_data_bus[1003]), .A2(n3383), .B1(
        i_data_bus[587]), .B2(n4050), .ZN(n3612) );
  AOI22D1BWP30P140LVT U3994 ( .A1(i_data_bus[939]), .A2(n4051), .B1(
        i_data_bus[971]), .B2(n4048), .ZN(n3611) );
  ND4D1BWP30P140LVT U3995 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), 
        .ZN(n3615) );
  INR4D0BWP30P140LVT U3996 ( .A1(n3618), .B1(n3617), .B2(n3616), .B3(n3615), 
        .ZN(n3619) );
  ND4D1BWP30P140LVT U3997 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), 
        .ZN(o_data_bus[75]) );
  AOI22D1BWP30P140LVT U3998 ( .A1(i_data_bus[268]), .A2(n4023), .B1(
        i_data_bus[332]), .B2(n3348), .ZN(n3642) );
  AOI22D1BWP30P140LVT U3999 ( .A1(i_data_bus[300]), .A2(n3347), .B1(
        i_data_bus[396]), .B2(n4022), .ZN(n3641) );
  AOI22D1BWP30P140LVT U4000 ( .A1(i_data_bus[76]), .A2(n4028), .B1(
        i_data_bus[844]), .B2(n4036), .ZN(n3626) );
  AOI22D1BWP30P140LVT U4001 ( .A1(i_data_bus[716]), .A2(n3360), .B1(
        i_data_bus[204]), .B2(n3351), .ZN(n3625) );
  AOI22D1BWP30P140LVT U4002 ( .A1(i_data_bus[684]), .A2(n4035), .B1(
        i_data_bus[236]), .B2(n3352), .ZN(n3624) );
  AOI22D1BWP30P140LVT U4003 ( .A1(i_data_bus[12]), .A2(n4038), .B1(
        i_data_bus[172]), .B2(n4037), .ZN(n3623) );
  AOI22D1BWP30P140LVT U4004 ( .A1(i_data_bus[364]), .A2(n4033), .B1(
        i_data_bus[428]), .B2(n4021), .ZN(n3638) );
  AOI22D1BWP30P140LVT U4005 ( .A1(i_data_bus[44]), .A2(n4025), .B1(
        i_data_bus[108]), .B2(n4026), .ZN(n3630) );
  AOI22D1BWP30P140LVT U4006 ( .A1(i_data_bus[812]), .A2(n4024), .B1(
        i_data_bus[876]), .B2(n4039), .ZN(n3629) );
  AOI22D1BWP30P140LVT U4007 ( .A1(i_data_bus[780]), .A2(n4027), .B1(
        i_data_bus[748]), .B2(n3353), .ZN(n3628) );
  AOI22D1BWP30P140LVT U4008 ( .A1(i_data_bus[140]), .A2(n3355), .B1(
        i_data_bus[652]), .B2(n4040), .ZN(n3627) );
  ND4D1BWP30P140LVT U4009 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), 
        .ZN(n3637) );
  INVD1BWP30P140LVT U4010 ( .I(i_data_bus[460]), .ZN(n5015) );
  OAI22D1BWP30P140LVT U4011 ( .A1(n5015), .A2(n4046), .B1(n5014), .B2(n3984), 
        .ZN(n3636) );
  AOI22D1BWP30P140LVT U4012 ( .A1(i_data_bus[940]), .A2(n4051), .B1(
        i_data_bus[972]), .B2(n4048), .ZN(n3634) );
  AOI22D1BWP30P140LVT U4013 ( .A1(i_data_bus[620]), .A2(n4049), .B1(
        i_data_bus[588]), .B2(n4050), .ZN(n3633) );
  AOI22D1BWP30P140LVT U4014 ( .A1(i_data_bus[908]), .A2(n3378), .B1(
        i_data_bus[1004]), .B2(n3383), .ZN(n3632) );
  AOI22D1BWP30P140LVT U4015 ( .A1(i_data_bus[556]), .A2(n4047), .B1(
        i_data_bus[524]), .B2(n4052), .ZN(n3631) );
  ND4D1BWP30P140LVT U4016 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), 
        .ZN(n3635) );
  INR4D0BWP30P140LVT U4017 ( .A1(n3638), .B1(n3637), .B2(n3636), .B3(n3635), 
        .ZN(n3639) );
  ND4D1BWP30P140LVT U4018 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), 
        .ZN(o_data_bus[76]) );
  AOI22D1BWP30P140LVT U4019 ( .A1(i_data_bus[365]), .A2(n4033), .B1(
        i_data_bus[461]), .B2(n4006), .ZN(n3662) );
  AOI22D1BWP30P140LVT U4020 ( .A1(i_data_bus[429]), .A2(n4021), .B1(
        i_data_bus[333]), .B2(n3348), .ZN(n3661) );
  AOI22D1BWP30P140LVT U4021 ( .A1(i_data_bus[525]), .A2(n4052), .B1(
        i_data_bus[621]), .B2(n4049), .ZN(n3646) );
  AOI22D1BWP30P140LVT U4022 ( .A1(i_data_bus[973]), .A2(n4048), .B1(
        i_data_bus[941]), .B2(n4051), .ZN(n3645) );
  AOI22D1BWP30P140LVT U4023 ( .A1(i_data_bus[557]), .A2(n4047), .B1(
        i_data_bus[1005]), .B2(n3383), .ZN(n3644) );
  AOI22D1BWP30P140LVT U4024 ( .A1(i_data_bus[909]), .A2(n3378), .B1(
        i_data_bus[589]), .B2(n4050), .ZN(n3643) );
  AOI22D1BWP30P140LVT U4025 ( .A1(i_data_bus[397]), .A2(n4022), .B1(
        i_data_bus[269]), .B2(n4023), .ZN(n3658) );
  MOAI22D1BWP30P140LVT U4026 ( .A1(n5036), .A2(n3984), .B1(i_data_bus[301]), 
        .B2(n3347), .ZN(n3657) );
  AOI22D1BWP30P140LVT U4027 ( .A1(i_data_bus[749]), .A2(n3353), .B1(
        i_data_bus[173]), .B2(n4037), .ZN(n3650) );
  AOI22D1BWP30P140LVT U4028 ( .A1(i_data_bus[77]), .A2(n4028), .B1(
        i_data_bus[141]), .B2(n3355), .ZN(n3649) );
  AOI22D1BWP30P140LVT U4029 ( .A1(i_data_bus[45]), .A2(n4025), .B1(
        i_data_bus[813]), .B2(n4024), .ZN(n3648) );
  AOI22D1BWP30P140LVT U4030 ( .A1(i_data_bus[781]), .A2(n4027), .B1(
        i_data_bus[205]), .B2(n3351), .ZN(n3647) );
  ND4D1BWP30P140LVT U4031 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), 
        .ZN(n3656) );
  AOI22D1BWP30P140LVT U4032 ( .A1(i_data_bus[685]), .A2(n4035), .B1(
        i_data_bus[717]), .B2(n3360), .ZN(n3654) );
  AOI22D1BWP30P140LVT U4033 ( .A1(i_data_bus[109]), .A2(n4026), .B1(
        i_data_bus[653]), .B2(n4040), .ZN(n3653) );
  AOI22D1BWP30P140LVT U4034 ( .A1(i_data_bus[13]), .A2(n4038), .B1(
        i_data_bus[877]), .B2(n4039), .ZN(n3652) );
  AOI22D1BWP30P140LVT U4035 ( .A1(i_data_bus[237]), .A2(n3352), .B1(
        i_data_bus[845]), .B2(n4036), .ZN(n3651) );
  ND4D1BWP30P140LVT U4036 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), 
        .ZN(n3655) );
  INR4D0BWP30P140LVT U4037 ( .A1(n3658), .B1(n3657), .B2(n3656), .B3(n3655), 
        .ZN(n3659) );
  ND4D1BWP30P140LVT U4038 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), 
        .ZN(o_data_bus[77]) );
  AOI22D1BWP30P140LVT U4039 ( .A1(i_data_bus[462]), .A2(n4006), .B1(
        i_data_bus[334]), .B2(n3348), .ZN(n3683) );
  AOI22D1BWP30P140LVT U4040 ( .A1(i_data_bus[270]), .A2(n4023), .B1(
        i_data_bus[302]), .B2(n3347), .ZN(n3682) );
  AOI22D1BWP30P140LVT U4041 ( .A1(i_data_bus[206]), .A2(n3351), .B1(
        i_data_bus[814]), .B2(n4024), .ZN(n3666) );
  AOI22D1BWP30P140LVT U4042 ( .A1(i_data_bus[238]), .A2(n3352), .B1(
        i_data_bus[654]), .B2(n4040), .ZN(n3665) );
  AOI22D1BWP30P140LVT U4043 ( .A1(i_data_bus[46]), .A2(n4025), .B1(
        i_data_bus[782]), .B2(n4027), .ZN(n3664) );
  AOI22D1BWP30P140LVT U4044 ( .A1(i_data_bus[14]), .A2(n4038), .B1(
        i_data_bus[718]), .B2(n3360), .ZN(n3663) );
  AOI22D1BWP30P140LVT U4045 ( .A1(i_data_bus[110]), .A2(n4026), .B1(
        i_data_bus[174]), .B2(n4037), .ZN(n3670) );
  AOI22D1BWP30P140LVT U4046 ( .A1(i_data_bus[78]), .A2(n4028), .B1(
        i_data_bus[750]), .B2(n3353), .ZN(n3669) );
  AOI22D1BWP30P140LVT U4047 ( .A1(i_data_bus[142]), .A2(n3355), .B1(
        i_data_bus[846]), .B2(n4036), .ZN(n3668) );
  AOI22D1BWP30P140LVT U4048 ( .A1(i_data_bus[878]), .A2(n4039), .B1(
        i_data_bus[686]), .B2(n4035), .ZN(n3667) );
  ND4D1BWP30P140LVT U4049 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), 
        .ZN(n3679) );
  MOAI22D1BWP30P140LVT U4050 ( .A1(n3671), .A2(n4007), .B1(i_data_bus[430]), 
        .B2(n4021), .ZN(n3678) );
  INVD1BWP30P140LVT U4051 ( .I(i_data_bus[494]), .ZN(n5792) );
  MOAI22D1BWP30P140LVT U4052 ( .A1(n5792), .A2(n3984), .B1(i_data_bus[366]), 
        .B2(n4033), .ZN(n3677) );
  AOI22D1BWP30P140LVT U4053 ( .A1(i_data_bus[974]), .A2(n4048), .B1(
        i_data_bus[942]), .B2(n4051), .ZN(n3675) );
  AOI22D1BWP30P140LVT U4054 ( .A1(i_data_bus[1006]), .A2(n3383), .B1(
        i_data_bus[558]), .B2(n4047), .ZN(n3674) );
  AOI22D1BWP30P140LVT U4055 ( .A1(i_data_bus[910]), .A2(n3378), .B1(
        i_data_bus[590]), .B2(n4050), .ZN(n3673) );
  AOI22D1BWP30P140LVT U4056 ( .A1(i_data_bus[622]), .A2(n4049), .B1(
        i_data_bus[526]), .B2(n4052), .ZN(n3672) );
  ND4D1BWP30P140LVT U4057 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), 
        .ZN(n3676) );
  NR4D0BWP30P140LVT U4058 ( .A1(n3679), .A2(n3678), .A3(n3677), .A4(n3676), 
        .ZN(n3680) );
  ND4D1BWP30P140LVT U4059 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), 
        .ZN(o_data_bus[78]) );
  AOI22D1BWP30P140LVT U4060 ( .A1(i_data_bus[271]), .A2(n4023), .B1(
        i_data_bus[303]), .B2(n3347), .ZN(n3704) );
  AOI22D1BWP30P140LVT U4061 ( .A1(i_data_bus[431]), .A2(n4021), .B1(
        i_data_bus[335]), .B2(n3348), .ZN(n3703) );
  AOI22D1BWP30P140LVT U4062 ( .A1(i_data_bus[911]), .A2(n3378), .B1(
        i_data_bus[623]), .B2(n4049), .ZN(n3687) );
  AOI22D1BWP30P140LVT U4063 ( .A1(i_data_bus[975]), .A2(n4048), .B1(
        i_data_bus[527]), .B2(n4052), .ZN(n3686) );
  AOI22D1BWP30P140LVT U4064 ( .A1(i_data_bus[1007]), .A2(n3383), .B1(
        i_data_bus[943]), .B2(n4051), .ZN(n3685) );
  AOI22D1BWP30P140LVT U4065 ( .A1(i_data_bus[591]), .A2(n4050), .B1(
        i_data_bus[559]), .B2(n4047), .ZN(n3684) );
  MOAI22D1BWP30P140LVT U4066 ( .A1(n3688), .A2(n4046), .B1(i_data_bus[495]), 
        .B2(n4020), .ZN(n3700) );
  INVD1BWP30P140LVT U4067 ( .I(i_data_bus[399]), .ZN(n5077) );
  INVD1BWP30P140LVT U4068 ( .I(i_data_bus[367]), .ZN(n5813) );
  OAI22D1BWP30P140LVT U4069 ( .A1(n5077), .A2(n4007), .B1(n5813), .B2(n3983), 
        .ZN(n3699) );
  AOI22D1BWP30P140LVT U4070 ( .A1(i_data_bus[143]), .A2(n3355), .B1(
        i_data_bus[655]), .B2(n4040), .ZN(n3692) );
  AOI22D1BWP30P140LVT U4071 ( .A1(i_data_bus[47]), .A2(n4025), .B1(
        i_data_bus[687]), .B2(n4035), .ZN(n3691) );
  AOI22D1BWP30P140LVT U4072 ( .A1(i_data_bus[15]), .A2(n4038), .B1(
        i_data_bus[239]), .B2(n3352), .ZN(n3690) );
  AOI22D1BWP30P140LVT U4073 ( .A1(i_data_bus[207]), .A2(n3351), .B1(
        i_data_bus[879]), .B2(n4039), .ZN(n3689) );
  ND4D1BWP30P140LVT U4074 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), 
        .ZN(n3698) );
  AOI22D1BWP30P140LVT U4075 ( .A1(i_data_bus[79]), .A2(n4028), .B1(
        i_data_bus[175]), .B2(n4037), .ZN(n3696) );
  AOI22D1BWP30P140LVT U4076 ( .A1(i_data_bus[719]), .A2(n3360), .B1(
        i_data_bus[783]), .B2(n4027), .ZN(n3695) );
  AOI22D1BWP30P140LVT U4077 ( .A1(i_data_bus[111]), .A2(n4026), .B1(
        i_data_bus[751]), .B2(n3353), .ZN(n3694) );
  AOI22D1BWP30P140LVT U4078 ( .A1(i_data_bus[847]), .A2(n4036), .B1(
        i_data_bus[815]), .B2(n4024), .ZN(n3693) );
  ND4D1BWP30P140LVT U4079 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), 
        .ZN(n3697) );
  NR4D0BWP30P140LVT U4080 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), 
        .ZN(n3701) );
  ND4D1BWP30P140LVT U4081 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), 
        .ZN(o_data_bus[79]) );
  AOI22D1BWP30P140LVT U4082 ( .A1(i_data_bus[304]), .A2(n3347), .B1(
        i_data_bus[368]), .B2(n4033), .ZN(n3725) );
  AOI22D1BWP30P140LVT U4083 ( .A1(i_data_bus[336]), .A2(n3348), .B1(
        i_data_bus[464]), .B2(n4006), .ZN(n3724) );
  AOI22D1BWP30P140LVT U4084 ( .A1(i_data_bus[528]), .A2(n4052), .B1(
        i_data_bus[912]), .B2(n3378), .ZN(n3708) );
  AOI22D1BWP30P140LVT U4085 ( .A1(i_data_bus[624]), .A2(n4049), .B1(
        i_data_bus[976]), .B2(n4048), .ZN(n3707) );
  AOI22D1BWP30P140LVT U4086 ( .A1(i_data_bus[944]), .A2(n4051), .B1(
        i_data_bus[592]), .B2(n4050), .ZN(n3706) );
  AOI22D1BWP30P140LVT U4087 ( .A1(i_data_bus[560]), .A2(n4047), .B1(
        i_data_bus[1008]), .B2(n3383), .ZN(n3705) );
  MOAI22D1BWP30P140LVT U4088 ( .A1(n3709), .A2(n3984), .B1(i_data_bus[272]), 
        .B2(n4023), .ZN(n3721) );
  INVD1BWP30P140LVT U4089 ( .I(i_data_bus[400]), .ZN(n5834) );
  MOAI22D1BWP30P140LVT U4090 ( .A1(n5834), .A2(n4007), .B1(i_data_bus[432]), 
        .B2(n4021), .ZN(n3720) );
  AOI22D1BWP30P140LVT U4091 ( .A1(i_data_bus[16]), .A2(n4038), .B1(
        i_data_bus[144]), .B2(n3355), .ZN(n3713) );
  AOI22D1BWP30P140LVT U4092 ( .A1(i_data_bus[752]), .A2(n3353), .B1(
        i_data_bus[816]), .B2(n4024), .ZN(n3712) );
  AOI22D1BWP30P140LVT U4093 ( .A1(i_data_bus[784]), .A2(n4027), .B1(
        i_data_bus[656]), .B2(n4040), .ZN(n3711) );
  AOI22D1BWP30P140LVT U4094 ( .A1(i_data_bus[880]), .A2(n4039), .B1(
        i_data_bus[688]), .B2(n4035), .ZN(n3710) );
  ND4D1BWP30P140LVT U4095 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), 
        .ZN(n3719) );
  AOI22D1BWP30P140LVT U4096 ( .A1(i_data_bus[80]), .A2(n4028), .B1(
        i_data_bus[848]), .B2(n4036), .ZN(n3717) );
  AOI22D1BWP30P140LVT U4097 ( .A1(i_data_bus[112]), .A2(n4026), .B1(
        i_data_bus[176]), .B2(n4037), .ZN(n3716) );
  AOI22D1BWP30P140LVT U4098 ( .A1(i_data_bus[48]), .A2(n4025), .B1(
        i_data_bus[720]), .B2(n3360), .ZN(n3715) );
  AOI22D1BWP30P140LVT U4099 ( .A1(i_data_bus[208]), .A2(n3351), .B1(
        i_data_bus[240]), .B2(n3352), .ZN(n3714) );
  ND4D1BWP30P140LVT U4100 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), 
        .ZN(n3718) );
  NR4D0BWP30P140LVT U4101 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), 
        .ZN(n3722) );
  ND4D1BWP30P140LVT U4102 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), 
        .ZN(o_data_bus[80]) );
  AOI22D1BWP30P140LVT U4103 ( .A1(i_data_bus[433]), .A2(n4021), .B1(
        i_data_bus[401]), .B2(n4022), .ZN(n3745) );
  AOI22D1BWP30P140LVT U4104 ( .A1(i_data_bus[465]), .A2(n4006), .B1(
        i_data_bus[497]), .B2(n4020), .ZN(n3744) );
  AOI22D1BWP30P140LVT U4105 ( .A1(i_data_bus[881]), .A2(n4039), .B1(
        i_data_bus[145]), .B2(n3355), .ZN(n3729) );
  AOI22D1BWP30P140LVT U4106 ( .A1(i_data_bus[657]), .A2(n4040), .B1(
        i_data_bus[753]), .B2(n3353), .ZN(n3728) );
  AOI22D1BWP30P140LVT U4107 ( .A1(i_data_bus[849]), .A2(n4036), .B1(
        i_data_bus[817]), .B2(n4024), .ZN(n3727) );
  AOI22D1BWP30P140LVT U4108 ( .A1(i_data_bus[785]), .A2(n4027), .B1(
        i_data_bus[721]), .B2(n3360), .ZN(n3726) );
  AOI22D1BWP30P140LVT U4109 ( .A1(i_data_bus[337]), .A2(n3348), .B1(
        i_data_bus[273]), .B2(n4023), .ZN(n3741) );
  AOI22D1BWP30P140LVT U4110 ( .A1(i_data_bus[17]), .A2(n4038), .B1(
        i_data_bus[49]), .B2(n4025), .ZN(n3733) );
  AOI22D1BWP30P140LVT U4111 ( .A1(i_data_bus[241]), .A2(n3352), .B1(
        i_data_bus[209]), .B2(n3351), .ZN(n3732) );
  AOI22D1BWP30P140LVT U4112 ( .A1(i_data_bus[81]), .A2(n4028), .B1(
        i_data_bus[689]), .B2(n4035), .ZN(n3731) );
  AOI22D1BWP30P140LVT U4113 ( .A1(i_data_bus[113]), .A2(n4026), .B1(
        i_data_bus[177]), .B2(n4037), .ZN(n3730) );
  ND4D1BWP30P140LVT U4114 ( .A1(n3733), .A2(n3732), .A3(n3731), .A4(n3730), 
        .ZN(n3740) );
  INVD1BWP30P140LVT U4115 ( .I(i_data_bus[369]), .ZN(n5855) );
  MOAI22D1BWP30P140LVT U4116 ( .A1(n5855), .A2(n3983), .B1(i_data_bus[305]), 
        .B2(n3347), .ZN(n3739) );
  AOI22D1BWP30P140LVT U4117 ( .A1(i_data_bus[625]), .A2(n4049), .B1(
        i_data_bus[1009]), .B2(n3383), .ZN(n3737) );
  AOI22D1BWP30P140LVT U4118 ( .A1(i_data_bus[593]), .A2(n4050), .B1(
        i_data_bus[529]), .B2(n4052), .ZN(n3736) );
  AOI22D1BWP30P140LVT U4119 ( .A1(i_data_bus[945]), .A2(n4051), .B1(
        i_data_bus[977]), .B2(n4048), .ZN(n3735) );
  AOI22D1BWP30P140LVT U4120 ( .A1(i_data_bus[913]), .A2(n3378), .B1(
        i_data_bus[561]), .B2(n4047), .ZN(n3734) );
  ND4D1BWP30P140LVT U4121 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), 
        .ZN(n3738) );
  INR4D0BWP30P140LVT U4122 ( .A1(n3741), .B1(n3740), .B2(n3739), .B3(n3738), 
        .ZN(n3742) );
  ND4D1BWP30P140LVT U4123 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), 
        .ZN(o_data_bus[81]) );
  AOI22D1BWP30P140LVT U4124 ( .A1(i_data_bus[498]), .A2(n4020), .B1(
        i_data_bus[306]), .B2(n3347), .ZN(n3765) );
  AOI22D1BWP30P140LVT U4125 ( .A1(i_data_bus[274]), .A2(n4023), .B1(
        i_data_bus[434]), .B2(n4021), .ZN(n3764) );
  AOI22D1BWP30P140LVT U4126 ( .A1(i_data_bus[18]), .A2(n4038), .B1(
        i_data_bus[690]), .B2(n4035), .ZN(n3749) );
  AOI22D1BWP30P140LVT U4127 ( .A1(i_data_bus[50]), .A2(n4025), .B1(
        i_data_bus[850]), .B2(n4036), .ZN(n3748) );
  AOI22D1BWP30P140LVT U4128 ( .A1(i_data_bus[82]), .A2(n4028), .B1(
        i_data_bus[754]), .B2(n3353), .ZN(n3747) );
  AOI22D1BWP30P140LVT U4129 ( .A1(i_data_bus[146]), .A2(n3355), .B1(
        i_data_bus[786]), .B2(n4027), .ZN(n3746) );
  AOI22D1BWP30P140LVT U4130 ( .A1(i_data_bus[402]), .A2(n4022), .B1(
        i_data_bus[370]), .B2(n4033), .ZN(n3761) );
  AO22D1BWP30P140LVT U4131 ( .A1(i_data_bus[466]), .A2(n4006), .B1(
        i_data_bus[338]), .B2(n3348), .Z(n3760) );
  AOI22D1BWP30P140LVT U4132 ( .A1(i_data_bus[242]), .A2(n3352), .B1(
        i_data_bus[178]), .B2(n4037), .ZN(n3753) );
  AOI22D1BWP30P140LVT U4133 ( .A1(i_data_bus[722]), .A2(n3360), .B1(
        i_data_bus[210]), .B2(n3351), .ZN(n3752) );
  AOI22D1BWP30P140LVT U4134 ( .A1(i_data_bus[818]), .A2(n4024), .B1(
        i_data_bus[658]), .B2(n4040), .ZN(n3751) );
  AOI22D1BWP30P140LVT U4135 ( .A1(i_data_bus[114]), .A2(n4026), .B1(
        i_data_bus[882]), .B2(n4039), .ZN(n3750) );
  ND4D1BWP30P140LVT U4136 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), 
        .ZN(n3759) );
  AOI22D1BWP30P140LVT U4137 ( .A1(i_data_bus[594]), .A2(n4050), .B1(
        i_data_bus[530]), .B2(n4052), .ZN(n3757) );
  AOI22D1BWP30P140LVT U4138 ( .A1(i_data_bus[562]), .A2(n4047), .B1(
        i_data_bus[946]), .B2(n4051), .ZN(n3756) );
  AOI22D1BWP30P140LVT U4139 ( .A1(i_data_bus[626]), .A2(n4049), .B1(
        i_data_bus[978]), .B2(n4048), .ZN(n3755) );
  AOI22D1BWP30P140LVT U4140 ( .A1(i_data_bus[1010]), .A2(n3383), .B1(
        i_data_bus[914]), .B2(n3378), .ZN(n3754) );
  ND4D1BWP30P140LVT U4141 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), 
        .ZN(n3758) );
  INR4D0BWP30P140LVT U4142 ( .A1(n3761), .B1(n3760), .B2(n3759), .B3(n3758), 
        .ZN(n3762) );
  ND4D1BWP30P140LVT U4143 ( .A1(n3765), .A2(n3764), .A3(n3763), .A4(n3762), 
        .ZN(o_data_bus[82]) );
  AOI22D1BWP30P140LVT U4144 ( .A1(i_data_bus[339]), .A2(n3348), .B1(
        i_data_bus[435]), .B2(n4021), .ZN(n3785) );
  AOI22D1BWP30P140LVT U4145 ( .A1(i_data_bus[371]), .A2(n4033), .B1(
        i_data_bus[403]), .B2(n4022), .ZN(n3784) );
  AOI22D1BWP30P140LVT U4146 ( .A1(i_data_bus[243]), .A2(n3352), .B1(
        i_data_bus[659]), .B2(n4040), .ZN(n3769) );
  AOI22D1BWP30P140LVT U4147 ( .A1(i_data_bus[19]), .A2(n4038), .B1(
        i_data_bus[883]), .B2(n4039), .ZN(n3768) );
  AOI22D1BWP30P140LVT U4148 ( .A1(i_data_bus[179]), .A2(n4037), .B1(
        i_data_bus[851]), .B2(n4036), .ZN(n3767) );
  AOI22D1BWP30P140LVT U4149 ( .A1(i_data_bus[211]), .A2(n3351), .B1(
        i_data_bus[787]), .B2(n4027), .ZN(n3766) );
  AOI22D1BWP30P140LVT U4150 ( .A1(i_data_bus[83]), .A2(n4028), .B1(
        i_data_bus[691]), .B2(n4035), .ZN(n3773) );
  AOI22D1BWP30P140LVT U4151 ( .A1(i_data_bus[115]), .A2(n4026), .B1(
        i_data_bus[755]), .B2(n3353), .ZN(n3772) );
  AOI22D1BWP30P140LVT U4152 ( .A1(i_data_bus[147]), .A2(n3355), .B1(
        i_data_bus[819]), .B2(n4024), .ZN(n3771) );
  AOI22D1BWP30P140LVT U4153 ( .A1(i_data_bus[51]), .A2(n4025), .B1(
        i_data_bus[723]), .B2(n3360), .ZN(n3770) );
  ND4D1BWP30P140LVT U4154 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), 
        .ZN(n3781) );
  INVD1BWP30P140LVT U4155 ( .I(i_data_bus[499]), .ZN(n5899) );
  MOAI22D1BWP30P140LVT U4156 ( .A1(n5899), .A2(n3984), .B1(i_data_bus[275]), 
        .B2(n4023), .ZN(n3780) );
  INVD1BWP30P140LVT U4157 ( .I(i_data_bus[307]), .ZN(n5158) );
  MOAI22D1BWP30P140LVT U4158 ( .A1(n5158), .A2(n3878), .B1(i_data_bus[467]), 
        .B2(n4006), .ZN(n3779) );
  AOI22D1BWP30P140LVT U4159 ( .A1(i_data_bus[627]), .A2(n4049), .B1(
        i_data_bus[595]), .B2(n4050), .ZN(n3777) );
  AOI22D1BWP30P140LVT U4160 ( .A1(i_data_bus[531]), .A2(n4052), .B1(
        i_data_bus[947]), .B2(n4051), .ZN(n3776) );
  AOI22D1BWP30P140LVT U4161 ( .A1(i_data_bus[979]), .A2(n4048), .B1(
        i_data_bus[1011]), .B2(n3383), .ZN(n3775) );
  AOI22D1BWP30P140LVT U4162 ( .A1(i_data_bus[563]), .A2(n4047), .B1(
        i_data_bus[915]), .B2(n3378), .ZN(n3774) );
  ND4D1BWP30P140LVT U4163 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), 
        .ZN(n3778) );
  NR4D0BWP30P140LVT U4164 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), 
        .ZN(n3782) );
  ND4D1BWP30P140LVT U4165 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), 
        .ZN(o_data_bus[83]) );
  AOI22D1BWP30P140LVT U4166 ( .A1(i_data_bus[404]), .A2(n4022), .B1(
        i_data_bus[500]), .B2(n4020), .ZN(n3806) );
  AOI22D1BWP30P140LVT U4167 ( .A1(i_data_bus[340]), .A2(n3348), .B1(
        i_data_bus[276]), .B2(n4023), .ZN(n3805) );
  AOI22D1BWP30P140LVT U4168 ( .A1(i_data_bus[948]), .A2(n4051), .B1(
        i_data_bus[916]), .B2(n3378), .ZN(n3789) );
  AOI22D1BWP30P140LVT U4169 ( .A1(i_data_bus[1012]), .A2(n3383), .B1(
        i_data_bus[564]), .B2(n4047), .ZN(n3788) );
  AOI22D1BWP30P140LVT U4170 ( .A1(i_data_bus[596]), .A2(n4050), .B1(
        i_data_bus[532]), .B2(n4052), .ZN(n3787) );
  AOI22D1BWP30P140LVT U4171 ( .A1(i_data_bus[980]), .A2(n4048), .B1(
        i_data_bus[628]), .B2(n4049), .ZN(n3786) );
  MOAI22D1BWP30P140LVT U4172 ( .A1(n3790), .A2(n4046), .B1(i_data_bus[372]), 
        .B2(n4033), .ZN(n3802) );
  INVD1BWP30P140LVT U4173 ( .I(i_data_bus[308]), .ZN(n5921) );
  MOAI22D1BWP30P140LVT U4174 ( .A1(n5921), .A2(n3878), .B1(i_data_bus[436]), 
        .B2(n4021), .ZN(n3801) );
  AOI22D1BWP30P140LVT U4175 ( .A1(i_data_bus[212]), .A2(n3351), .B1(
        i_data_bus[180]), .B2(n4037), .ZN(n3794) );
  AOI22D1BWP30P140LVT U4176 ( .A1(i_data_bus[52]), .A2(n4025), .B1(
        i_data_bus[788]), .B2(n4027), .ZN(n3793) );
  AOI22D1BWP30P140LVT U4177 ( .A1(i_data_bus[852]), .A2(n4036), .B1(
        i_data_bus[148]), .B2(n3355), .ZN(n3792) );
  AOI22D1BWP30P140LVT U4178 ( .A1(i_data_bus[884]), .A2(n4039), .B1(
        i_data_bus[660]), .B2(n4040), .ZN(n3791) );
  ND4D1BWP30P140LVT U4179 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), 
        .ZN(n3800) );
  AOI22D1BWP30P140LVT U4180 ( .A1(i_data_bus[20]), .A2(n4038), .B1(
        i_data_bus[724]), .B2(n3360), .ZN(n3798) );
  AOI22D1BWP30P140LVT U4181 ( .A1(i_data_bus[244]), .A2(n3352), .B1(
        i_data_bus[756]), .B2(n3353), .ZN(n3797) );
  AOI22D1BWP30P140LVT U4182 ( .A1(i_data_bus[116]), .A2(n4026), .B1(
        i_data_bus[820]), .B2(n4024), .ZN(n3796) );
  AOI22D1BWP30P140LVT U4183 ( .A1(i_data_bus[84]), .A2(n4028), .B1(
        i_data_bus[692]), .B2(n4035), .ZN(n3795) );
  ND4D1BWP30P140LVT U4184 ( .A1(n3795), .A2(n3797), .A3(n3796), .A4(n3798), 
        .ZN(n3799) );
  NR4D0BWP30P140LVT U4185 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), 
        .ZN(n3803) );
  ND4D1BWP30P140LVT U4186 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), 
        .ZN(o_data_bus[84]) );
  AOI22D1BWP30P140LVT U4187 ( .A1(i_data_bus[437]), .A2(n4021), .B1(
        i_data_bus[501]), .B2(n4020), .ZN(n3827) );
  AOI22D1BWP30P140LVT U4188 ( .A1(i_data_bus[341]), .A2(n3348), .B1(
        i_data_bus[277]), .B2(n4023), .ZN(n3826) );
  AOI22D1BWP30P140LVT U4189 ( .A1(i_data_bus[981]), .A2(n4048), .B1(
        i_data_bus[1013]), .B2(n3383), .ZN(n3810) );
  AOI22D1BWP30P140LVT U4190 ( .A1(i_data_bus[949]), .A2(n4051), .B1(
        i_data_bus[917]), .B2(n3378), .ZN(n3809) );
  AOI22D1BWP30P140LVT U4191 ( .A1(i_data_bus[629]), .A2(n4049), .B1(
        i_data_bus[565]), .B2(n4047), .ZN(n3808) );
  AOI22D1BWP30P140LVT U4192 ( .A1(i_data_bus[597]), .A2(n4050), .B1(
        i_data_bus[533]), .B2(n4052), .ZN(n3807) );
  INVD1BWP30P140LVT U4193 ( .I(i_data_bus[373]), .ZN(n5942) );
  MOAI22D1BWP30P140LVT U4194 ( .A1(n5942), .A2(n3983), .B1(i_data_bus[469]), 
        .B2(n4006), .ZN(n3823) );
  INVD1BWP30P140LVT U4195 ( .I(i_data_bus[309]), .ZN(n5199) );
  OAI22D1BWP30P140LVT U4196 ( .A1(n5199), .A2(n3878), .B1(n3811), .B2(n4007), 
        .ZN(n3822) );
  AOI22D1BWP30P140LVT U4197 ( .A1(i_data_bus[821]), .A2(n4024), .B1(
        i_data_bus[725]), .B2(n3360), .ZN(n3815) );
  AOI22D1BWP30P140LVT U4198 ( .A1(i_data_bus[181]), .A2(n4037), .B1(
        i_data_bus[213]), .B2(n3351), .ZN(n3814) );
  AOI22D1BWP30P140LVT U4199 ( .A1(i_data_bus[21]), .A2(n4038), .B1(
        i_data_bus[149]), .B2(n3355), .ZN(n3813) );
  AOI22D1BWP30P140LVT U4200 ( .A1(i_data_bus[853]), .A2(n4036), .B1(
        i_data_bus[789]), .B2(n4027), .ZN(n3812) );
  ND4D1BWP30P140LVT U4201 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), 
        .ZN(n3821) );
  AOI22D1BWP30P140LVT U4202 ( .A1(i_data_bus[117]), .A2(n4026), .B1(
        i_data_bus[693]), .B2(n4035), .ZN(n3819) );
  AOI22D1BWP30P140LVT U4203 ( .A1(i_data_bus[757]), .A2(n3353), .B1(
        i_data_bus[885]), .B2(n4039), .ZN(n3818) );
  AOI22D1BWP30P140LVT U4204 ( .A1(i_data_bus[85]), .A2(n4028), .B1(
        i_data_bus[661]), .B2(n4040), .ZN(n3817) );
  AOI22D1BWP30P140LVT U4205 ( .A1(i_data_bus[53]), .A2(n4025), .B1(
        i_data_bus[245]), .B2(n3352), .ZN(n3816) );
  ND4D1BWP30P140LVT U4206 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), 
        .ZN(n3820) );
  NR4D0BWP30P140LVT U4207 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), 
        .ZN(n3824) );
  ND4D1BWP30P140LVT U4208 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), 
        .ZN(o_data_bus[85]) );
  AOI22D1BWP30P140LVT U4209 ( .A1(i_data_bus[438]), .A2(n4021), .B1(
        i_data_bus[502]), .B2(n4020), .ZN(n3847) );
  AOI22D1BWP30P140LVT U4210 ( .A1(i_data_bus[310]), .A2(n3347), .B1(
        i_data_bus[278]), .B2(n4023), .ZN(n3846) );
  AOI22D1BWP30P140LVT U4211 ( .A1(i_data_bus[822]), .A2(n4024), .B1(
        i_data_bus[246]), .B2(n3352), .ZN(n3831) );
  AOI22D1BWP30P140LVT U4212 ( .A1(i_data_bus[758]), .A2(n3353), .B1(
        i_data_bus[886]), .B2(n4039), .ZN(n3829) );
  AOI22D1BWP30P140LVT U4213 ( .A1(i_data_bus[182]), .A2(n4037), .B1(
        i_data_bus[214]), .B2(n3351), .ZN(n3828) );
  AOI22D1BWP30P140LVT U4214 ( .A1(i_data_bus[22]), .A2(n4038), .B1(
        i_data_bus[662]), .B2(n4040), .ZN(n3835) );
  AOI22D1BWP30P140LVT U4215 ( .A1(i_data_bus[54]), .A2(n4025), .B1(
        i_data_bus[150]), .B2(n3355), .ZN(n3834) );
  AOI22D1BWP30P140LVT U4216 ( .A1(i_data_bus[694]), .A2(n4035), .B1(
        i_data_bus[726]), .B2(n3360), .ZN(n3833) );
  AOI22D1BWP30P140LVT U4217 ( .A1(i_data_bus[790]), .A2(n4027), .B1(
        i_data_bus[854]), .B2(n4036), .ZN(n3832) );
  ND4D1BWP30P140LVT U4218 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), 
        .ZN(n3843) );
  MOAI22D1BWP30P140LVT U4219 ( .A1(n5222), .A2(n4046), .B1(i_data_bus[374]), 
        .B2(n4033), .ZN(n3842) );
  INVD1BWP30P140LVT U4220 ( .I(i_data_bus[342]), .ZN(n5221) );
  MOAI22D1BWP30P140LVT U4221 ( .A1(n5221), .A2(n3961), .B1(i_data_bus[406]), 
        .B2(n4022), .ZN(n3841) );
  AOI22D1BWP30P140LVT U4222 ( .A1(i_data_bus[534]), .A2(n4052), .B1(
        i_data_bus[918]), .B2(n3378), .ZN(n3839) );
  AOI22D1BWP30P140LVT U4223 ( .A1(i_data_bus[566]), .A2(n4047), .B1(
        i_data_bus[982]), .B2(n4048), .ZN(n3838) );
  AOI22D1BWP30P140LVT U4224 ( .A1(i_data_bus[1014]), .A2(n3383), .B1(
        i_data_bus[598]), .B2(n4050), .ZN(n3837) );
  AOI22D1BWP30P140LVT U4225 ( .A1(i_data_bus[950]), .A2(n4051), .B1(
        i_data_bus[630]), .B2(n4049), .ZN(n3836) );
  ND4D1BWP30P140LVT U4226 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), 
        .ZN(n3840) );
  NR4D0BWP30P140LVT U4227 ( .A1(n3843), .A2(n3842), .A3(n3841), .A4(n3840), 
        .ZN(n3844) );
  ND4D1BWP30P140LVT U4228 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), 
        .ZN(o_data_bus[86]) );
  AOI22D1BWP30P140LVT U4229 ( .A1(i_data_bus[503]), .A2(n4020), .B1(
        i_data_bus[343]), .B2(n3348), .ZN(n3868) );
  AOI22D1BWP30P140LVT U4230 ( .A1(i_data_bus[311]), .A2(n3347), .B1(
        i_data_bus[407]), .B2(n4022), .ZN(n3867) );
  AOI22D1BWP30P140LVT U4231 ( .A1(i_data_bus[183]), .A2(n4037), .B1(
        i_data_bus[151]), .B2(n3355), .ZN(n3851) );
  AOI22D1BWP30P140LVT U4232 ( .A1(i_data_bus[55]), .A2(n4025), .B1(
        i_data_bus[727]), .B2(n3360), .ZN(n3850) );
  AOI22D1BWP30P140LVT U4233 ( .A1(i_data_bus[759]), .A2(n3353), .B1(
        i_data_bus[663]), .B2(n4040), .ZN(n3849) );
  AOI22D1BWP30P140LVT U4234 ( .A1(i_data_bus[23]), .A2(n4038), .B1(
        i_data_bus[823]), .B2(n4024), .ZN(n3848) );
  AOI22D1BWP30P140LVT U4235 ( .A1(i_data_bus[87]), .A2(n4028), .B1(
        i_data_bus[119]), .B2(n4026), .ZN(n3855) );
  AOI22D1BWP30P140LVT U4236 ( .A1(i_data_bus[695]), .A2(n4035), .B1(
        i_data_bus[791]), .B2(n4027), .ZN(n3854) );
  AOI22D1BWP30P140LVT U4237 ( .A1(i_data_bus[247]), .A2(n3352), .B1(
        i_data_bus[215]), .B2(n3351), .ZN(n3853) );
  AOI22D1BWP30P140LVT U4238 ( .A1(i_data_bus[887]), .A2(n4039), .B1(
        i_data_bus[855]), .B2(n4036), .ZN(n3852) );
  ND4D1BWP30P140LVT U4239 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), 
        .ZN(n3864) );
  INVD1BWP30P140LVT U4240 ( .I(i_data_bus[375]), .ZN(n5985) );
  OAI22D1BWP30P140LVT U4241 ( .A1(n5243), .A2(n4046), .B1(n5985), .B2(n3983), 
        .ZN(n3863) );
  INVD1BWP30P140LVT U4242 ( .I(i_data_bus[439]), .ZN(n5987) );
  MOAI22D1BWP30P140LVT U4243 ( .A1(n5987), .A2(n3856), .B1(i_data_bus[279]), 
        .B2(n4023), .ZN(n3862) );
  AOI22D1BWP30P140LVT U4244 ( .A1(i_data_bus[1015]), .A2(n3383), .B1(
        i_data_bus[567]), .B2(n4047), .ZN(n3860) );
  AOI22D1BWP30P140LVT U4245 ( .A1(i_data_bus[631]), .A2(n4049), .B1(
        i_data_bus[919]), .B2(n3378), .ZN(n3859) );
  AOI22D1BWP30P140LVT U4246 ( .A1(i_data_bus[983]), .A2(n4048), .B1(
        i_data_bus[535]), .B2(n4052), .ZN(n3858) );
  AOI22D1BWP30P140LVT U4247 ( .A1(i_data_bus[599]), .A2(n4050), .B1(
        i_data_bus[951]), .B2(n4051), .ZN(n3857) );
  ND4D1BWP30P140LVT U4248 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), 
        .ZN(n3861) );
  NR4D0BWP30P140LVT U4249 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), 
        .ZN(n3865) );
  ND4D1BWP30P140LVT U4250 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), 
        .ZN(o_data_bus[87]) );
  AOI22D1BWP30P140LVT U4251 ( .A1(i_data_bus[344]), .A2(n3348), .B1(
        i_data_bus[408]), .B2(n4022), .ZN(n3890) );
  AOI22D1BWP30P140LVT U4252 ( .A1(i_data_bus[440]), .A2(n4021), .B1(
        i_data_bus[472]), .B2(n4006), .ZN(n3889) );
  AOI22D1BWP30P140LVT U4253 ( .A1(i_data_bus[696]), .A2(n4035), .B1(
        i_data_bus[760]), .B2(n3353), .ZN(n3872) );
  AOI22D1BWP30P140LVT U4254 ( .A1(i_data_bus[248]), .A2(n3352), .B1(
        i_data_bus[888]), .B2(n4039), .ZN(n3871) );
  AOI22D1BWP30P140LVT U4255 ( .A1(i_data_bus[88]), .A2(n4028), .B1(
        i_data_bus[216]), .B2(n3351), .ZN(n3870) );
  AOI22D1BWP30P140LVT U4256 ( .A1(i_data_bus[824]), .A2(n4024), .B1(
        i_data_bus[184]), .B2(n4037), .ZN(n3869) );
  AOI22D1BWP30P140LVT U4257 ( .A1(i_data_bus[24]), .A2(n4038), .B1(
        i_data_bus[728]), .B2(n3360), .ZN(n3876) );
  AOI22D1BWP30P140LVT U4258 ( .A1(i_data_bus[856]), .A2(n4036), .B1(
        i_data_bus[664]), .B2(n4040), .ZN(n3875) );
  AOI22D1BWP30P140LVT U4259 ( .A1(i_data_bus[120]), .A2(n4026), .B1(
        i_data_bus[56]), .B2(n4025), .ZN(n3874) );
  AOI22D1BWP30P140LVT U4260 ( .A1(i_data_bus[792]), .A2(n4027), .B1(
        i_data_bus[152]), .B2(n3355), .ZN(n3873) );
  ND4D1BWP30P140LVT U4261 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), 
        .ZN(n3886) );
  MOAI22D1BWP30P140LVT U4262 ( .A1(n3877), .A2(n3984), .B1(i_data_bus[376]), 
        .B2(n4033), .ZN(n3885) );
  INVD1BWP30P140LVT U4263 ( .I(i_data_bus[280]), .ZN(n6008) );
  INVD1BWP30P140LVT U4264 ( .I(i_data_bus[312]), .ZN(n5265) );
  OAI22D1BWP30P140LVT U4265 ( .A1(n6008), .A2(n3982), .B1(n5265), .B2(n3878), 
        .ZN(n3884) );
  AOI22D1BWP30P140LVT U4266 ( .A1(i_data_bus[984]), .A2(n4048), .B1(
        i_data_bus[568]), .B2(n4047), .ZN(n3882) );
  AOI22D1BWP30P140LVT U4267 ( .A1(i_data_bus[1016]), .A2(n3383), .B1(
        i_data_bus[920]), .B2(n3378), .ZN(n3881) );
  AOI22D1BWP30P140LVT U4268 ( .A1(i_data_bus[632]), .A2(n4049), .B1(
        i_data_bus[536]), .B2(n4052), .ZN(n3880) );
  AOI22D1BWP30P140LVT U4269 ( .A1(i_data_bus[600]), .A2(n4050), .B1(
        i_data_bus[952]), .B2(n4051), .ZN(n3879) );
  ND4D1BWP30P140LVT U4270 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), 
        .ZN(n3883) );
  NR4D0BWP30P140LVT U4271 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), 
        .ZN(n3887) );
  ND4D1BWP30P140LVT U4272 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), 
        .ZN(o_data_bus[88]) );
  AOI22D1BWP30P140LVT U4273 ( .A1(i_data_bus[377]), .A2(n4033), .B1(
        i_data_bus[473]), .B2(n4006), .ZN(n3910) );
  AOI22D1BWP30P140LVT U4274 ( .A1(i_data_bus[345]), .A2(n3348), .B1(
        i_data_bus[313]), .B2(n3347), .ZN(n3909) );
  AOI22D1BWP30P140LVT U4275 ( .A1(i_data_bus[921]), .A2(n3378), .B1(
        i_data_bus[985]), .B2(n4048), .ZN(n3894) );
  AOI22D1BWP30P140LVT U4276 ( .A1(i_data_bus[537]), .A2(n4052), .B1(
        i_data_bus[953]), .B2(n4051), .ZN(n3893) );
  AOI22D1BWP30P140LVT U4277 ( .A1(i_data_bus[1017]), .A2(n3383), .B1(
        i_data_bus[633]), .B2(n4049), .ZN(n3892) );
  AOI22D1BWP30P140LVT U4278 ( .A1(i_data_bus[569]), .A2(n4047), .B1(
        i_data_bus[601]), .B2(n4050), .ZN(n3891) );
  MOAI22D1BWP30P140LVT U4279 ( .A1(n6029), .A2(n4007), .B1(i_data_bus[281]), 
        .B2(n4023), .ZN(n3906) );
  MOAI22D1BWP30P140LVT U4280 ( .A1(n5286), .A2(n3984), .B1(i_data_bus[441]), 
        .B2(n4021), .ZN(n3905) );
  AOI22D1BWP30P140LVT U4281 ( .A1(i_data_bus[121]), .A2(n4026), .B1(
        i_data_bus[249]), .B2(n3352), .ZN(n3898) );
  AOI22D1BWP30P140LVT U4282 ( .A1(i_data_bus[57]), .A2(n4025), .B1(
        i_data_bus[857]), .B2(n4036), .ZN(n3897) );
  AOI22D1BWP30P140LVT U4283 ( .A1(i_data_bus[153]), .A2(n3355), .B1(
        i_data_bus[889]), .B2(n4039), .ZN(n3896) );
  AOI22D1BWP30P140LVT U4284 ( .A1(i_data_bus[89]), .A2(n4028), .B1(
        i_data_bus[217]), .B2(n3351), .ZN(n3895) );
  ND4D1BWP30P140LVT U4285 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), 
        .ZN(n3904) );
  AOI22D1BWP30P140LVT U4286 ( .A1(i_data_bus[729]), .A2(n3360), .B1(
        i_data_bus[793]), .B2(n4027), .ZN(n3902) );
  AOI22D1BWP30P140LVT U4287 ( .A1(i_data_bus[697]), .A2(n4035), .B1(
        i_data_bus[185]), .B2(n4037), .ZN(n3901) );
  AOI22D1BWP30P140LVT U4288 ( .A1(i_data_bus[25]), .A2(n4038), .B1(
        i_data_bus[825]), .B2(n4024), .ZN(n3900) );
  AOI22D1BWP30P140LVT U4289 ( .A1(i_data_bus[665]), .A2(n4040), .B1(
        i_data_bus[761]), .B2(n3353), .ZN(n3899) );
  ND4D1BWP30P140LVT U4290 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), 
        .ZN(n3903) );
  NR4D0BWP30P140LVT U4291 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), 
        .ZN(n3907) );
  ND4D1BWP30P140LVT U4292 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), 
        .ZN(o_data_bus[89]) );
  AOI22D1BWP30P140LVT U4293 ( .A1(i_data_bus[442]), .A2(n4021), .B1(
        i_data_bus[282]), .B2(n4023), .ZN(n3930) );
  AOI22D1BWP30P140LVT U4294 ( .A1(i_data_bus[314]), .A2(n3347), .B1(
        i_data_bus[346]), .B2(n3348), .ZN(n3929) );
  AOI22D1BWP30P140LVT U4295 ( .A1(i_data_bus[250]), .A2(n3352), .B1(
        i_data_bus[666]), .B2(n4040), .ZN(n3914) );
  AOI22D1BWP30P140LVT U4296 ( .A1(i_data_bus[826]), .A2(n4024), .B1(
        i_data_bus[186]), .B2(n4037), .ZN(n3913) );
  AOI22D1BWP30P140LVT U4297 ( .A1(i_data_bus[218]), .A2(n3351), .B1(
        i_data_bus[858]), .B2(n4036), .ZN(n3912) );
  AOI22D1BWP30P140LVT U4298 ( .A1(i_data_bus[698]), .A2(n4035), .B1(
        i_data_bus[762]), .B2(n3353), .ZN(n3911) );
  AOI22D1BWP30P140LVT U4299 ( .A1(i_data_bus[58]), .A2(n4025), .B1(
        i_data_bus[794]), .B2(n4027), .ZN(n3918) );
  AOI22D1BWP30P140LVT U4300 ( .A1(i_data_bus[26]), .A2(n4038), .B1(
        i_data_bus[154]), .B2(n3355), .ZN(n3917) );
  AOI22D1BWP30P140LVT U4301 ( .A1(i_data_bus[122]), .A2(n4026), .B1(
        i_data_bus[90]), .B2(n4028), .ZN(n3916) );
  AOI22D1BWP30P140LVT U4302 ( .A1(i_data_bus[890]), .A2(n4039), .B1(
        i_data_bus[730]), .B2(n3360), .ZN(n3915) );
  ND4D1BWP30P140LVT U4303 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), 
        .ZN(n3926) );
  INVD1BWP30P140LVT U4304 ( .I(i_data_bus[378]), .ZN(n6050) );
  MOAI22D1BWP30P140LVT U4305 ( .A1(n6050), .A2(n3983), .B1(i_data_bus[474]), 
        .B2(n4006), .ZN(n3925) );
  INVD1BWP30P140LVT U4306 ( .I(i_data_bus[506]), .ZN(n5309) );
  OAI22D1BWP30P140LVT U4307 ( .A1(n5309), .A2(n3984), .B1(n5307), .B2(n4007), 
        .ZN(n3924) );
  AOI22D1BWP30P140LVT U4308 ( .A1(i_data_bus[602]), .A2(n4050), .B1(
        i_data_bus[954]), .B2(n4051), .ZN(n3922) );
  AOI22D1BWP30P140LVT U4309 ( .A1(i_data_bus[986]), .A2(n4048), .B1(
        i_data_bus[922]), .B2(n3378), .ZN(n3921) );
  AOI22D1BWP30P140LVT U4310 ( .A1(i_data_bus[1018]), .A2(n3383), .B1(
        i_data_bus[570]), .B2(n4047), .ZN(n3920) );
  AOI22D1BWP30P140LVT U4311 ( .A1(i_data_bus[538]), .A2(n4052), .B1(
        i_data_bus[634]), .B2(n4049), .ZN(n3919) );
  ND4D1BWP30P140LVT U4312 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), 
        .ZN(n3923) );
  NR4D0BWP30P140LVT U4313 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), 
        .ZN(n3927) );
  AOI22D1BWP30P140LVT U4314 ( .A1(i_data_bus[315]), .A2(n3347), .B1(
        i_data_bus[475]), .B2(n4006), .ZN(n3951) );
  AOI22D1BWP30P140LVT U4315 ( .A1(i_data_bus[443]), .A2(n4021), .B1(
        i_data_bus[283]), .B2(n4023), .ZN(n3950) );
  AOI22D1BWP30P140LVT U4316 ( .A1(i_data_bus[891]), .A2(n4039), .B1(
        i_data_bus[859]), .B2(n4036), .ZN(n3934) );
  AOI22D1BWP30P140LVT U4317 ( .A1(i_data_bus[59]), .A2(n4025), .B1(
        i_data_bus[763]), .B2(n3353), .ZN(n3933) );
  AOI22D1BWP30P140LVT U4318 ( .A1(i_data_bus[219]), .A2(n3351), .B1(
        i_data_bus[187]), .B2(n4037), .ZN(n3932) );
  AOI22D1BWP30P140LVT U4319 ( .A1(i_data_bus[667]), .A2(n4040), .B1(
        i_data_bus[699]), .B2(n4035), .ZN(n3931) );
  AOI22D1BWP30P140LVT U4320 ( .A1(i_data_bus[123]), .A2(n4026), .B1(
        i_data_bus[795]), .B2(n4027), .ZN(n3938) );
  AOI22D1BWP30P140LVT U4321 ( .A1(i_data_bus[27]), .A2(n4038), .B1(
        i_data_bus[731]), .B2(n3360), .ZN(n3937) );
  AOI22D1BWP30P140LVT U4322 ( .A1(i_data_bus[91]), .A2(n4028), .B1(
        i_data_bus[251]), .B2(n3352), .ZN(n3936) );
  AOI22D1BWP30P140LVT U4323 ( .A1(i_data_bus[827]), .A2(n4024), .B1(
        i_data_bus[155]), .B2(n3355), .ZN(n3935) );
  ND4D1BWP30P140LVT U4324 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), 
        .ZN(n3947) );
  MOAI22D1BWP30P140LVT U4325 ( .A1(n3939), .A2(n3983), .B1(i_data_bus[507]), 
        .B2(n4020), .ZN(n3946) );
  INVD1BWP30P140LVT U4326 ( .I(i_data_bus[347]), .ZN(n6072) );
  MOAI22D1BWP30P140LVT U4327 ( .A1(n6072), .A2(n3961), .B1(i_data_bus[411]), 
        .B2(n4022), .ZN(n3945) );
  AOI22D1BWP30P140LVT U4328 ( .A1(i_data_bus[571]), .A2(n4047), .B1(
        i_data_bus[539]), .B2(n4052), .ZN(n3943) );
  AOI22D1BWP30P140LVT U4329 ( .A1(i_data_bus[987]), .A2(n4048), .B1(
        i_data_bus[603]), .B2(n4050), .ZN(n3942) );
  AOI22D1BWP30P140LVT U4330 ( .A1(i_data_bus[635]), .A2(n4049), .B1(
        i_data_bus[923]), .B2(n3378), .ZN(n3941) );
  AOI22D1BWP30P140LVT U4331 ( .A1(i_data_bus[1019]), .A2(n3383), .B1(
        i_data_bus[955]), .B2(n4051), .ZN(n3940) );
  ND4D1BWP30P140LVT U4332 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), 
        .ZN(n3944) );
  NR4D0BWP30P140LVT U4333 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), 
        .ZN(n3948) );
  ND4D1BWP30P140LVT U4334 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), 
        .ZN(o_data_bus[91]) );
  AOI22D1BWP30P140LVT U4335 ( .A1(i_data_bus[380]), .A2(n4033), .B1(
        i_data_bus[444]), .B2(n4021), .ZN(n3973) );
  AOI22D1BWP30P140LVT U4336 ( .A1(i_data_bus[508]), .A2(n4020), .B1(
        i_data_bus[316]), .B2(n3347), .ZN(n3972) );
  AOI22D1BWP30P140LVT U4337 ( .A1(i_data_bus[92]), .A2(n4028), .B1(
        i_data_bus[892]), .B2(n4039), .ZN(n3955) );
  AOI22D1BWP30P140LVT U4338 ( .A1(i_data_bus[764]), .A2(n3353), .B1(
        i_data_bus[860]), .B2(n4036), .ZN(n3954) );
  AOI22D1BWP30P140LVT U4339 ( .A1(i_data_bus[124]), .A2(n4026), .B1(
        i_data_bus[700]), .B2(n4035), .ZN(n3953) );
  AOI22D1BWP30P140LVT U4340 ( .A1(i_data_bus[796]), .A2(n4027), .B1(
        i_data_bus[156]), .B2(n3355), .ZN(n3952) );
  AOI22D1BWP30P140LVT U4341 ( .A1(i_data_bus[60]), .A2(n4025), .B1(
        i_data_bus[252]), .B2(n3352), .ZN(n3959) );
  AOI22D1BWP30P140LVT U4342 ( .A1(i_data_bus[28]), .A2(n4038), .B1(
        i_data_bus[668]), .B2(n4040), .ZN(n3958) );
  AOI22D1BWP30P140LVT U4343 ( .A1(i_data_bus[828]), .A2(n4024), .B1(
        i_data_bus[220]), .B2(n3351), .ZN(n3957) );
  AOI22D1BWP30P140LVT U4344 ( .A1(i_data_bus[732]), .A2(n3360), .B1(
        i_data_bus[188]), .B2(n4037), .ZN(n3956) );
  ND4D1BWP30P140LVT U4345 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), 
        .ZN(n3969) );
  INVD1BWP30P140LVT U4346 ( .I(i_data_bus[284]), .ZN(n5330) );
  OAI22D1BWP30P140LVT U4347 ( .A1(n3960), .A2(n4046), .B1(n5330), .B2(n3982), 
        .ZN(n3968) );
  INVD1BWP30P140LVT U4348 ( .I(i_data_bus[348]), .ZN(n6095) );
  INVD1BWP30P140LVT U4349 ( .I(i_data_bus[412]), .ZN(n6093) );
  AOI22D1BWP30P140LVT U4350 ( .A1(i_data_bus[988]), .A2(n4048), .B1(
        i_data_bus[956]), .B2(n4051), .ZN(n3965) );
  AOI22D1BWP30P140LVT U4351 ( .A1(i_data_bus[540]), .A2(n4052), .B1(
        i_data_bus[604]), .B2(n4050), .ZN(n3964) );
  AOI22D1BWP30P140LVT U4352 ( .A1(i_data_bus[924]), .A2(n3378), .B1(
        i_data_bus[1020]), .B2(n3383), .ZN(n3963) );
  AOI22D1BWP30P140LVT U4353 ( .A1(i_data_bus[636]), .A2(n4049), .B1(
        i_data_bus[572]), .B2(n4047), .ZN(n3962) );
  ND4D1BWP30P140LVT U4354 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), 
        .ZN(n3966) );
  NR4D0BWP30P140LVT U4355 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), 
        .ZN(n3970) );
  ND4D1BWP30P140LVT U4356 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), 
        .ZN(o_data_bus[92]) );
  AOI22D1BWP30P140LVT U4357 ( .A1(i_data_bus[445]), .A2(n4021), .B1(
        i_data_bus[413]), .B2(n4022), .ZN(n3997) );
  AOI22D1BWP30P140LVT U4358 ( .A1(i_data_bus[349]), .A2(n3348), .B1(
        i_data_bus[477]), .B2(n4006), .ZN(n3996) );
  AOI22D1BWP30P140LVT U4359 ( .A1(i_data_bus[765]), .A2(n3353), .B1(
        i_data_bus[733]), .B2(n3360), .ZN(n3977) );
  AOI22D1BWP30P140LVT U4360 ( .A1(i_data_bus[29]), .A2(n4038), .B1(
        i_data_bus[61]), .B2(n4025), .ZN(n3976) );
  AOI22D1BWP30P140LVT U4361 ( .A1(i_data_bus[701]), .A2(n4035), .B1(
        i_data_bus[669]), .B2(n4040), .ZN(n3975) );
  AOI22D1BWP30P140LVT U4362 ( .A1(i_data_bus[861]), .A2(n4036), .B1(
        i_data_bus[221]), .B2(n3351), .ZN(n3974) );
  AOI22D1BWP30P140LVT U4363 ( .A1(i_data_bus[125]), .A2(n4026), .B1(
        i_data_bus[893]), .B2(n4039), .ZN(n3981) );
  AOI22D1BWP30P140LVT U4364 ( .A1(i_data_bus[93]), .A2(n4028), .B1(
        i_data_bus[797]), .B2(n4027), .ZN(n3980) );
  AOI22D1BWP30P140LVT U4365 ( .A1(i_data_bus[189]), .A2(n4037), .B1(
        i_data_bus[253]), .B2(n3352), .ZN(n3979) );
  AOI22D1BWP30P140LVT U4366 ( .A1(i_data_bus[157]), .A2(n3355), .B1(
        i_data_bus[829]), .B2(n4024), .ZN(n3978) );
  ND4D1BWP30P140LVT U4367 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), 
        .ZN(n3993) );
  INVD1BWP30P140LVT U4368 ( .I(i_data_bus[381]), .ZN(n6117) );
  INVD1BWP30P140LVT U4369 ( .I(i_data_bus[285]), .ZN(n5352) );
  OAI22D1BWP30P140LVT U4370 ( .A1(n6117), .A2(n3983), .B1(n5352), .B2(n3982), 
        .ZN(n3992) );
  MOAI22D1BWP30P140LVT U4371 ( .A1(n3985), .A2(n3984), .B1(i_data_bus[317]), 
        .B2(n3347), .ZN(n3991) );
  AOI22D1BWP30P140LVT U4372 ( .A1(i_data_bus[1021]), .A2(n3383), .B1(
        i_data_bus[541]), .B2(n4052), .ZN(n3989) );
  AOI22D1BWP30P140LVT U4373 ( .A1(i_data_bus[637]), .A2(n4049), .B1(
        i_data_bus[989]), .B2(n4048), .ZN(n3988) );
  AOI22D1BWP30P140LVT U4374 ( .A1(i_data_bus[925]), .A2(n3378), .B1(
        i_data_bus[605]), .B2(n4050), .ZN(n3987) );
  AOI22D1BWP30P140LVT U4375 ( .A1(i_data_bus[957]), .A2(n4051), .B1(
        i_data_bus[573]), .B2(n4047), .ZN(n3986) );
  ND4D1BWP30P140LVT U4376 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), 
        .ZN(n3990) );
  NR4D0BWP30P140LVT U4377 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), 
        .ZN(n3994) );
  ND4D1BWP30P140LVT U4378 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), 
        .ZN(o_data_bus[93]) );
  AOI22D1BWP30P140LVT U4379 ( .A1(i_data_bus[446]), .A2(n4021), .B1(
        i_data_bus[510]), .B2(n4020), .ZN(n4019) );
  AOI22D1BWP30P140LVT U4380 ( .A1(i_data_bus[350]), .A2(n3348), .B1(
        i_data_bus[318]), .B2(n3347), .ZN(n4018) );
  AOI22D1BWP30P140LVT U4381 ( .A1(i_data_bus[766]), .A2(n3353), .B1(
        i_data_bus[830]), .B2(n4024), .ZN(n4001) );
  AOI22D1BWP30P140LVT U4382 ( .A1(i_data_bus[670]), .A2(n4040), .B1(
        i_data_bus[190]), .B2(n4037), .ZN(n4000) );
  AOI22D1BWP30P140LVT U4383 ( .A1(i_data_bus[862]), .A2(n4036), .B1(
        i_data_bus[798]), .B2(n4027), .ZN(n3999) );
  AOI22D1BWP30P140LVT U4384 ( .A1(i_data_bus[62]), .A2(n4025), .B1(
        i_data_bus[894]), .B2(n4039), .ZN(n3998) );
  AOI22D1BWP30P140LVT U4385 ( .A1(i_data_bus[286]), .A2(n4023), .B1(
        i_data_bus[382]), .B2(n4033), .ZN(n4015) );
  AOI22D1BWP30P140LVT U4386 ( .A1(i_data_bus[734]), .A2(n3360), .B1(
        i_data_bus[158]), .B2(n3355), .ZN(n4005) );
  AOI22D1BWP30P140LVT U4387 ( .A1(i_data_bus[126]), .A2(n4026), .B1(
        i_data_bus[254]), .B2(n3352), .ZN(n4004) );
  AOI22D1BWP30P140LVT U4388 ( .A1(i_data_bus[94]), .A2(n4028), .B1(
        i_data_bus[222]), .B2(n3351), .ZN(n4003) );
  AOI22D1BWP30P140LVT U4389 ( .A1(i_data_bus[30]), .A2(n4038), .B1(
        i_data_bus[702]), .B2(n4035), .ZN(n4002) );
  ND4D1BWP30P140LVT U4390 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), 
        .ZN(n4014) );
  MOAI22D1BWP30P140LVT U4391 ( .A1(n6138), .A2(n4007), .B1(i_data_bus[478]), 
        .B2(n4006), .ZN(n4013) );
  AOI22D1BWP30P140LVT U4392 ( .A1(i_data_bus[958]), .A2(n4051), .B1(
        i_data_bus[1022]), .B2(n3383), .ZN(n4011) );
  AOI22D1BWP30P140LVT U4393 ( .A1(i_data_bus[926]), .A2(n3378), .B1(
        i_data_bus[990]), .B2(n4048), .ZN(n4010) );
  AOI22D1BWP30P140LVT U4394 ( .A1(i_data_bus[606]), .A2(n4050), .B1(
        i_data_bus[638]), .B2(n4049), .ZN(n4009) );
  AOI22D1BWP30P140LVT U4395 ( .A1(i_data_bus[542]), .A2(n4052), .B1(
        i_data_bus[574]), .B2(n4047), .ZN(n4008) );
  ND4D1BWP30P140LVT U4396 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), 
        .ZN(n4012) );
  INR4D0BWP30P140LVT U4397 ( .A1(n4015), .B1(n4014), .B2(n4013), .B3(n4012), 
        .ZN(n4016) );
  ND4D1BWP30P140LVT U4398 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), 
        .ZN(o_data_bus[94]) );
  AOI22D1BWP30P140LVT U4399 ( .A1(i_data_bus[447]), .A2(n4021), .B1(
        i_data_bus[511]), .B2(n4020), .ZN(n4064) );
  AOI22D1BWP30P140LVT U4400 ( .A1(i_data_bus[287]), .A2(n4023), .B1(
        i_data_bus[415]), .B2(n4022), .ZN(n4063) );
  AOI22D1BWP30P140LVT U4401 ( .A1(i_data_bus[63]), .A2(n4025), .B1(
        i_data_bus[831]), .B2(n4024), .ZN(n4032) );
  AOI22D1BWP30P140LVT U4402 ( .A1(i_data_bus[735]), .A2(n3360), .B1(
        i_data_bus[767]), .B2(n3353), .ZN(n4031) );
  AOI22D1BWP30P140LVT U4403 ( .A1(i_data_bus[127]), .A2(n4026), .B1(
        i_data_bus[223]), .B2(n3351), .ZN(n4030) );
  AOI22D1BWP30P140LVT U4404 ( .A1(i_data_bus[95]), .A2(n4028), .B1(
        i_data_bus[799]), .B2(n4027), .ZN(n4029) );
  AOI22D1BWP30P140LVT U4405 ( .A1(i_data_bus[319]), .A2(n3347), .B1(
        i_data_bus[383]), .B2(n4033), .ZN(n4060) );
  AOI22D1BWP30P140LVT U4406 ( .A1(i_data_bus[863]), .A2(n4036), .B1(
        i_data_bus[703]), .B2(n4035), .ZN(n4044) );
  AOI22D1BWP30P140LVT U4407 ( .A1(i_data_bus[159]), .A2(n3355), .B1(
        i_data_bus[255]), .B2(n3352), .ZN(n4043) );
  AOI22D1BWP30P140LVT U4408 ( .A1(i_data_bus[31]), .A2(n4038), .B1(
        i_data_bus[191]), .B2(n4037), .ZN(n4042) );
  AOI22D1BWP30P140LVT U4409 ( .A1(i_data_bus[671]), .A2(n4040), .B1(
        i_data_bus[895]), .B2(n4039), .ZN(n4041) );
  ND4D1BWP30P140LVT U4410 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), 
        .ZN(n4059) );
  INVD1BWP30P140LVT U4411 ( .I(i_data_bus[479]), .ZN(n5409) );
  MOAI22D1BWP30P140LVT U4412 ( .A1(n5409), .A2(n4046), .B1(i_data_bus[351]), 
        .B2(n3348), .ZN(n4058) );
  AOI22D1BWP30P140LVT U4413 ( .A1(i_data_bus[991]), .A2(n4048), .B1(
        i_data_bus[575]), .B2(n4047), .ZN(n4056) );
  AOI22D1BWP30P140LVT U4414 ( .A1(i_data_bus[927]), .A2(n3378), .B1(
        i_data_bus[639]), .B2(n4049), .ZN(n4055) );
  AOI22D1BWP30P140LVT U4415 ( .A1(i_data_bus[1023]), .A2(n3383), .B1(
        i_data_bus[607]), .B2(n4050), .ZN(n4054) );
  AOI22D1BWP30P140LVT U4416 ( .A1(i_data_bus[543]), .A2(n4052), .B1(
        i_data_bus[959]), .B2(n4051), .ZN(n4053) );
  ND4D1BWP30P140LVT U4417 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), 
        .ZN(n4057) );
  INR4D0BWP30P140LVT U4418 ( .A1(n4060), .B1(n4059), .B2(n4058), .B3(n4057), 
        .ZN(n4061) );
  ND4D1BWP30P140LVT U4419 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), 
        .ZN(o_data_bus[95]) );
  AOI22D1BWP30P140LVT U4420 ( .A1(i_data_bus[992]), .A2(n4066), .B1(
        i_data_bus[960]), .B2(n4068), .ZN(n4080) );
  AOI22D1BWP30P140LVT U4421 ( .A1(i_data_bus[928]), .A2(n4070), .B1(
        i_data_bus[896]), .B2(n4073), .ZN(n4079) );
  INR3D2BWP30P140LVT U4422 ( .A1(i_cmd[94]), .B1(n4074), .B2(n4094), .ZN(n4739) );
  AOI22D1BWP30P140LVT U4423 ( .A1(i_data_bus[352]), .A2(n4739), .B1(
        i_data_bus[672]), .B2(n4075), .ZN(n4078) );
  INR3D2BWP30P140LVT U4424 ( .A1(i_cmd[158]), .B1(n5478), .B2(n4102), .ZN(
        n4733) );
  AOI22D1BWP30P140LVT U4425 ( .A1(i_data_bus[608]), .A2(n4733), .B1(
        i_data_bus[800]), .B2(n4076), .ZN(n4077) );
  ND4D1BWP30P140LVT U4426 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), 
        .ZN(n4120) );
  INR3D2BWP30P140LVT U4427 ( .A1(i_cmd[150]), .B1(n5481), .B2(n4102), .ZN(
        n4742) );
  INVD1BWP30P140LVT U4428 ( .I(i_cmd[70]), .ZN(n4081) );
  NR3D0P7BWP30P140LVT U4429 ( .A1(n5497), .A2(n4081), .A3(n4094), .ZN(n4082)
         );
  AOI22D1BWP30P140LVT U4430 ( .A1(i_data_bus[576]), .A2(n4742), .B1(
        i_data_bus[256]), .B2(n4731), .ZN(n4092) );
  INR3D2BWP30P140LVT U4431 ( .A1(i_cmd[118]), .B1(n4083), .B2(n4109), .ZN(
        n4751) );
  INR3D2BWP30P140LVT U4432 ( .A1(i_cmd[86]), .B1(n4084), .B2(n4094), .ZN(n4729) );
  AOI22D1BWP30P140LVT U4433 ( .A1(i_data_bus[448]), .A2(n4751), .B1(
        i_data_bus[320]), .B2(n4729), .ZN(n4091) );
  INR3D2BWP30P140LVT U4434 ( .A1(i_cmd[110]), .B1(n4085), .B2(n4109), .ZN(
        n4732) );
  INVD1BWP30P140LVT U4435 ( .I(i_cmd[166]), .ZN(n4086) );
  NR3D0P7BWP30P140LVT U4436 ( .A1(n5455), .A2(n4086), .A3(n4093), .ZN(n4087)
         );
  BUFFD2BWP30P140LVT U4437 ( .I(n4087), .Z(n4730) );
  AOI22D1BWP30P140LVT U4438 ( .A1(i_data_bus[416]), .A2(n4732), .B1(
        i_data_bus[640]), .B2(n4730), .ZN(n4090) );
  INR3D2BWP30P140LVT U4439 ( .A1(i_cmd[62]), .B1(n5471), .B2(n4112), .ZN(n4749) );
  AOI22D1BWP30P140LVT U4440 ( .A1(i_data_bus[736]), .A2(n4088), .B1(
        i_data_bus[224]), .B2(n4749), .ZN(n4089) );
  ND4D1BWP30P140LVT U4441 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), 
        .ZN(n4119) );
  INR3D2BWP30P140LVT U4442 ( .A1(i_cmd[14]), .B1(n5442), .B2(n4107), .ZN(n4740) );
  INR3D2BWP30P140LVT U4443 ( .A1(i_cmd[182]), .B1(n5448), .B2(n4093), .ZN(
        n4753) );
  AOI22D1BWP30P140LVT U4444 ( .A1(i_data_bus[32]), .A2(n4740), .B1(
        i_data_bus[704]), .B2(n4753), .ZN(n4101) );
  INR3D2BWP30P140LVT U4445 ( .A1(i_cmd[142]), .B1(n5479), .B2(n4102), .ZN(
        n4723) );
  INR3D2BWP30P140LVT U4446 ( .A1(i_cmd[78]), .B1(n4095), .B2(n4094), .ZN(n4741) );
  AOI22D1BWP30P140LVT U4447 ( .A1(i_data_bus[544]), .A2(n4723), .B1(
        i_data_bus[288]), .B2(n4741), .ZN(n4100) );
  NR3D1P5BWP30P140LVT U4448 ( .A1(n5476), .A2(n132), .A3(n4109), .ZN(n4752) );
  AOI22D1BWP30P140LVT U4449 ( .A1(i_data_bus[384]), .A2(n4752), .B1(
        i_data_bus[832]), .B2(n4096), .ZN(n4099) );
  INR3D2BWP30P140LVT U4450 ( .A1(i_cmd[54]), .B1(n5494), .B2(n4112), .ZN(n4744) );
  AOI22D1BWP30P140LVT U4451 ( .A1(i_data_bus[0]), .A2(n4097), .B1(
        i_data_bus[192]), .B2(n4744), .ZN(n4098) );
  ND4D1BWP30P140LVT U4452 ( .A1(n4101), .A2(n4100), .A3(n4099), .A4(n4098), 
        .ZN(n4118) );
  INVD1BWP30P140LVT U4453 ( .I(i_cmd[134]), .ZN(n4103) );
  INVD1BWP30P140LVT U4454 ( .I(i_cmd[198]), .ZN(n4104) );
  NR3D0P7BWP30P140LVT U4455 ( .A1(n5444), .A2(n4104), .A3(n4106), .ZN(n4105)
         );
  AOI22D1BWP30P140LVT U4456 ( .A1(i_data_bus[512]), .A2(n4722), .B1(
        i_data_bus[768]), .B2(n4721), .ZN(n4116) );
  INR3D2BWP30P140LVT U4457 ( .A1(i_cmd[30]), .B1(n5446), .B2(n4107), .ZN(n4750) );
  INR3D2BWP30P140LVT U4458 ( .A1(i_cmd[222]), .B1(n5457), .B2(n4106), .ZN(
        n4743) );
  AOI22D1BWP30P140LVT U4459 ( .A1(i_data_bus[96]), .A2(n4750), .B1(
        i_data_bus[864]), .B2(n4743), .ZN(n4115) );
  INR3D2BWP30P140LVT U4460 ( .A1(i_cmd[22]), .B1(n5451), .B2(n4107), .ZN(n4724) );
  AOI22D1BWP30P140LVT U4461 ( .A1(i_data_bus[64]), .A2(n4724), .B1(
        i_data_bus[128]), .B2(n4108), .ZN(n4114) );
  INR3D2BWP30P140LVT U4462 ( .A1(i_cmd[46]), .B1(n5487), .B2(n4112), .ZN(n4738) );
  AOI22D1BWP30P140LVT U4463 ( .A1(i_data_bus[480]), .A2(n4111), .B1(
        i_data_bus[160]), .B2(n4738), .ZN(n4113) );
  ND4D1BWP30P140LVT U4464 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), 
        .ZN(n4117) );
  OR4D1BWP30P140LVT U4465 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), 
        .Z(o_data_bus[192]) );
  AOI22D1BWP30P140LVT U4466 ( .A1(i_data_bus[897]), .A2(n4073), .B1(
        i_data_bus[993]), .B2(n4066), .ZN(n4124) );
  AOI22D1BWP30P140LVT U4467 ( .A1(i_data_bus[961]), .A2(n4068), .B1(
        i_data_bus[929]), .B2(n4070), .ZN(n4123) );
  AOI22D1BWP30P140LVT U4468 ( .A1(i_data_bus[193]), .A2(n4744), .B1(
        i_data_bus[833]), .B2(n4096), .ZN(n4122) );
  AOI22D1BWP30P140LVT U4469 ( .A1(i_data_bus[609]), .A2(n4733), .B1(
        i_data_bus[353]), .B2(n4739), .ZN(n4121) );
  ND4D1BWP30P140LVT U4470 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), 
        .ZN(n4140) );
  AOI22D1BWP30P140LVT U4471 ( .A1(i_data_bus[65]), .A2(n4724), .B1(
        i_data_bus[417]), .B2(n4732), .ZN(n4128) );
  AOI22D1BWP30P140LVT U4472 ( .A1(i_data_bus[289]), .A2(n4741), .B1(
        i_data_bus[321]), .B2(n4729), .ZN(n4127) );
  AOI22D1BWP30P140LVT U4473 ( .A1(i_data_bus[97]), .A2(n4750), .B1(
        i_data_bus[769]), .B2(n4721), .ZN(n4126) );
  AOI22D1BWP30P140LVT U4474 ( .A1(i_data_bus[513]), .A2(n4722), .B1(
        i_data_bus[673]), .B2(n4075), .ZN(n4125) );
  ND4D1BWP30P140LVT U4475 ( .A1(n4128), .A2(n4127), .A3(n4126), .A4(n4125), 
        .ZN(n4139) );
  AOI22D1BWP30P140LVT U4476 ( .A1(i_data_bus[1]), .A2(n4097), .B1(
        i_data_bus[257]), .B2(n4731), .ZN(n4132) );
  AOI22D1BWP30P140LVT U4477 ( .A1(i_data_bus[33]), .A2(n4740), .B1(
        i_data_bus[449]), .B2(n4751), .ZN(n4131) );
  AOI22D1BWP30P140LVT U4478 ( .A1(i_data_bus[705]), .A2(n4753), .B1(
        i_data_bus[865]), .B2(n4743), .ZN(n4130) );
  AOI22D1BWP30P140LVT U4479 ( .A1(i_data_bus[577]), .A2(n4742), .B1(
        i_data_bus[161]), .B2(n4738), .ZN(n4129) );
  ND4D1BWP30P140LVT U4480 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), 
        .ZN(n4138) );
  AOI22D1BWP30P140LVT U4481 ( .A1(i_data_bus[641]), .A2(n4730), .B1(
        i_data_bus[481]), .B2(n4111), .ZN(n4136) );
  AOI22D1BWP30P140LVT U4482 ( .A1(i_data_bus[385]), .A2(n4752), .B1(
        i_data_bus[737]), .B2(n4088), .ZN(n4135) );
  AOI22D1BWP30P140LVT U4483 ( .A1(i_data_bus[801]), .A2(n4076), .B1(
        i_data_bus[225]), .B2(n4749), .ZN(n4134) );
  AOI22D1BWP30P140LVT U4484 ( .A1(i_data_bus[545]), .A2(n4723), .B1(
        i_data_bus[129]), .B2(n4108), .ZN(n4133) );
  ND4D1BWP30P140LVT U4485 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), 
        .ZN(n4137) );
  OR4D1BWP30P140LVT U4486 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), 
        .Z(o_data_bus[193]) );
  AOI22D1BWP30P140LVT U4487 ( .A1(i_data_bus[962]), .A2(n4068), .B1(
        i_data_bus[930]), .B2(n4070), .ZN(n4144) );
  AOI22D1BWP30P140LVT U4488 ( .A1(i_data_bus[898]), .A2(n4073), .B1(
        i_data_bus[994]), .B2(n4066), .ZN(n4143) );
  AOI22D1BWP30P140LVT U4489 ( .A1(i_data_bus[674]), .A2(n4075), .B1(
        i_data_bus[770]), .B2(n4721), .ZN(n4142) );
  AOI22D1BWP30P140LVT U4490 ( .A1(i_data_bus[98]), .A2(n4750), .B1(
        i_data_bus[226]), .B2(n4749), .ZN(n4141) );
  ND4D1BWP30P140LVT U4491 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), 
        .ZN(n4160) );
  AOI22D1BWP30P140LVT U4492 ( .A1(i_data_bus[546]), .A2(n4723), .B1(
        i_data_bus[706]), .B2(n4753), .ZN(n4148) );
  AOI22D1BWP30P140LVT U4493 ( .A1(i_data_bus[610]), .A2(n4733), .B1(
        i_data_bus[834]), .B2(n4096), .ZN(n4147) );
  AOI22D1BWP30P140LVT U4494 ( .A1(i_data_bus[66]), .A2(n4724), .B1(
        i_data_bus[514]), .B2(n4722), .ZN(n4146) );
  AOI22D1BWP30P140LVT U4495 ( .A1(i_data_bus[34]), .A2(n4740), .B1(
        i_data_bus[354]), .B2(n4739), .ZN(n4145) );
  ND4D1BWP30P140LVT U4496 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), 
        .ZN(n4159) );
  AOI22D1BWP30P140LVT U4497 ( .A1(i_data_bus[290]), .A2(n4741), .B1(
        i_data_bus[802]), .B2(n4076), .ZN(n4152) );
  AOI22D1BWP30P140LVT U4498 ( .A1(i_data_bus[162]), .A2(n4738), .B1(
        i_data_bus[258]), .B2(n4731), .ZN(n4151) );
  AOI22D1BWP30P140LVT U4499 ( .A1(i_data_bus[194]), .A2(n4744), .B1(
        i_data_bus[322]), .B2(n4729), .ZN(n4150) );
  AOI22D1BWP30P140LVT U4500 ( .A1(i_data_bus[2]), .A2(n4097), .B1(
        i_data_bus[418]), .B2(n4732), .ZN(n4149) );
  ND4D1BWP30P140LVT U4501 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), 
        .ZN(n4158) );
  AOI22D1BWP30P140LVT U4502 ( .A1(i_data_bus[578]), .A2(n4742), .B1(
        i_data_bus[866]), .B2(n4743), .ZN(n4156) );
  AOI22D1BWP30P140LVT U4503 ( .A1(i_data_bus[386]), .A2(n4752), .B1(
        i_data_bus[738]), .B2(n4088), .ZN(n4155) );
  AOI22D1BWP30P140LVT U4504 ( .A1(i_data_bus[450]), .A2(n4751), .B1(
        i_data_bus[130]), .B2(n4108), .ZN(n4154) );
  AOI22D1BWP30P140LVT U4505 ( .A1(i_data_bus[482]), .A2(n4111), .B1(
        i_data_bus[642]), .B2(n4730), .ZN(n4153) );
  ND4D1BWP30P140LVT U4506 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), 
        .ZN(n4157) );
  OR4D1BWP30P140LVT U4507 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), 
        .Z(o_data_bus[194]) );
  AOI22D1BWP30P140LVT U4508 ( .A1(i_data_bus[963]), .A2(n4068), .B1(
        i_data_bus[995]), .B2(n4066), .ZN(n4164) );
  AOI22D1BWP30P140LVT U4509 ( .A1(i_data_bus[899]), .A2(n4073), .B1(
        i_data_bus[931]), .B2(n4070), .ZN(n4163) );
  AOI22D1BWP30P140LVT U4510 ( .A1(i_data_bus[3]), .A2(n4097), .B1(
        i_data_bus[323]), .B2(n4729), .ZN(n4162) );
  AOI22D1BWP30P140LVT U4511 ( .A1(i_data_bus[99]), .A2(n4750), .B1(
        i_data_bus[387]), .B2(n4752), .ZN(n4161) );
  ND4D1BWP30P140LVT U4512 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), 
        .ZN(n4180) );
  AOI22D1BWP30P140LVT U4513 ( .A1(i_data_bus[67]), .A2(n4724), .B1(
        i_data_bus[483]), .B2(n4111), .ZN(n4168) );
  AOI22D1BWP30P140LVT U4514 ( .A1(i_data_bus[163]), .A2(n4738), .B1(
        i_data_bus[707]), .B2(n4753), .ZN(n4167) );
  AOI22D1BWP30P140LVT U4515 ( .A1(i_data_bus[547]), .A2(n4723), .B1(
        i_data_bus[643]), .B2(n4730), .ZN(n4166) );
  AOI22D1BWP30P140LVT U4516 ( .A1(i_data_bus[771]), .A2(n4721), .B1(
        i_data_bus[867]), .B2(n4743), .ZN(n4165) );
  ND4D1BWP30P140LVT U4517 ( .A1(n4168), .A2(n4167), .A3(n4166), .A4(n4165), 
        .ZN(n4179) );
  AOI22D1BWP30P140LVT U4518 ( .A1(i_data_bus[675]), .A2(n4075), .B1(
        i_data_bus[451]), .B2(n4751), .ZN(n4172) );
  AOI22D1BWP30P140LVT U4519 ( .A1(i_data_bus[739]), .A2(n4088), .B1(
        i_data_bus[227]), .B2(n4749), .ZN(n4171) );
  AOI22D1BWP30P140LVT U4520 ( .A1(i_data_bus[355]), .A2(n4739), .B1(
        i_data_bus[803]), .B2(n4076), .ZN(n4170) );
  AOI22D1BWP30P140LVT U4521 ( .A1(i_data_bus[611]), .A2(n4733), .B1(
        i_data_bus[259]), .B2(n4731), .ZN(n4169) );
  ND4D1BWP30P140LVT U4522 ( .A1(n4172), .A2(n4171), .A3(n4170), .A4(n4169), 
        .ZN(n4178) );
  AOI22D1BWP30P140LVT U4523 ( .A1(i_data_bus[579]), .A2(n4742), .B1(
        i_data_bus[835]), .B2(n4096), .ZN(n4176) );
  AOI22D1BWP30P140LVT U4524 ( .A1(i_data_bus[515]), .A2(n4722), .B1(
        i_data_bus[35]), .B2(n4740), .ZN(n4175) );
  AOI22D1BWP30P140LVT U4525 ( .A1(i_data_bus[419]), .A2(n4732), .B1(
        i_data_bus[291]), .B2(n4741), .ZN(n4174) );
  AOI22D1BWP30P140LVT U4526 ( .A1(i_data_bus[131]), .A2(n4108), .B1(
        i_data_bus[195]), .B2(n4744), .ZN(n4173) );
  ND4D1BWP30P140LVT U4527 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), 
        .ZN(n4177) );
  OR4D1BWP30P140LVT U4528 ( .A1(n4180), .A2(n4179), .A3(n4178), .A4(n4177), 
        .Z(o_data_bus[195]) );
  AOI22D1BWP30P140LVT U4529 ( .A1(i_data_bus[964]), .A2(n4068), .B1(
        i_data_bus[996]), .B2(n4066), .ZN(n4184) );
  AOI22D1BWP30P140LVT U4530 ( .A1(i_data_bus[932]), .A2(n4070), .B1(
        i_data_bus[900]), .B2(n4073), .ZN(n4183) );
  AOI22D1BWP30P140LVT U4531 ( .A1(i_data_bus[740]), .A2(n4088), .B1(
        i_data_bus[676]), .B2(n4075), .ZN(n4182) );
  AOI22D1BWP30P140LVT U4532 ( .A1(i_data_bus[100]), .A2(n4750), .B1(
        i_data_bus[196]), .B2(n4744), .ZN(n4181) );
  ND4D1BWP30P140LVT U4533 ( .A1(n4184), .A2(n4183), .A3(n4182), .A4(n4181), 
        .ZN(n4200) );
  AOI22D1BWP30P140LVT U4534 ( .A1(i_data_bus[548]), .A2(n4723), .B1(
        i_data_bus[420]), .B2(n4732), .ZN(n4188) );
  AOI22D1BWP30P140LVT U4535 ( .A1(i_data_bus[708]), .A2(n4753), .B1(
        i_data_bus[228]), .B2(n4749), .ZN(n4187) );
  AOI22D1BWP30P140LVT U4536 ( .A1(i_data_bus[4]), .A2(n4097), .B1(
        i_data_bus[260]), .B2(n4731), .ZN(n4186) );
  AOI22D1BWP30P140LVT U4537 ( .A1(i_data_bus[292]), .A2(n4741), .B1(
        i_data_bus[644]), .B2(n4730), .ZN(n4185) );
  ND4D1BWP30P140LVT U4538 ( .A1(n4188), .A2(n4187), .A3(n4186), .A4(n4185), 
        .ZN(n4199) );
  AOI22D1BWP30P140LVT U4539 ( .A1(i_data_bus[324]), .A2(n4729), .B1(
        i_data_bus[356]), .B2(n4739), .ZN(n4192) );
  AOI22D1BWP30P140LVT U4540 ( .A1(i_data_bus[612]), .A2(n4733), .B1(
        i_data_bus[772]), .B2(n4721), .ZN(n4191) );
  AOI22D1BWP30P140LVT U4541 ( .A1(i_data_bus[132]), .A2(n4108), .B1(
        i_data_bus[388]), .B2(n4752), .ZN(n4190) );
  AOI22D1BWP30P140LVT U4542 ( .A1(i_data_bus[580]), .A2(n4742), .B1(
        i_data_bus[804]), .B2(n4076), .ZN(n4189) );
  ND4D1BWP30P140LVT U4543 ( .A1(n4192), .A2(n4191), .A3(n4190), .A4(n4189), 
        .ZN(n4198) );
  AOI22D1BWP30P140LVT U4544 ( .A1(i_data_bus[452]), .A2(n4751), .B1(
        i_data_bus[868]), .B2(n4743), .ZN(n4196) );
  AOI22D1BWP30P140LVT U4545 ( .A1(i_data_bus[164]), .A2(n4738), .B1(
        i_data_bus[836]), .B2(n4096), .ZN(n4195) );
  AOI22D1BWP30P140LVT U4546 ( .A1(i_data_bus[68]), .A2(n4724), .B1(
        i_data_bus[36]), .B2(n4740), .ZN(n4194) );
  AOI22D1BWP30P140LVT U4547 ( .A1(i_data_bus[516]), .A2(n4722), .B1(
        i_data_bus[484]), .B2(n4111), .ZN(n4193) );
  ND4D1BWP30P140LVT U4548 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), 
        .ZN(n4197) );
  OR4D1BWP30P140LVT U4549 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), 
        .Z(o_data_bus[196]) );
  AOI22D1BWP30P140LVT U4550 ( .A1(i_data_bus[933]), .A2(n4070), .B1(
        i_data_bus[997]), .B2(n4066), .ZN(n4204) );
  AOI22D1BWP30P140LVT U4551 ( .A1(i_data_bus[901]), .A2(n4073), .B1(
        i_data_bus[965]), .B2(n4068), .ZN(n4203) );
  AOI22D1BWP30P140LVT U4552 ( .A1(i_data_bus[517]), .A2(n4722), .B1(
        i_data_bus[261]), .B2(n4731), .ZN(n4202) );
  AOI22D1BWP30P140LVT U4553 ( .A1(i_data_bus[165]), .A2(n4738), .B1(
        i_data_bus[293]), .B2(n4741), .ZN(n4201) );
  ND4D1BWP30P140LVT U4554 ( .A1(n4204), .A2(n4203), .A3(n4202), .A4(n4201), 
        .ZN(n4220) );
  AOI22D1BWP30P140LVT U4555 ( .A1(i_data_bus[613]), .A2(n4733), .B1(
        i_data_bus[837]), .B2(n4096), .ZN(n4208) );
  AOI22D1BWP30P140LVT U4556 ( .A1(i_data_bus[805]), .A2(n4076), .B1(
        i_data_bus[741]), .B2(n4088), .ZN(n4207) );
  AOI22D1BWP30P140LVT U4557 ( .A1(i_data_bus[69]), .A2(n4724), .B1(
        i_data_bus[485]), .B2(n4111), .ZN(n4206) );
  AOI22D1BWP30P140LVT U4558 ( .A1(i_data_bus[709]), .A2(n4753), .B1(
        i_data_bus[133]), .B2(n4108), .ZN(n4205) );
  ND4D1BWP30P140LVT U4559 ( .A1(n4208), .A2(n4207), .A3(n4206), .A4(n4205), 
        .ZN(n4219) );
  AOI22D1BWP30P140LVT U4560 ( .A1(i_data_bus[869]), .A2(n4743), .B1(
        i_data_bus[325]), .B2(n4729), .ZN(n4212) );
  AOI22D1BWP30P140LVT U4561 ( .A1(i_data_bus[197]), .A2(n4744), .B1(
        i_data_bus[645]), .B2(n4730), .ZN(n4211) );
  AOI22D1BWP30P140LVT U4562 ( .A1(i_data_bus[581]), .A2(n4742), .B1(
        i_data_bus[773]), .B2(n4721), .ZN(n4210) );
  AOI22D1BWP30P140LVT U4563 ( .A1(i_data_bus[453]), .A2(n4751), .B1(
        i_data_bus[389]), .B2(n4752), .ZN(n4209) );
  ND4D1BWP30P140LVT U4564 ( .A1(n4212), .A2(n4211), .A3(n4210), .A4(n4209), 
        .ZN(n4218) );
  AOI22D1BWP30P140LVT U4565 ( .A1(i_data_bus[37]), .A2(n4740), .B1(
        i_data_bus[101]), .B2(n4750), .ZN(n4216) );
  AOI22D1BWP30P140LVT U4566 ( .A1(i_data_bus[357]), .A2(n4739), .B1(
        i_data_bus[229]), .B2(n4749), .ZN(n4215) );
  AOI22D1BWP30P140LVT U4567 ( .A1(i_data_bus[5]), .A2(n4097), .B1(
        i_data_bus[421]), .B2(n4732), .ZN(n4214) );
  AOI22D1BWP30P140LVT U4568 ( .A1(i_data_bus[549]), .A2(n4723), .B1(
        i_data_bus[677]), .B2(n4075), .ZN(n4213) );
  ND4D1BWP30P140LVT U4569 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), 
        .ZN(n4217) );
  OR4D1BWP30P140LVT U4570 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), 
        .Z(o_data_bus[197]) );
  AOI22D1BWP30P140LVT U4571 ( .A1(i_data_bus[934]), .A2(n4070), .B1(
        i_data_bus[902]), .B2(n4073), .ZN(n4224) );
  AOI22D1BWP30P140LVT U4572 ( .A1(i_data_bus[966]), .A2(n4068), .B1(
        i_data_bus[998]), .B2(n4066), .ZN(n4223) );
  AOI22D1BWP30P140LVT U4573 ( .A1(i_data_bus[6]), .A2(n4097), .B1(
        i_data_bus[806]), .B2(n4076), .ZN(n4222) );
  AOI22D1BWP30P140LVT U4574 ( .A1(i_data_bus[742]), .A2(n4088), .B1(
        i_data_bus[326]), .B2(n4729), .ZN(n4221) );
  ND4D1BWP30P140LVT U4575 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), 
        .ZN(n4240) );
  AOI22D1BWP30P140LVT U4576 ( .A1(i_data_bus[70]), .A2(n4724), .B1(
        i_data_bus[678]), .B2(n4075), .ZN(n4228) );
  AOI22D1BWP30P140LVT U4577 ( .A1(i_data_bus[550]), .A2(n4723), .B1(
        i_data_bus[710]), .B2(n4753), .ZN(n4227) );
  AOI22D1BWP30P140LVT U4578 ( .A1(i_data_bus[38]), .A2(n4740), .B1(
        i_data_bus[134]), .B2(n4108), .ZN(n4226) );
  AOI22D1BWP30P140LVT U4579 ( .A1(i_data_bus[486]), .A2(n4111), .B1(
        i_data_bus[230]), .B2(n4749), .ZN(n4225) );
  ND4D1BWP30P140LVT U4580 ( .A1(n4228), .A2(n4227), .A3(n4226), .A4(n4225), 
        .ZN(n4239) );
  AOI22D1BWP30P140LVT U4581 ( .A1(i_data_bus[838]), .A2(n4096), .B1(
        i_data_bus[166]), .B2(n4738), .ZN(n4232) );
  AOI22D1BWP30P140LVT U4582 ( .A1(i_data_bus[582]), .A2(n4742), .B1(
        i_data_bus[454]), .B2(n4751), .ZN(n4231) );
  AOI22D1BWP30P140LVT U4583 ( .A1(i_data_bus[870]), .A2(n4743), .B1(
        i_data_bus[294]), .B2(n4741), .ZN(n4230) );
  AOI22D1BWP30P140LVT U4584 ( .A1(i_data_bus[102]), .A2(n4750), .B1(
        i_data_bus[358]), .B2(n4739), .ZN(n4229) );
  ND4D1BWP30P140LVT U4585 ( .A1(n4232), .A2(n4231), .A3(n4230), .A4(n4229), 
        .ZN(n4238) );
  AOI22D1BWP30P140LVT U4586 ( .A1(i_data_bus[646]), .A2(n4730), .B1(
        i_data_bus[774]), .B2(n4721), .ZN(n4236) );
  AOI22D1BWP30P140LVT U4587 ( .A1(i_data_bus[390]), .A2(n4752), .B1(
        i_data_bus[198]), .B2(n4744), .ZN(n4235) );
  AOI22D1BWP30P140LVT U4588 ( .A1(i_data_bus[614]), .A2(n4733), .B1(
        i_data_bus[262]), .B2(n4731), .ZN(n4234) );
  AOI22D1BWP30P140LVT U4589 ( .A1(i_data_bus[518]), .A2(n4722), .B1(
        i_data_bus[422]), .B2(n4732), .ZN(n4233) );
  ND4D1BWP30P140LVT U4590 ( .A1(n4236), .A2(n4235), .A3(n4234), .A4(n4233), 
        .ZN(n4237) );
  OR4D1BWP30P140LVT U4591 ( .A1(n4240), .A2(n4239), .A3(n4238), .A4(n4237), 
        .Z(o_data_bus[198]) );
  AOI22D1BWP30P140LVT U4592 ( .A1(i_data_bus[903]), .A2(n4073), .B1(
        i_data_bus[935]), .B2(n4070), .ZN(n4244) );
  AOI22D1BWP30P140LVT U4593 ( .A1(i_data_bus[967]), .A2(n4068), .B1(
        i_data_bus[999]), .B2(n4066), .ZN(n4243) );
  AOI22D1BWP30P140LVT U4594 ( .A1(i_data_bus[615]), .A2(n4733), .B1(
        i_data_bus[487]), .B2(n4111), .ZN(n4242) );
  AOI22D1BWP30P140LVT U4595 ( .A1(i_data_bus[167]), .A2(n4738), .B1(
        i_data_bus[423]), .B2(n4732), .ZN(n4241) );
  ND4D1BWP30P140LVT U4596 ( .A1(n4244), .A2(n4243), .A3(n4242), .A4(n4241), 
        .ZN(n4260) );
  AOI22D1BWP30P140LVT U4597 ( .A1(i_data_bus[7]), .A2(n4097), .B1(
        i_data_bus[327]), .B2(n4729), .ZN(n4248) );
  AOI22D1BWP30P140LVT U4598 ( .A1(i_data_bus[519]), .A2(n4722), .B1(
        i_data_bus[455]), .B2(n4751), .ZN(n4247) );
  AOI22D1BWP30P140LVT U4599 ( .A1(i_data_bus[103]), .A2(n4750), .B1(
        i_data_bus[839]), .B2(n4096), .ZN(n4246) );
  AOI22D1BWP30P140LVT U4600 ( .A1(i_data_bus[71]), .A2(n4724), .B1(
        i_data_bus[775]), .B2(n4721), .ZN(n4245) );
  ND4D1BWP30P140LVT U4601 ( .A1(n4248), .A2(n4247), .A3(n4246), .A4(n4245), 
        .ZN(n4259) );
  AOI22D1BWP30P140LVT U4602 ( .A1(i_data_bus[39]), .A2(n4740), .B1(
        i_data_bus[295]), .B2(n4741), .ZN(n4252) );
  AOI22D1BWP30P140LVT U4603 ( .A1(i_data_bus[391]), .A2(n4752), .B1(
        i_data_bus[199]), .B2(n4744), .ZN(n4251) );
  AOI22D1BWP30P140LVT U4604 ( .A1(i_data_bus[583]), .A2(n4742), .B1(
        i_data_bus[359]), .B2(n4739), .ZN(n4250) );
  AOI22D1BWP30P140LVT U4605 ( .A1(i_data_bus[679]), .A2(n4075), .B1(
        i_data_bus[807]), .B2(n4076), .ZN(n4249) );
  ND4D1BWP30P140LVT U4606 ( .A1(n4252), .A2(n4251), .A3(n4250), .A4(n4249), 
        .ZN(n4258) );
  AOI22D1BWP30P140LVT U4607 ( .A1(i_data_bus[263]), .A2(n4731), .B1(
        i_data_bus[711]), .B2(n4753), .ZN(n4256) );
  AOI22D1BWP30P140LVT U4608 ( .A1(i_data_bus[871]), .A2(n4743), .B1(
        i_data_bus[231]), .B2(n4749), .ZN(n4255) );
  AOI22D1BWP30P140LVT U4609 ( .A1(i_data_bus[743]), .A2(n4088), .B1(
        i_data_bus[135]), .B2(n4108), .ZN(n4254) );
  AOI22D1BWP30P140LVT U4610 ( .A1(i_data_bus[551]), .A2(n4723), .B1(
        i_data_bus[647]), .B2(n4730), .ZN(n4253) );
  ND4D1BWP30P140LVT U4611 ( .A1(n4256), .A2(n4255), .A3(n4254), .A4(n4253), 
        .ZN(n4257) );
  OR4D1BWP30P140LVT U4612 ( .A1(n4260), .A2(n4259), .A3(n4258), .A4(n4257), 
        .Z(o_data_bus[199]) );
  AOI22D1BWP30P140LVT U4613 ( .A1(i_data_bus[936]), .A2(n4070), .B1(
        i_data_bus[904]), .B2(n4073), .ZN(n4264) );
  AOI22D1BWP30P140LVT U4614 ( .A1(i_data_bus[968]), .A2(n4068), .B1(
        i_data_bus[1000]), .B2(n4066), .ZN(n4263) );
  AOI22D1BWP30P140LVT U4615 ( .A1(i_data_bus[264]), .A2(n4731), .B1(
        i_data_bus[392]), .B2(n4752), .ZN(n4262) );
  AOI22D1BWP30P140LVT U4616 ( .A1(i_data_bus[488]), .A2(n4111), .B1(
        i_data_bus[232]), .B2(n4749), .ZN(n4261) );
  ND4D1BWP30P140LVT U4617 ( .A1(n4264), .A2(n4263), .A3(n4262), .A4(n4261), 
        .ZN(n4280) );
  AOI22D1BWP30P140LVT U4618 ( .A1(i_data_bus[72]), .A2(n4724), .B1(
        i_data_bus[168]), .B2(n4738), .ZN(n4268) );
  AOI22D1BWP30P140LVT U4619 ( .A1(i_data_bus[8]), .A2(n4097), .B1(
        i_data_bus[872]), .B2(n4743), .ZN(n4267) );
  AOI22D1BWP30P140LVT U4620 ( .A1(i_data_bus[520]), .A2(n4722), .B1(
        i_data_bus[200]), .B2(n4744), .ZN(n4266) );
  AOI22D1BWP30P140LVT U4621 ( .A1(i_data_bus[456]), .A2(n4751), .B1(
        i_data_bus[296]), .B2(n4741), .ZN(n4265) );
  ND4D1BWP30P140LVT U4622 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), 
        .ZN(n4279) );
  AOI22D1BWP30P140LVT U4623 ( .A1(i_data_bus[840]), .A2(n4096), .B1(
        i_data_bus[648]), .B2(n4730), .ZN(n4272) );
  AOI22D1BWP30P140LVT U4624 ( .A1(i_data_bus[328]), .A2(n4729), .B1(
        i_data_bus[360]), .B2(n4739), .ZN(n4271) );
  AOI22D1BWP30P140LVT U4625 ( .A1(i_data_bus[424]), .A2(n4732), .B1(
        i_data_bus[712]), .B2(n4753), .ZN(n4270) );
  AOI22D1BWP30P140LVT U4626 ( .A1(i_data_bus[680]), .A2(n4075), .B1(
        i_data_bus[776]), .B2(n4721), .ZN(n4269) );
  ND4D1BWP30P140LVT U4627 ( .A1(n4272), .A2(n4271), .A3(n4270), .A4(n4269), 
        .ZN(n4278) );
  AOI22D1BWP30P140LVT U4628 ( .A1(i_data_bus[744]), .A2(n4088), .B1(
        i_data_bus[808]), .B2(n4076), .ZN(n4276) );
  AOI22D1BWP30P140LVT U4629 ( .A1(i_data_bus[616]), .A2(n4733), .B1(
        i_data_bus[40]), .B2(n4740), .ZN(n4275) );
  AOI22D1BWP30P140LVT U4630 ( .A1(i_data_bus[104]), .A2(n4750), .B1(
        i_data_bus[552]), .B2(n4723), .ZN(n4274) );
  AOI22D1BWP30P140LVT U4631 ( .A1(i_data_bus[584]), .A2(n4742), .B1(
        i_data_bus[136]), .B2(n4108), .ZN(n4273) );
  ND4D1BWP30P140LVT U4632 ( .A1(n4276), .A2(n4275), .A3(n4274), .A4(n4273), 
        .ZN(n4277) );
  OR4D1BWP30P140LVT U4633 ( .A1(n4280), .A2(n4279), .A3(n4278), .A4(n4277), 
        .Z(o_data_bus[200]) );
  AOI22D1BWP30P140LVT U4634 ( .A1(i_data_bus[969]), .A2(n4068), .B1(
        i_data_bus[1001]), .B2(n4066), .ZN(n4284) );
  AOI22D1BWP30P140LVT U4635 ( .A1(i_data_bus[905]), .A2(n4073), .B1(
        i_data_bus[937]), .B2(n4070), .ZN(n4283) );
  AOI22D1BWP30P140LVT U4636 ( .A1(i_data_bus[9]), .A2(n4097), .B1(
        i_data_bus[105]), .B2(n4750), .ZN(n4282) );
  AOI22D1BWP30P140LVT U4637 ( .A1(i_data_bus[489]), .A2(n4111), .B1(
        i_data_bus[425]), .B2(n4732), .ZN(n4281) );
  ND4D1BWP30P140LVT U4638 ( .A1(n4284), .A2(n4283), .A3(n4282), .A4(n4281), 
        .ZN(n4300) );
  AOI22D1BWP30P140LVT U4639 ( .A1(i_data_bus[265]), .A2(n4731), .B1(
        i_data_bus[777]), .B2(n4721), .ZN(n4288) );
  AOI22D1BWP30P140LVT U4640 ( .A1(i_data_bus[41]), .A2(n4740), .B1(
        i_data_bus[137]), .B2(n4108), .ZN(n4287) );
  AOI22D1BWP30P140LVT U4641 ( .A1(i_data_bus[585]), .A2(n4742), .B1(
        i_data_bus[329]), .B2(n4729), .ZN(n4286) );
  AOI22D1BWP30P140LVT U4642 ( .A1(i_data_bus[713]), .A2(n4753), .B1(
        i_data_bus[457]), .B2(n4751), .ZN(n4285) );
  ND4D1BWP30P140LVT U4643 ( .A1(n4288), .A2(n4287), .A3(n4286), .A4(n4285), 
        .ZN(n4299) );
  AOI22D1BWP30P140LVT U4644 ( .A1(i_data_bus[201]), .A2(n4744), .B1(
        i_data_bus[393]), .B2(n4752), .ZN(n4292) );
  AOI22D1BWP30P140LVT U4645 ( .A1(i_data_bus[745]), .A2(n4088), .B1(
        i_data_bus[809]), .B2(n4076), .ZN(n4291) );
  AOI22D1BWP30P140LVT U4646 ( .A1(i_data_bus[841]), .A2(n4096), .B1(
        i_data_bus[649]), .B2(n4730), .ZN(n4290) );
  AOI22D1BWP30P140LVT U4647 ( .A1(i_data_bus[617]), .A2(n4733), .B1(
        i_data_bus[233]), .B2(n4749), .ZN(n4289) );
  ND4D1BWP30P140LVT U4648 ( .A1(n4292), .A2(n4291), .A3(n4290), .A4(n4289), 
        .ZN(n4298) );
  AOI22D1BWP30P140LVT U4649 ( .A1(i_data_bus[297]), .A2(n4741), .B1(
        i_data_bus[361]), .B2(n4739), .ZN(n4296) );
  AOI22D1BWP30P140LVT U4650 ( .A1(i_data_bus[553]), .A2(n4723), .B1(
        i_data_bus[169]), .B2(n4738), .ZN(n4295) );
  AOI22D1BWP30P140LVT U4651 ( .A1(i_data_bus[73]), .A2(n4724), .B1(
        i_data_bus[873]), .B2(n4743), .ZN(n4294) );
  AOI22D1BWP30P140LVT U4652 ( .A1(i_data_bus[521]), .A2(n4722), .B1(
        i_data_bus[681]), .B2(n4075), .ZN(n4293) );
  ND4D1BWP30P140LVT U4653 ( .A1(n4296), .A2(n4295), .A3(n4294), .A4(n4293), 
        .ZN(n4297) );
  OR4D1BWP30P140LVT U4654 ( .A1(n4300), .A2(n4299), .A3(n4298), .A4(n4297), 
        .Z(o_data_bus[201]) );
  AOI22D1BWP30P140LVT U4655 ( .A1(i_data_bus[970]), .A2(n4068), .B1(
        i_data_bus[906]), .B2(n4073), .ZN(n4304) );
  AOI22D1BWP30P140LVT U4656 ( .A1(i_data_bus[1002]), .A2(n4066), .B1(
        i_data_bus[938]), .B2(n4070), .ZN(n4303) );
  AOI22D1BWP30P140LVT U4657 ( .A1(i_data_bus[522]), .A2(n4722), .B1(
        i_data_bus[202]), .B2(n4744), .ZN(n4302) );
  AOI22D1BWP30P140LVT U4658 ( .A1(i_data_bus[490]), .A2(n4111), .B1(
        i_data_bus[682]), .B2(n4075), .ZN(n4301) );
  ND4D1BWP30P140LVT U4659 ( .A1(n4304), .A2(n4303), .A3(n4302), .A4(n4301), 
        .ZN(n4320) );
  AOI22D1BWP30P140LVT U4660 ( .A1(i_data_bus[42]), .A2(n4740), .B1(
        i_data_bus[650]), .B2(n4730), .ZN(n4308) );
  AOI22D1BWP30P140LVT U4661 ( .A1(i_data_bus[170]), .A2(n4738), .B1(
        i_data_bus[266]), .B2(n4731), .ZN(n4307) );
  AOI22D1BWP30P140LVT U4662 ( .A1(i_data_bus[554]), .A2(n4723), .B1(
        i_data_bus[74]), .B2(n4724), .ZN(n4306) );
  AOI22D1BWP30P140LVT U4663 ( .A1(i_data_bus[842]), .A2(n4096), .B1(
        i_data_bus[298]), .B2(n4741), .ZN(n4305) );
  ND4D1BWP30P140LVT U4664 ( .A1(n4308), .A2(n4307), .A3(n4306), .A4(n4305), 
        .ZN(n4319) );
  AOI22D1BWP30P140LVT U4665 ( .A1(i_data_bus[778]), .A2(n4721), .B1(
        i_data_bus[362]), .B2(n4739), .ZN(n4312) );
  AOI22D1BWP30P140LVT U4666 ( .A1(i_data_bus[458]), .A2(n4751), .B1(
        i_data_bus[138]), .B2(n4108), .ZN(n4311) );
  AOI22D1BWP30P140LVT U4667 ( .A1(i_data_bus[234]), .A2(n4749), .B1(
        i_data_bus[394]), .B2(n4752), .ZN(n4310) );
  AOI22D1BWP30P140LVT U4668 ( .A1(i_data_bus[586]), .A2(n4742), .B1(
        i_data_bus[330]), .B2(n4729), .ZN(n4309) );
  ND4D1BWP30P140LVT U4669 ( .A1(n4312), .A2(n4311), .A3(n4310), .A4(n4309), 
        .ZN(n4318) );
  AOI22D1BWP30P140LVT U4670 ( .A1(i_data_bus[10]), .A2(n4097), .B1(
        i_data_bus[426]), .B2(n4732), .ZN(n4316) );
  AOI22D1BWP30P140LVT U4671 ( .A1(i_data_bus[714]), .A2(n4753), .B1(
        i_data_bus[746]), .B2(n4088), .ZN(n4315) );
  AOI22D1BWP30P140LVT U4672 ( .A1(i_data_bus[618]), .A2(n4733), .B1(
        i_data_bus[874]), .B2(n4743), .ZN(n4314) );
  AOI22D1BWP30P140LVT U4673 ( .A1(i_data_bus[106]), .A2(n4750), .B1(
        i_data_bus[810]), .B2(n4076), .ZN(n4313) );
  ND4D1BWP30P140LVT U4674 ( .A1(n4316), .A2(n4315), .A3(n4314), .A4(n4313), 
        .ZN(n4317) );
  OR4D1BWP30P140LVT U4675 ( .A1(n4320), .A2(n4319), .A3(n4318), .A4(n4317), 
        .Z(o_data_bus[202]) );
  AOI22D1BWP30P140LVT U4676 ( .A1(i_data_bus[907]), .A2(n4073), .B1(
        i_data_bus[1003]), .B2(n4066), .ZN(n4324) );
  AOI22D1BWP30P140LVT U4677 ( .A1(i_data_bus[939]), .A2(n4070), .B1(
        i_data_bus[971]), .B2(n4068), .ZN(n4323) );
  AOI22D1BWP30P140LVT U4678 ( .A1(i_data_bus[811]), .A2(n4076), .B1(
        i_data_bus[331]), .B2(n4729), .ZN(n4322) );
  AOI22D1BWP30P140LVT U4679 ( .A1(i_data_bus[139]), .A2(n4108), .B1(
        i_data_bus[715]), .B2(n4753), .ZN(n4321) );
  ND4D1BWP30P140LVT U4680 ( .A1(n4324), .A2(n4323), .A3(n4322), .A4(n4321), 
        .ZN(n4340) );
  AOI22D1BWP30P140LVT U4681 ( .A1(i_data_bus[875]), .A2(n4743), .B1(
        i_data_bus[747]), .B2(n4088), .ZN(n4328) );
  AOI22D1BWP30P140LVT U4682 ( .A1(i_data_bus[75]), .A2(n4724), .B1(
        i_data_bus[235]), .B2(n4749), .ZN(n4327) );
  AOI22D1BWP30P140LVT U4683 ( .A1(i_data_bus[43]), .A2(n4740), .B1(
        i_data_bus[843]), .B2(n4096), .ZN(n4326) );
  AOI22D1BWP30P140LVT U4684 ( .A1(i_data_bus[587]), .A2(n4742), .B1(
        i_data_bus[427]), .B2(n4732), .ZN(n4325) );
  ND4D1BWP30P140LVT U4685 ( .A1(n4328), .A2(n4327), .A3(n4326), .A4(n4325), 
        .ZN(n4339) );
  AOI22D1BWP30P140LVT U4686 ( .A1(i_data_bus[619]), .A2(n4733), .B1(
        i_data_bus[555]), .B2(n4723), .ZN(n4332) );
  AOI22D1BWP30P140LVT U4687 ( .A1(i_data_bus[11]), .A2(n4097), .B1(
        i_data_bus[203]), .B2(n4744), .ZN(n4331) );
  AOI22D1BWP30P140LVT U4688 ( .A1(i_data_bus[107]), .A2(n4750), .B1(
        i_data_bus[299]), .B2(n4741), .ZN(n4330) );
  AOI22D1BWP30P140LVT U4689 ( .A1(i_data_bus[523]), .A2(n4722), .B1(
        i_data_bus[491]), .B2(n4111), .ZN(n4329) );
  ND4D1BWP30P140LVT U4690 ( .A1(n4332), .A2(n4331), .A3(n4330), .A4(n4329), 
        .ZN(n4338) );
  AOI22D1BWP30P140LVT U4691 ( .A1(i_data_bus[171]), .A2(n4738), .B1(
        i_data_bus[651]), .B2(n4730), .ZN(n4336) );
  AOI22D1BWP30P140LVT U4692 ( .A1(i_data_bus[363]), .A2(n4739), .B1(
        i_data_bus[459]), .B2(n4751), .ZN(n4335) );
  AOI22D1BWP30P140LVT U4693 ( .A1(i_data_bus[779]), .A2(n4721), .B1(
        i_data_bus[267]), .B2(n4731), .ZN(n4334) );
  AOI22D1BWP30P140LVT U4694 ( .A1(i_data_bus[395]), .A2(n4752), .B1(
        i_data_bus[683]), .B2(n4075), .ZN(n4333) );
  ND4D1BWP30P140LVT U4695 ( .A1(n4336), .A2(n4335), .A3(n4334), .A4(n4333), 
        .ZN(n4337) );
  OR4D1BWP30P140LVT U4696 ( .A1(n4340), .A2(n4339), .A3(n4338), .A4(n4337), 
        .Z(o_data_bus[203]) );
  AOI22D1BWP30P140LVT U4697 ( .A1(i_data_bus[908]), .A2(n4073), .B1(
        i_data_bus[1004]), .B2(n4066), .ZN(n4344) );
  AOI22D1BWP30P140LVT U4698 ( .A1(i_data_bus[940]), .A2(n4070), .B1(
        i_data_bus[972]), .B2(n4068), .ZN(n4343) );
  AOI22D1BWP30P140LVT U4699 ( .A1(i_data_bus[524]), .A2(n4722), .B1(
        i_data_bus[652]), .B2(n4730), .ZN(n4342) );
  AOI22D1BWP30P140LVT U4700 ( .A1(i_data_bus[716]), .A2(n4753), .B1(
        i_data_bus[268]), .B2(n4731), .ZN(n4341) );
  ND4D1BWP30P140LVT U4701 ( .A1(n4344), .A2(n4343), .A3(n4342), .A4(n4341), 
        .ZN(n4360) );
  AOI22D1BWP30P140LVT U4702 ( .A1(i_data_bus[140]), .A2(n4108), .B1(
        i_data_bus[236]), .B2(n4749), .ZN(n4348) );
  AOI22D1BWP30P140LVT U4703 ( .A1(i_data_bus[556]), .A2(n4723), .B1(
        i_data_bus[460]), .B2(n4751), .ZN(n4347) );
  AOI22D1BWP30P140LVT U4704 ( .A1(i_data_bus[108]), .A2(n4750), .B1(
        i_data_bus[300]), .B2(n4741), .ZN(n4346) );
  AOI22D1BWP30P140LVT U4705 ( .A1(i_data_bus[428]), .A2(n4732), .B1(
        i_data_bus[844]), .B2(n4096), .ZN(n4345) );
  ND4D1BWP30P140LVT U4706 ( .A1(n4348), .A2(n4347), .A3(n4346), .A4(n4345), 
        .ZN(n4359) );
  AOI22D1BWP30P140LVT U4707 ( .A1(i_data_bus[780]), .A2(n4721), .B1(
        i_data_bus[332]), .B2(n4729), .ZN(n4352) );
  AOI22D1BWP30P140LVT U4708 ( .A1(i_data_bus[588]), .A2(n4742), .B1(
        i_data_bus[684]), .B2(n4075), .ZN(n4351) );
  AOI22D1BWP30P140LVT U4709 ( .A1(i_data_bus[620]), .A2(n4733), .B1(
        i_data_bus[876]), .B2(n4743), .ZN(n4350) );
  AOI22D1BWP30P140LVT U4710 ( .A1(i_data_bus[44]), .A2(n4740), .B1(
        i_data_bus[172]), .B2(n4738), .ZN(n4349) );
  ND4D1BWP30P140LVT U4711 ( .A1(n4352), .A2(n4351), .A3(n4350), .A4(n4349), 
        .ZN(n4358) );
  AOI22D1BWP30P140LVT U4712 ( .A1(i_data_bus[204]), .A2(n4744), .B1(
        i_data_bus[492]), .B2(n4111), .ZN(n4356) );
  AOI22D1BWP30P140LVT U4713 ( .A1(i_data_bus[364]), .A2(n4739), .B1(
        i_data_bus[396]), .B2(n4752), .ZN(n4355) );
  AOI22D1BWP30P140LVT U4714 ( .A1(i_data_bus[76]), .A2(n4724), .B1(
        i_data_bus[812]), .B2(n4076), .ZN(n4354) );
  AOI22D1BWP30P140LVT U4715 ( .A1(i_data_bus[12]), .A2(n4097), .B1(
        i_data_bus[748]), .B2(n4088), .ZN(n4353) );
  ND4D1BWP30P140LVT U4716 ( .A1(n4356), .A2(n4355), .A3(n4354), .A4(n4353), 
        .ZN(n4357) );
  OR4D1BWP30P140LVT U4717 ( .A1(n4360), .A2(n4359), .A3(n4358), .A4(n4357), 
        .Z(o_data_bus[204]) );
  AOI22D1BWP30P140LVT U4718 ( .A1(i_data_bus[973]), .A2(n4068), .B1(
        i_data_bus[941]), .B2(n4070), .ZN(n4364) );
  AOI22D1BWP30P140LVT U4719 ( .A1(i_data_bus[909]), .A2(n4073), .B1(
        i_data_bus[1005]), .B2(n4066), .ZN(n4363) );
  AOI22D1BWP30P140LVT U4720 ( .A1(i_data_bus[77]), .A2(n4724), .B1(
        i_data_bus[749]), .B2(n4088), .ZN(n4362) );
  AOI22D1BWP30P140LVT U4721 ( .A1(i_data_bus[109]), .A2(n4750), .B1(
        i_data_bus[877]), .B2(n4743), .ZN(n4361) );
  ND4D1BWP30P140LVT U4722 ( .A1(n4364), .A2(n4363), .A3(n4362), .A4(n4361), 
        .ZN(n4380) );
  AOI22D1BWP30P140LVT U4723 ( .A1(i_data_bus[589]), .A2(n4742), .B1(
        i_data_bus[685]), .B2(n4075), .ZN(n4368) );
  AOI22D1BWP30P140LVT U4724 ( .A1(i_data_bus[365]), .A2(n4739), .B1(
        i_data_bus[781]), .B2(n4721), .ZN(n4367) );
  AOI22D1BWP30P140LVT U4725 ( .A1(i_data_bus[621]), .A2(n4733), .B1(
        i_data_bus[301]), .B2(n4741), .ZN(n4366) );
  AOI22D1BWP30P140LVT U4726 ( .A1(i_data_bus[237]), .A2(n4749), .B1(
        i_data_bus[653]), .B2(n4730), .ZN(n4365) );
  ND4D1BWP30P140LVT U4727 ( .A1(n4368), .A2(n4367), .A3(n4366), .A4(n4365), 
        .ZN(n4379) );
  AOI22D1BWP30P140LVT U4728 ( .A1(i_data_bus[397]), .A2(n4752), .B1(
        i_data_bus[429]), .B2(n4732), .ZN(n4372) );
  AOI22D1BWP30P140LVT U4729 ( .A1(i_data_bus[845]), .A2(n4096), .B1(
        i_data_bus[813]), .B2(n4076), .ZN(n4371) );
  AOI22D1BWP30P140LVT U4730 ( .A1(i_data_bus[45]), .A2(n4740), .B1(
        i_data_bus[173]), .B2(n4738), .ZN(n4370) );
  AOI22D1BWP30P140LVT U4731 ( .A1(i_data_bus[525]), .A2(n4722), .B1(
        i_data_bus[269]), .B2(n4731), .ZN(n4369) );
  ND4D1BWP30P140LVT U4732 ( .A1(n4372), .A2(n4371), .A3(n4370), .A4(n4369), 
        .ZN(n4378) );
  AOI22D1BWP30P140LVT U4733 ( .A1(i_data_bus[333]), .A2(n4729), .B1(
        i_data_bus[717]), .B2(n4753), .ZN(n4376) );
  AOI22D1BWP30P140LVT U4734 ( .A1(i_data_bus[13]), .A2(n4097), .B1(
        i_data_bus[461]), .B2(n4751), .ZN(n4375) );
  AOI22D1BWP30P140LVT U4735 ( .A1(i_data_bus[557]), .A2(n4723), .B1(
        i_data_bus[205]), .B2(n4744), .ZN(n4374) );
  AOI22D1BWP30P140LVT U4736 ( .A1(i_data_bus[493]), .A2(n4111), .B1(
        i_data_bus[141]), .B2(n4108), .ZN(n4373) );
  ND4D1BWP30P140LVT U4737 ( .A1(n4376), .A2(n4375), .A3(n4374), .A4(n4373), 
        .ZN(n4377) );
  OR4D1BWP30P140LVT U4738 ( .A1(n4380), .A2(n4379), .A3(n4378), .A4(n4377), 
        .Z(o_data_bus[205]) );
  AOI22D1BWP30P140LVT U4739 ( .A1(i_data_bus[1006]), .A2(n4066), .B1(
        i_data_bus[974]), .B2(n4068), .ZN(n4384) );
  AOI22D1BWP30P140LVT U4740 ( .A1(i_data_bus[910]), .A2(n4073), .B1(
        i_data_bus[942]), .B2(n4070), .ZN(n4383) );
  AOI22D1BWP30P140LVT U4741 ( .A1(i_data_bus[46]), .A2(n4740), .B1(
        i_data_bus[206]), .B2(n4744), .ZN(n4382) );
  AOI22D1BWP30P140LVT U4742 ( .A1(i_data_bus[430]), .A2(n4732), .B1(
        i_data_bus[750]), .B2(n4088), .ZN(n4381) );
  ND4D1BWP30P140LVT U4743 ( .A1(n4384), .A2(n4383), .A3(n4382), .A4(n4381), 
        .ZN(n4400) );
  AOI22D1BWP30P140LVT U4744 ( .A1(i_data_bus[302]), .A2(n4741), .B1(
        i_data_bus[782]), .B2(n4721), .ZN(n4388) );
  AOI22D1BWP30P140LVT U4745 ( .A1(i_data_bus[590]), .A2(n4742), .B1(
        i_data_bus[558]), .B2(n4723), .ZN(n4387) );
  AOI22D1BWP30P140LVT U4746 ( .A1(i_data_bus[174]), .A2(n4738), .B1(
        i_data_bus[686]), .B2(n4075), .ZN(n4386) );
  AOI22D1BWP30P140LVT U4747 ( .A1(i_data_bus[622]), .A2(n4733), .B1(
        i_data_bus[238]), .B2(n4749), .ZN(n4385) );
  ND4D1BWP30P140LVT U4748 ( .A1(n4388), .A2(n4387), .A3(n4386), .A4(n4385), 
        .ZN(n4399) );
  AOI22D1BWP30P140LVT U4749 ( .A1(i_data_bus[78]), .A2(n4724), .B1(
        i_data_bus[366]), .B2(n4739), .ZN(n4392) );
  AOI22D1BWP30P140LVT U4750 ( .A1(i_data_bus[526]), .A2(n4722), .B1(
        i_data_bus[334]), .B2(n4729), .ZN(n4391) );
  AOI22D1BWP30P140LVT U4751 ( .A1(i_data_bus[14]), .A2(n4097), .B1(
        i_data_bus[270]), .B2(n4731), .ZN(n4390) );
  AOI22D1BWP30P140LVT U4752 ( .A1(i_data_bus[462]), .A2(n4751), .B1(
        i_data_bus[846]), .B2(n4096), .ZN(n4389) );
  ND4D1BWP30P140LVT U4753 ( .A1(n4392), .A2(n4391), .A3(n4390), .A4(n4389), 
        .ZN(n4398) );
  AOI22D1BWP30P140LVT U4754 ( .A1(i_data_bus[110]), .A2(n4750), .B1(
        i_data_bus[398]), .B2(n4752), .ZN(n4396) );
  AOI22D1BWP30P140LVT U4755 ( .A1(i_data_bus[814]), .A2(n4076), .B1(
        i_data_bus[878]), .B2(n4743), .ZN(n4395) );
  AOI22D1BWP30P140LVT U4756 ( .A1(i_data_bus[494]), .A2(n4111), .B1(
        i_data_bus[654]), .B2(n4730), .ZN(n4394) );
  AOI22D1BWP30P140LVT U4757 ( .A1(i_data_bus[142]), .A2(n4108), .B1(
        i_data_bus[718]), .B2(n4753), .ZN(n4393) );
  ND4D1BWP30P140LVT U4758 ( .A1(n4396), .A2(n4395), .A3(n4394), .A4(n4393), 
        .ZN(n4397) );
  OR4D1BWP30P140LVT U4759 ( .A1(n4400), .A2(n4399), .A3(n4398), .A4(n4397), 
        .Z(o_data_bus[206]) );
  AOI22D1BWP30P140LVT U4760 ( .A1(i_data_bus[1007]), .A2(n4066), .B1(
        i_data_bus[943]), .B2(n4070), .ZN(n4404) );
  AOI22D1BWP30P140LVT U4761 ( .A1(i_data_bus[975]), .A2(n4068), .B1(
        i_data_bus[911]), .B2(n4073), .ZN(n4403) );
  AOI22D1BWP30P140LVT U4762 ( .A1(i_data_bus[111]), .A2(n4750), .B1(
        i_data_bus[335]), .B2(n4729), .ZN(n4402) );
  AOI22D1BWP30P140LVT U4763 ( .A1(i_data_bus[271]), .A2(n4731), .B1(
        i_data_bus[815]), .B2(n4076), .ZN(n4401) );
  ND4D1BWP30P140LVT U4764 ( .A1(n4404), .A2(n4403), .A3(n4402), .A4(n4401), 
        .ZN(n4420) );
  AOI22D1BWP30P140LVT U4765 ( .A1(i_data_bus[47]), .A2(n4740), .B1(
        i_data_bus[207]), .B2(n4744), .ZN(n4408) );
  AOI22D1BWP30P140LVT U4766 ( .A1(i_data_bus[79]), .A2(n4724), .B1(
        i_data_bus[431]), .B2(n4732), .ZN(n4407) );
  AOI22D1BWP30P140LVT U4767 ( .A1(i_data_bus[847]), .A2(n4096), .B1(
        i_data_bus[143]), .B2(n4108), .ZN(n4406) );
  AOI22D1BWP30P140LVT U4768 ( .A1(i_data_bus[15]), .A2(n4097), .B1(
        i_data_bus[175]), .B2(n4738), .ZN(n4405) );
  ND4D1BWP30P140LVT U4769 ( .A1(n4408), .A2(n4407), .A3(n4406), .A4(n4405), 
        .ZN(n4419) );
  AOI22D1BWP30P140LVT U4770 ( .A1(i_data_bus[463]), .A2(n4751), .B1(
        i_data_bus[399]), .B2(n4752), .ZN(n4412) );
  AOI22D1BWP30P140LVT U4771 ( .A1(i_data_bus[527]), .A2(n4722), .B1(
        i_data_bus[623]), .B2(n4733), .ZN(n4411) );
  AOI22D1BWP30P140LVT U4772 ( .A1(i_data_bus[559]), .A2(n4723), .B1(
        i_data_bus[303]), .B2(n4741), .ZN(n4410) );
  AOI22D1BWP30P140LVT U4773 ( .A1(i_data_bus[719]), .A2(n4753), .B1(
        i_data_bus[239]), .B2(n4749), .ZN(n4409) );
  ND4D1BWP30P140LVT U4774 ( .A1(n4412), .A2(n4411), .A3(n4410), .A4(n4409), 
        .ZN(n4418) );
  AOI22D1BWP30P140LVT U4775 ( .A1(i_data_bus[655]), .A2(n4730), .B1(
        i_data_bus[783]), .B2(n4721), .ZN(n4416) );
  AOI22D1BWP30P140LVT U4776 ( .A1(i_data_bus[495]), .A2(n4111), .B1(
        i_data_bus[879]), .B2(n4743), .ZN(n4415) );
  AOI22D1BWP30P140LVT U4777 ( .A1(i_data_bus[751]), .A2(n4088), .B1(
        i_data_bus[687]), .B2(n4075), .ZN(n4414) );
  AOI22D1BWP30P140LVT U4778 ( .A1(i_data_bus[591]), .A2(n4742), .B1(
        i_data_bus[367]), .B2(n4739), .ZN(n4413) );
  ND4D1BWP30P140LVT U4779 ( .A1(n4416), .A2(n4415), .A3(n4414), .A4(n4413), 
        .ZN(n4417) );
  OR4D1BWP30P140LVT U4780 ( .A1(n4420), .A2(n4419), .A3(n4418), .A4(n4417), 
        .Z(o_data_bus[207]) );
  AOI22D1BWP30P140LVT U4781 ( .A1(i_data_bus[944]), .A2(n4070), .B1(
        i_data_bus[976]), .B2(n4068), .ZN(n4424) );
  AOI22D1BWP30P140LVT U4782 ( .A1(i_data_bus[912]), .A2(n4073), .B1(
        i_data_bus[1008]), .B2(n4066), .ZN(n4423) );
  AOI22D1BWP30P140LVT U4783 ( .A1(i_data_bus[496]), .A2(n4111), .B1(
        i_data_bus[720]), .B2(n4753), .ZN(n4422) );
  AOI22D1BWP30P140LVT U4784 ( .A1(i_data_bus[528]), .A2(n4722), .B1(
        i_data_bus[144]), .B2(n4108), .ZN(n4421) );
  ND4D1BWP30P140LVT U4785 ( .A1(n4424), .A2(n4423), .A3(n4422), .A4(n4421), 
        .ZN(n4440) );
  AOI22D1BWP30P140LVT U4786 ( .A1(i_data_bus[80]), .A2(n4724), .B1(
        i_data_bus[112]), .B2(n4750), .ZN(n4428) );
  AOI22D1BWP30P140LVT U4787 ( .A1(i_data_bus[304]), .A2(n4741), .B1(
        i_data_bus[208]), .B2(n4744), .ZN(n4427) );
  AOI22D1BWP30P140LVT U4788 ( .A1(i_data_bus[784]), .A2(n4721), .B1(
        i_data_bus[400]), .B2(n4752), .ZN(n4426) );
  AOI22D1BWP30P140LVT U4789 ( .A1(i_data_bus[560]), .A2(n4723), .B1(
        i_data_bus[880]), .B2(n4743), .ZN(n4425) );
  ND4D1BWP30P140LVT U4790 ( .A1(n4428), .A2(n4427), .A3(n4426), .A4(n4425), 
        .ZN(n4439) );
  AOI22D1BWP30P140LVT U4791 ( .A1(i_data_bus[432]), .A2(n4732), .B1(
        i_data_bus[752]), .B2(n4088), .ZN(n4432) );
  AOI22D1BWP30P140LVT U4792 ( .A1(i_data_bus[656]), .A2(n4730), .B1(
        i_data_bus[176]), .B2(n4738), .ZN(n4431) );
  AOI22D1BWP30P140LVT U4793 ( .A1(i_data_bus[624]), .A2(n4733), .B1(
        i_data_bus[816]), .B2(n4076), .ZN(n4430) );
  AOI22D1BWP30P140LVT U4794 ( .A1(i_data_bus[336]), .A2(n4729), .B1(
        i_data_bus[848]), .B2(n4096), .ZN(n4429) );
  ND4D1BWP30P140LVT U4795 ( .A1(n4432), .A2(n4431), .A3(n4430), .A4(n4429), 
        .ZN(n4438) );
  AOI22D1BWP30P140LVT U4796 ( .A1(i_data_bus[592]), .A2(n4742), .B1(
        i_data_bus[688]), .B2(n4075), .ZN(n4436) );
  AOI22D1BWP30P140LVT U4797 ( .A1(i_data_bus[16]), .A2(n4097), .B1(
        i_data_bus[464]), .B2(n4751), .ZN(n4435) );
  AOI22D1BWP30P140LVT U4798 ( .A1(i_data_bus[48]), .A2(n4740), .B1(
        i_data_bus[368]), .B2(n4739), .ZN(n4434) );
  AOI22D1BWP30P140LVT U4799 ( .A1(i_data_bus[272]), .A2(n4731), .B1(
        i_data_bus[240]), .B2(n4749), .ZN(n4433) );
  ND4D1BWP30P140LVT U4800 ( .A1(n4436), .A2(n4435), .A3(n4434), .A4(n4433), 
        .ZN(n4437) );
  OR4D1BWP30P140LVT U4801 ( .A1(n4440), .A2(n4439), .A3(n4438), .A4(n4437), 
        .Z(o_data_bus[208]) );
  AOI22D1BWP30P140LVT U4802 ( .A1(i_data_bus[1009]), .A2(n4066), .B1(
        i_data_bus[913]), .B2(n4073), .ZN(n4444) );
  AOI22D1BWP30P140LVT U4803 ( .A1(i_data_bus[945]), .A2(n4070), .B1(
        i_data_bus[977]), .B2(n4068), .ZN(n4443) );
  AOI22D1BWP30P140LVT U4804 ( .A1(i_data_bus[49]), .A2(n4740), .B1(
        i_data_bus[145]), .B2(n4108), .ZN(n4442) );
  AOI22D1BWP30P140LVT U4805 ( .A1(i_data_bus[401]), .A2(n4752), .B1(
        i_data_bus[209]), .B2(n4744), .ZN(n4441) );
  ND4D1BWP30P140LVT U4806 ( .A1(n4444), .A2(n4443), .A3(n4442), .A4(n4441), 
        .ZN(n4460) );
  AOI22D1BWP30P140LVT U4807 ( .A1(i_data_bus[721]), .A2(n4753), .B1(
        i_data_bus[657]), .B2(n4730), .ZN(n4448) );
  AOI22D1BWP30P140LVT U4808 ( .A1(i_data_bus[753]), .A2(n4088), .B1(
        i_data_bus[465]), .B2(n4751), .ZN(n4447) );
  AOI22D1BWP30P140LVT U4809 ( .A1(i_data_bus[273]), .A2(n4731), .B1(
        i_data_bus[369]), .B2(n4739), .ZN(n4446) );
  AOI22D1BWP30P140LVT U4810 ( .A1(i_data_bus[529]), .A2(n4722), .B1(
        i_data_bus[433]), .B2(n4732), .ZN(n4445) );
  ND4D1BWP30P140LVT U4811 ( .A1(n4448), .A2(n4447), .A3(n4446), .A4(n4445), 
        .ZN(n4459) );
  AOI22D1BWP30P140LVT U4812 ( .A1(i_data_bus[881]), .A2(n4743), .B1(
        i_data_bus[305]), .B2(n4741), .ZN(n4452) );
  AOI22D1BWP30P140LVT U4813 ( .A1(i_data_bus[241]), .A2(n4749), .B1(
        i_data_bus[817]), .B2(n4076), .ZN(n4451) );
  AOI22D1BWP30P140LVT U4814 ( .A1(i_data_bus[625]), .A2(n4733), .B1(
        i_data_bus[81]), .B2(n4724), .ZN(n4450) );
  AOI22D1BWP30P140LVT U4815 ( .A1(i_data_bus[113]), .A2(n4750), .B1(
        i_data_bus[177]), .B2(n4738), .ZN(n4449) );
  ND4D1BWP30P140LVT U4816 ( .A1(n4452), .A2(n4451), .A3(n4450), .A4(n4449), 
        .ZN(n4458) );
  AOI22D1BWP30P140LVT U4817 ( .A1(i_data_bus[689]), .A2(n4075), .B1(
        i_data_bus[785]), .B2(n4721), .ZN(n4456) );
  AOI22D1BWP30P140LVT U4818 ( .A1(i_data_bus[17]), .A2(n4097), .B1(
        i_data_bus[497]), .B2(n4111), .ZN(n4455) );
  AOI22D1BWP30P140LVT U4819 ( .A1(i_data_bus[593]), .A2(n4742), .B1(
        i_data_bus[849]), .B2(n4096), .ZN(n4454) );
  AOI22D1BWP30P140LVT U4820 ( .A1(i_data_bus[561]), .A2(n4723), .B1(
        i_data_bus[337]), .B2(n4729), .ZN(n4453) );
  ND4D1BWP30P140LVT U4821 ( .A1(n4456), .A2(n4455), .A3(n4454), .A4(n4453), 
        .ZN(n4457) );
  OR4D1BWP30P140LVT U4822 ( .A1(n4460), .A2(n4459), .A3(n4458), .A4(n4457), 
        .Z(o_data_bus[209]) );
  AOI22D1BWP30P140LVT U4823 ( .A1(i_data_bus[978]), .A2(n4068), .B1(
        i_data_bus[914]), .B2(n4073), .ZN(n4464) );
  AOI22D1BWP30P140LVT U4824 ( .A1(i_data_bus[1010]), .A2(n4066), .B1(
        i_data_bus[946]), .B2(n4070), .ZN(n4463) );
  AOI22D1BWP30P140LVT U4825 ( .A1(i_data_bus[370]), .A2(n4739), .B1(
        i_data_bus[434]), .B2(n4732), .ZN(n4462) );
  AOI22D1BWP30P140LVT U4826 ( .A1(i_data_bus[626]), .A2(n4733), .B1(
        i_data_bus[146]), .B2(n4108), .ZN(n4461) );
  ND4D1BWP30P140LVT U4827 ( .A1(n4464), .A2(n4463), .A3(n4462), .A4(n4461), 
        .ZN(n4480) );
  AOI22D1BWP30P140LVT U4828 ( .A1(i_data_bus[882]), .A2(n4743), .B1(
        i_data_bus[690]), .B2(n4075), .ZN(n4468) );
  AOI22D1BWP30P140LVT U4829 ( .A1(i_data_bus[594]), .A2(n4742), .B1(
        i_data_bus[18]), .B2(n4097), .ZN(n4467) );
  AOI22D1BWP30P140LVT U4830 ( .A1(i_data_bus[402]), .A2(n4752), .B1(
        i_data_bus[498]), .B2(n4111), .ZN(n4466) );
  AOI22D1BWP30P140LVT U4831 ( .A1(i_data_bus[850]), .A2(n4096), .B1(
        i_data_bus[274]), .B2(n4731), .ZN(n4465) );
  ND4D1BWP30P140LVT U4832 ( .A1(n4468), .A2(n4467), .A3(n4466), .A4(n4465), 
        .ZN(n4479) );
  AOI22D1BWP30P140LVT U4833 ( .A1(i_data_bus[50]), .A2(n4740), .B1(
        i_data_bus[114]), .B2(n4750), .ZN(n4472) );
  AOI22D1BWP30P140LVT U4834 ( .A1(i_data_bus[82]), .A2(n4724), .B1(
        i_data_bus[658]), .B2(n4730), .ZN(n4471) );
  AOI22D1BWP30P140LVT U4835 ( .A1(i_data_bus[562]), .A2(n4723), .B1(
        i_data_bus[210]), .B2(n4744), .ZN(n4470) );
  AOI22D1BWP30P140LVT U4836 ( .A1(i_data_bus[178]), .A2(n4738), .B1(
        i_data_bus[754]), .B2(n4088), .ZN(n4469) );
  ND4D1BWP30P140LVT U4837 ( .A1(n4472), .A2(n4471), .A3(n4470), .A4(n4469), 
        .ZN(n4478) );
  AOI22D1BWP30P140LVT U4838 ( .A1(i_data_bus[242]), .A2(n4749), .B1(
        i_data_bus[306]), .B2(n4741), .ZN(n4476) );
  AOI22D1BWP30P140LVT U4839 ( .A1(i_data_bus[818]), .A2(n4076), .B1(
        i_data_bus[338]), .B2(n4729), .ZN(n4475) );
  AOI22D1BWP30P140LVT U4840 ( .A1(i_data_bus[530]), .A2(n4722), .B1(
        i_data_bus[722]), .B2(n4753), .ZN(n4474) );
  AOI22D1BWP30P140LVT U4841 ( .A1(i_data_bus[466]), .A2(n4751), .B1(
        i_data_bus[786]), .B2(n4721), .ZN(n4473) );
  ND4D1BWP30P140LVT U4842 ( .A1(n4476), .A2(n4475), .A3(n4474), .A4(n4473), 
        .ZN(n4477) );
  OR4D1BWP30P140LVT U4843 ( .A1(n4480), .A2(n4479), .A3(n4478), .A4(n4477), 
        .Z(o_data_bus[210]) );
  AOI22D1BWP30P140LVT U4844 ( .A1(i_data_bus[979]), .A2(n4068), .B1(
        i_data_bus[915]), .B2(n4073), .ZN(n4484) );
  AOI22D1BWP30P140LVT U4845 ( .A1(i_data_bus[1011]), .A2(n4066), .B1(
        i_data_bus[947]), .B2(n4070), .ZN(n4483) );
  AOI22D1BWP30P140LVT U4846 ( .A1(i_data_bus[211]), .A2(n4744), .B1(
        i_data_bus[307]), .B2(n4741), .ZN(n4482) );
  AOI22D1BWP30P140LVT U4847 ( .A1(i_data_bus[755]), .A2(n4088), .B1(
        i_data_bus[659]), .B2(n4730), .ZN(n4481) );
  ND4D1BWP30P140LVT U4848 ( .A1(n4484), .A2(n4483), .A3(n4482), .A4(n4481), 
        .ZN(n4500) );
  AOI22D1BWP30P140LVT U4849 ( .A1(i_data_bus[531]), .A2(n4722), .B1(
        i_data_bus[19]), .B2(n4097), .ZN(n4488) );
  AOI22D1BWP30P140LVT U4850 ( .A1(i_data_bus[51]), .A2(n4740), .B1(
        i_data_bus[595]), .B2(n4742), .ZN(n4487) );
  AOI22D1BWP30P140LVT U4851 ( .A1(i_data_bus[563]), .A2(n4723), .B1(
        i_data_bus[787]), .B2(n4721), .ZN(n4486) );
  AOI22D1BWP30P140LVT U4852 ( .A1(i_data_bus[627]), .A2(n4733), .B1(
        i_data_bus[723]), .B2(n4753), .ZN(n4485) );
  ND4D1BWP30P140LVT U4853 ( .A1(n4488), .A2(n4487), .A3(n4486), .A4(n4485), 
        .ZN(n4499) );
  AOI22D1BWP30P140LVT U4854 ( .A1(i_data_bus[115]), .A2(n4750), .B1(
        i_data_bus[275]), .B2(n4731), .ZN(n4492) );
  AOI22D1BWP30P140LVT U4855 ( .A1(i_data_bus[371]), .A2(n4739), .B1(
        i_data_bus[467]), .B2(n4751), .ZN(n4491) );
  AOI22D1BWP30P140LVT U4856 ( .A1(i_data_bus[243]), .A2(n4749), .B1(
        i_data_bus[819]), .B2(n4076), .ZN(n4490) );
  AOI22D1BWP30P140LVT U4857 ( .A1(i_data_bus[339]), .A2(n4729), .B1(
        i_data_bus[435]), .B2(n4732), .ZN(n4489) );
  ND4D1BWP30P140LVT U4858 ( .A1(n4492), .A2(n4491), .A3(n4490), .A4(n4489), 
        .ZN(n4498) );
  AOI22D1BWP30P140LVT U4859 ( .A1(i_data_bus[883]), .A2(n4743), .B1(
        i_data_bus[691]), .B2(n4075), .ZN(n4496) );
  AOI22D1BWP30P140LVT U4860 ( .A1(i_data_bus[403]), .A2(n4752), .B1(
        i_data_bus[851]), .B2(n4096), .ZN(n4495) );
  AOI22D1BWP30P140LVT U4861 ( .A1(i_data_bus[83]), .A2(n4724), .B1(
        i_data_bus[147]), .B2(n4108), .ZN(n4494) );
  AOI22D1BWP30P140LVT U4862 ( .A1(i_data_bus[179]), .A2(n4738), .B1(
        i_data_bus[499]), .B2(n4111), .ZN(n4493) );
  ND4D1BWP30P140LVT U4863 ( .A1(n4496), .A2(n4495), .A3(n4494), .A4(n4493), 
        .ZN(n4497) );
  OR4D1BWP30P140LVT U4864 ( .A1(n4500), .A2(n4499), .A3(n4498), .A4(n4497), 
        .Z(o_data_bus[211]) );
  AOI22D1BWP30P140LVT U4865 ( .A1(i_data_bus[980]), .A2(n4068), .B1(
        i_data_bus[916]), .B2(n4073), .ZN(n4504) );
  AOI22D1BWP30P140LVT U4866 ( .A1(i_data_bus[1012]), .A2(n4066), .B1(
        i_data_bus[948]), .B2(n4070), .ZN(n4503) );
  AOI22D1BWP30P140LVT U4867 ( .A1(i_data_bus[788]), .A2(n4721), .B1(
        i_data_bus[372]), .B2(n4739), .ZN(n4502) );
  AOI22D1BWP30P140LVT U4868 ( .A1(i_data_bus[212]), .A2(n4744), .B1(
        i_data_bus[660]), .B2(n4730), .ZN(n4501) );
  ND4D1BWP30P140LVT U4869 ( .A1(n4504), .A2(n4503), .A3(n4502), .A4(n4501), 
        .ZN(n4520) );
  AOI22D1BWP30P140LVT U4870 ( .A1(i_data_bus[628]), .A2(n4733), .B1(
        i_data_bus[436]), .B2(n4732), .ZN(n4508) );
  AOI22D1BWP30P140LVT U4871 ( .A1(i_data_bus[596]), .A2(n4742), .B1(
        i_data_bus[852]), .B2(n4096), .ZN(n4507) );
  AOI22D1BWP30P140LVT U4872 ( .A1(i_data_bus[532]), .A2(n4722), .B1(
        i_data_bus[884]), .B2(n4743), .ZN(n4506) );
  AOI22D1BWP30P140LVT U4873 ( .A1(i_data_bus[52]), .A2(n4740), .B1(
        i_data_bus[276]), .B2(n4731), .ZN(n4505) );
  ND4D1BWP30P140LVT U4874 ( .A1(n4508), .A2(n4507), .A3(n4506), .A4(n4505), 
        .ZN(n4519) );
  AOI22D1BWP30P140LVT U4875 ( .A1(i_data_bus[756]), .A2(n4088), .B1(
        i_data_bus[692]), .B2(n4075), .ZN(n4512) );
  AOI22D1BWP30P140LVT U4876 ( .A1(i_data_bus[20]), .A2(n4097), .B1(
        i_data_bus[820]), .B2(n4076), .ZN(n4511) );
  AOI22D1BWP30P140LVT U4877 ( .A1(i_data_bus[84]), .A2(n4724), .B1(
        i_data_bus[468]), .B2(n4751), .ZN(n4510) );
  AOI22D1BWP30P140LVT U4878 ( .A1(i_data_bus[244]), .A2(n4749), .B1(
        i_data_bus[308]), .B2(n4741), .ZN(n4509) );
  ND4D1BWP30P140LVT U4879 ( .A1(n4512), .A2(n4511), .A3(n4510), .A4(n4509), 
        .ZN(n4518) );
  AOI22D1BWP30P140LVT U4880 ( .A1(i_data_bus[116]), .A2(n4750), .B1(
        i_data_bus[180]), .B2(n4738), .ZN(n4516) );
  AOI22D1BWP30P140LVT U4881 ( .A1(i_data_bus[724]), .A2(n4753), .B1(
        i_data_bus[500]), .B2(n4111), .ZN(n4515) );
  AOI22D1BWP30P140LVT U4882 ( .A1(i_data_bus[404]), .A2(n4752), .B1(
        i_data_bus[148]), .B2(n4108), .ZN(n4514) );
  AOI22D1BWP30P140LVT U4883 ( .A1(i_data_bus[564]), .A2(n4723), .B1(
        i_data_bus[340]), .B2(n4729), .ZN(n4513) );
  ND4D1BWP30P140LVT U4884 ( .A1(n4516), .A2(n4515), .A3(n4514), .A4(n4513), 
        .ZN(n4517) );
  OR4D1BWP30P140LVT U4885 ( .A1(n4520), .A2(n4519), .A3(n4518), .A4(n4517), 
        .Z(o_data_bus[212]) );
  AOI22D1BWP30P140LVT U4886 ( .A1(i_data_bus[917]), .A2(n4073), .B1(
        i_data_bus[1013]), .B2(n4066), .ZN(n4524) );
  AOI22D1BWP30P140LVT U4887 ( .A1(i_data_bus[949]), .A2(n4070), .B1(
        i_data_bus[981]), .B2(n4068), .ZN(n4523) );
  AOI22D1BWP30P140LVT U4888 ( .A1(i_data_bus[501]), .A2(n4111), .B1(
        i_data_bus[373]), .B2(n4739), .ZN(n4522) );
  AOI22D1BWP30P140LVT U4889 ( .A1(i_data_bus[565]), .A2(n4723), .B1(
        i_data_bus[853]), .B2(n4096), .ZN(n4521) );
  ND4D1BWP30P140LVT U4890 ( .A1(n4524), .A2(n4523), .A3(n4522), .A4(n4521), 
        .ZN(n4540) );
  AOI22D1BWP30P140LVT U4891 ( .A1(i_data_bus[53]), .A2(n4740), .B1(
        i_data_bus[885]), .B2(n4743), .ZN(n4528) );
  AOI22D1BWP30P140LVT U4892 ( .A1(i_data_bus[629]), .A2(n4733), .B1(
        i_data_bus[533]), .B2(n4722), .ZN(n4527) );
  AOI22D1BWP30P140LVT U4893 ( .A1(i_data_bus[597]), .A2(n4742), .B1(
        i_data_bus[277]), .B2(n4731), .ZN(n4526) );
  AOI22D1BWP30P140LVT U4894 ( .A1(i_data_bus[341]), .A2(n4729), .B1(
        i_data_bus[309]), .B2(n4741), .ZN(n4525) );
  ND4D1BWP30P140LVT U4895 ( .A1(n4528), .A2(n4527), .A3(n4526), .A4(n4525), 
        .ZN(n4539) );
  AOI22D1BWP30P140LVT U4896 ( .A1(i_data_bus[213]), .A2(n4744), .B1(
        i_data_bus[469]), .B2(n4751), .ZN(n4532) );
  AOI22D1BWP30P140LVT U4897 ( .A1(i_data_bus[789]), .A2(n4721), .B1(
        i_data_bus[149]), .B2(n4108), .ZN(n4531) );
  AOI22D1BWP30P140LVT U4898 ( .A1(i_data_bus[85]), .A2(n4724), .B1(
        i_data_bus[661]), .B2(n4730), .ZN(n4530) );
  AOI22D1BWP30P140LVT U4899 ( .A1(i_data_bus[21]), .A2(n4097), .B1(
        i_data_bus[725]), .B2(n4753), .ZN(n4529) );
  ND4D1BWP30P140LVT U4900 ( .A1(n4532), .A2(n4531), .A3(n4530), .A4(n4529), 
        .ZN(n4538) );
  AOI22D1BWP30P140LVT U4901 ( .A1(i_data_bus[757]), .A2(n4088), .B1(
        i_data_bus[821]), .B2(n4076), .ZN(n4536) );
  AOI22D1BWP30P140LVT U4902 ( .A1(i_data_bus[245]), .A2(n4749), .B1(
        i_data_bus[405]), .B2(n4752), .ZN(n4535) );
  AOI22D1BWP30P140LVT U4903 ( .A1(i_data_bus[117]), .A2(n4750), .B1(
        i_data_bus[437]), .B2(n4732), .ZN(n4534) );
  AOI22D1BWP30P140LVT U4904 ( .A1(i_data_bus[181]), .A2(n4738), .B1(
        i_data_bus[693]), .B2(n4075), .ZN(n4533) );
  ND4D1BWP30P140LVT U4905 ( .A1(n4536), .A2(n4535), .A3(n4534), .A4(n4533), 
        .ZN(n4537) );
  OR4D1BWP30P140LVT U4906 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), 
        .Z(o_data_bus[213]) );
  AOI22D1BWP30P140LVT U4907 ( .A1(i_data_bus[1014]), .A2(n4066), .B1(
        i_data_bus[918]), .B2(n4073), .ZN(n4544) );
  AOI22D1BWP30P140LVT U4908 ( .A1(i_data_bus[950]), .A2(n4070), .B1(
        i_data_bus[982]), .B2(n4068), .ZN(n4543) );
  AOI22D1BWP30P140LVT U4909 ( .A1(i_data_bus[822]), .A2(n4076), .B1(
        i_data_bus[246]), .B2(n4749), .ZN(n4542) );
  AOI22D1BWP30P140LVT U4910 ( .A1(i_data_bus[374]), .A2(n4739), .B1(
        i_data_bus[150]), .B2(n4108), .ZN(n4541) );
  ND4D1BWP30P140LVT U4911 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), 
        .ZN(n4560) );
  AOI22D1BWP30P140LVT U4912 ( .A1(i_data_bus[406]), .A2(n4752), .B1(
        i_data_bus[662]), .B2(n4730), .ZN(n4548) );
  AOI22D1BWP30P140LVT U4913 ( .A1(i_data_bus[630]), .A2(n4733), .B1(
        i_data_bus[214]), .B2(n4744), .ZN(n4547) );
  AOI22D1BWP30P140LVT U4914 ( .A1(i_data_bus[118]), .A2(n4750), .B1(
        i_data_bus[310]), .B2(n4741), .ZN(n4546) );
  AOI22D1BWP30P140LVT U4915 ( .A1(i_data_bus[598]), .A2(n4742), .B1(
        i_data_bus[854]), .B2(n4096), .ZN(n4545) );
  ND4D1BWP30P140LVT U4916 ( .A1(n4548), .A2(n4547), .A3(n4546), .A4(n4545), 
        .ZN(n4559) );
  AOI22D1BWP30P140LVT U4917 ( .A1(i_data_bus[54]), .A2(n4740), .B1(
        i_data_bus[566]), .B2(n4723), .ZN(n4552) );
  AOI22D1BWP30P140LVT U4918 ( .A1(i_data_bus[502]), .A2(n4111), .B1(
        i_data_bus[470]), .B2(n4751), .ZN(n4551) );
  AOI22D1BWP30P140LVT U4919 ( .A1(i_data_bus[726]), .A2(n4753), .B1(
        i_data_bus[278]), .B2(n4731), .ZN(n4550) );
  AOI22D1BWP30P140LVT U4920 ( .A1(i_data_bus[22]), .A2(n4097), .B1(
        i_data_bus[342]), .B2(n4729), .ZN(n4549) );
  ND4D1BWP30P140LVT U4921 ( .A1(n4552), .A2(n4551), .A3(n4550), .A4(n4549), 
        .ZN(n4558) );
  AOI22D1BWP30P140LVT U4922 ( .A1(i_data_bus[86]), .A2(n4724), .B1(
        i_data_bus[886]), .B2(n4743), .ZN(n4556) );
  AOI22D1BWP30P140LVT U4923 ( .A1(i_data_bus[534]), .A2(n4722), .B1(
        i_data_bus[438]), .B2(n4732), .ZN(n4555) );
  AOI22D1BWP30P140LVT U4924 ( .A1(i_data_bus[790]), .A2(n4721), .B1(
        i_data_bus[182]), .B2(n4738), .ZN(n4554) );
  AOI22D1BWP30P140LVT U4925 ( .A1(i_data_bus[694]), .A2(n4075), .B1(
        i_data_bus[758]), .B2(n4088), .ZN(n4553) );
  ND4D1BWP30P140LVT U4926 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), 
        .ZN(n4557) );
  OR4D1BWP30P140LVT U4927 ( .A1(n4560), .A2(n4559), .A3(n4558), .A4(n4557), 
        .Z(o_data_bus[214]) );
  AOI22D1BWP30P140LVT U4928 ( .A1(i_data_bus[951]), .A2(n4070), .B1(
        i_data_bus[919]), .B2(n4073), .ZN(n4564) );
  AOI22D1BWP30P140LVT U4929 ( .A1(i_data_bus[1015]), .A2(n4066), .B1(
        i_data_bus[983]), .B2(n4068), .ZN(n4563) );
  AOI22D1BWP30P140LVT U4930 ( .A1(i_data_bus[727]), .A2(n4753), .B1(
        i_data_bus[823]), .B2(n4076), .ZN(n4562) );
  AOI22D1BWP30P140LVT U4931 ( .A1(i_data_bus[535]), .A2(n4722), .B1(
        i_data_bus[151]), .B2(n4108), .ZN(n4561) );
  ND4D1BWP30P140LVT U4932 ( .A1(n4564), .A2(n4563), .A3(n4562), .A4(n4561), 
        .ZN(n4580) );
  AOI22D1BWP30P140LVT U4933 ( .A1(i_data_bus[503]), .A2(n4111), .B1(
        i_data_bus[407]), .B2(n4752), .ZN(n4568) );
  AOI22D1BWP30P140LVT U4934 ( .A1(i_data_bus[119]), .A2(n4750), .B1(
        i_data_bus[759]), .B2(n4088), .ZN(n4567) );
  AOI22D1BWP30P140LVT U4935 ( .A1(i_data_bus[695]), .A2(n4075), .B1(
        i_data_bus[663]), .B2(n4730), .ZN(n4566) );
  AOI22D1BWP30P140LVT U4936 ( .A1(i_data_bus[471]), .A2(n4751), .B1(
        i_data_bus[855]), .B2(n4096), .ZN(n4565) );
  ND4D1BWP30P140LVT U4937 ( .A1(n4568), .A2(n4567), .A3(n4566), .A4(n4565), 
        .ZN(n4579) );
  AOI22D1BWP30P140LVT U4938 ( .A1(i_data_bus[599]), .A2(n4742), .B1(
        i_data_bus[887]), .B2(n4743), .ZN(n4572) );
  AOI22D1BWP30P140LVT U4939 ( .A1(i_data_bus[311]), .A2(n4741), .B1(
        i_data_bus[343]), .B2(n4729), .ZN(n4571) );
  AOI22D1BWP30P140LVT U4940 ( .A1(i_data_bus[247]), .A2(n4749), .B1(
        i_data_bus[791]), .B2(n4721), .ZN(n4570) );
  AOI22D1BWP30P140LVT U4941 ( .A1(i_data_bus[23]), .A2(n4097), .B1(
        i_data_bus[567]), .B2(n4723), .ZN(n4569) );
  ND4D1BWP30P140LVT U4942 ( .A1(n4572), .A2(n4571), .A3(n4570), .A4(n4569), 
        .ZN(n4578) );
  AOI22D1BWP30P140LVT U4943 ( .A1(i_data_bus[87]), .A2(n4724), .B1(
        i_data_bus[183]), .B2(n4738), .ZN(n4576) );
  AOI22D1BWP30P140LVT U4944 ( .A1(i_data_bus[55]), .A2(n4740), .B1(
        i_data_bus[375]), .B2(n4739), .ZN(n4575) );
  AOI22D1BWP30P140LVT U4945 ( .A1(i_data_bus[279]), .A2(n4731), .B1(
        i_data_bus[215]), .B2(n4744), .ZN(n4574) );
  AOI22D1BWP30P140LVT U4946 ( .A1(i_data_bus[631]), .A2(n4733), .B1(
        i_data_bus[439]), .B2(n4732), .ZN(n4573) );
  ND4D1BWP30P140LVT U4947 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), 
        .ZN(n4577) );
  OR4D1BWP30P140LVT U4948 ( .A1(n4580), .A2(n4579), .A3(n4578), .A4(n4577), 
        .Z(o_data_bus[215]) );
  AOI22D1BWP30P140LVT U4949 ( .A1(i_data_bus[952]), .A2(n4070), .B1(
        i_data_bus[920]), .B2(n4073), .ZN(n4584) );
  AOI22D1BWP30P140LVT U4950 ( .A1(i_data_bus[984]), .A2(n4068), .B1(
        i_data_bus[1016]), .B2(n4066), .ZN(n4583) );
  AOI22D1BWP30P140LVT U4951 ( .A1(i_data_bus[600]), .A2(n4742), .B1(
        i_data_bus[472]), .B2(n4751), .ZN(n4582) );
  AOI22D1BWP30P140LVT U4952 ( .A1(i_data_bus[568]), .A2(n4723), .B1(
        i_data_bus[504]), .B2(n4111), .ZN(n4581) );
  ND4D1BWP30P140LVT U4953 ( .A1(n4584), .A2(n4583), .A3(n4582), .A4(n4581), 
        .ZN(n4600) );
  AOI22D1BWP30P140LVT U4954 ( .A1(i_data_bus[440]), .A2(n4732), .B1(
        i_data_bus[728]), .B2(n4753), .ZN(n4588) );
  AOI22D1BWP30P140LVT U4955 ( .A1(i_data_bus[632]), .A2(n4733), .B1(
        i_data_bus[88]), .B2(n4724), .ZN(n4587) );
  AOI22D1BWP30P140LVT U4956 ( .A1(i_data_bus[408]), .A2(n4752), .B1(
        i_data_bus[184]), .B2(n4738), .ZN(n4586) );
  AOI22D1BWP30P140LVT U4957 ( .A1(i_data_bus[856]), .A2(n4096), .B1(
        i_data_bus[824]), .B2(n4076), .ZN(n4585) );
  ND4D1BWP30P140LVT U4958 ( .A1(n4588), .A2(n4587), .A3(n4586), .A4(n4585), 
        .ZN(n4599) );
  AOI22D1BWP30P140LVT U4959 ( .A1(i_data_bus[120]), .A2(n4750), .B1(
        i_data_bus[280]), .B2(n4731), .ZN(n4592) );
  AOI22D1BWP30P140LVT U4960 ( .A1(i_data_bus[24]), .A2(n4097), .B1(
        i_data_bus[376]), .B2(n4739), .ZN(n4591) );
  AOI22D1BWP30P140LVT U4961 ( .A1(i_data_bus[536]), .A2(n4722), .B1(
        i_data_bus[792]), .B2(n4721), .ZN(n4590) );
  AOI22D1BWP30P140LVT U4962 ( .A1(i_data_bus[248]), .A2(n4749), .B1(
        i_data_bus[152]), .B2(n4108), .ZN(n4589) );
  ND4D1BWP30P140LVT U4963 ( .A1(n4592), .A2(n4591), .A3(n4590), .A4(n4589), 
        .ZN(n4598) );
  AOI22D1BWP30P140LVT U4964 ( .A1(i_data_bus[344]), .A2(n4729), .B1(
        i_data_bus[312]), .B2(n4741), .ZN(n4596) );
  AOI22D1BWP30P140LVT U4965 ( .A1(i_data_bus[56]), .A2(n4740), .B1(
        i_data_bus[696]), .B2(n4075), .ZN(n4595) );
  AOI22D1BWP30P140LVT U4966 ( .A1(i_data_bus[888]), .A2(n4743), .B1(
        i_data_bus[760]), .B2(n4088), .ZN(n4594) );
  AOI22D1BWP30P140LVT U4967 ( .A1(i_data_bus[664]), .A2(n4730), .B1(
        i_data_bus[216]), .B2(n4744), .ZN(n4593) );
  ND4D1BWP30P140LVT U4968 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), 
        .ZN(n4597) );
  OR4D1BWP30P140LVT U4969 ( .A1(n4600), .A2(n4599), .A3(n4598), .A4(n4597), 
        .Z(o_data_bus[216]) );
  AOI22D1BWP30P140LVT U4970 ( .A1(i_data_bus[1017]), .A2(n4066), .B1(
        i_data_bus[921]), .B2(n4073), .ZN(n4604) );
  AOI22D1BWP30P140LVT U4971 ( .A1(i_data_bus[985]), .A2(n4068), .B1(
        i_data_bus[953]), .B2(n4070), .ZN(n4603) );
  AOI22D1BWP30P140LVT U4972 ( .A1(i_data_bus[665]), .A2(n4730), .B1(
        i_data_bus[153]), .B2(n4108), .ZN(n4602) );
  AOI22D1BWP30P140LVT U4973 ( .A1(i_data_bus[601]), .A2(n4742), .B1(
        i_data_bus[281]), .B2(n4731), .ZN(n4601) );
  ND4D1BWP30P140LVT U4974 ( .A1(n4604), .A2(n4603), .A3(n4602), .A4(n4601), 
        .ZN(n4620) );
  AOI22D1BWP30P140LVT U4975 ( .A1(i_data_bus[761]), .A2(n4088), .B1(
        i_data_bus[505]), .B2(n4111), .ZN(n4608) );
  AOI22D1BWP30P140LVT U4976 ( .A1(i_data_bus[633]), .A2(n4733), .B1(
        i_data_bus[345]), .B2(n4729), .ZN(n4607) );
  AOI22D1BWP30P140LVT U4977 ( .A1(i_data_bus[729]), .A2(n4753), .B1(
        i_data_bus[441]), .B2(n4732), .ZN(n4606) );
  AOI22D1BWP30P140LVT U4978 ( .A1(i_data_bus[537]), .A2(n4722), .B1(
        i_data_bus[857]), .B2(n4096), .ZN(n4605) );
  ND4D1BWP30P140LVT U4979 ( .A1(n4608), .A2(n4607), .A3(n4606), .A4(n4605), 
        .ZN(n4619) );
  AOI22D1BWP30P140LVT U4980 ( .A1(i_data_bus[89]), .A2(n4724), .B1(
        i_data_bus[409]), .B2(n4752), .ZN(n4612) );
  AOI22D1BWP30P140LVT U4981 ( .A1(i_data_bus[25]), .A2(n4097), .B1(
        i_data_bus[313]), .B2(n4741), .ZN(n4611) );
  AOI22D1BWP30P140LVT U4982 ( .A1(i_data_bus[473]), .A2(n4751), .B1(
        i_data_bus[249]), .B2(n4749), .ZN(n4610) );
  AOI22D1BWP30P140LVT U4983 ( .A1(i_data_bus[793]), .A2(n4721), .B1(
        i_data_bus[377]), .B2(n4739), .ZN(n4609) );
  ND4D1BWP30P140LVT U4984 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n4609), 
        .ZN(n4618) );
  AOI22D1BWP30P140LVT U4985 ( .A1(i_data_bus[57]), .A2(n4740), .B1(
        i_data_bus[185]), .B2(n4738), .ZN(n4616) );
  AOI22D1BWP30P140LVT U4986 ( .A1(i_data_bus[697]), .A2(n4075), .B1(
        i_data_bus[217]), .B2(n4744), .ZN(n4615) );
  AOI22D1BWP30P140LVT U4987 ( .A1(i_data_bus[825]), .A2(n4076), .B1(
        i_data_bus[889]), .B2(n4743), .ZN(n4614) );
  AOI22D1BWP30P140LVT U4988 ( .A1(i_data_bus[569]), .A2(n4723), .B1(
        i_data_bus[121]), .B2(n4750), .ZN(n4613) );
  ND4D1BWP30P140LVT U4989 ( .A1(n4616), .A2(n4615), .A3(n4614), .A4(n4613), 
        .ZN(n4617) );
  OR4D1BWP30P140LVT U4990 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), 
        .Z(o_data_bus[217]) );
  AOI22D1BWP30P140LVT U4991 ( .A1(i_data_bus[954]), .A2(n4070), .B1(
        i_data_bus[986]), .B2(n4068), .ZN(n4624) );
  AOI22D1BWP30P140LVT U4992 ( .A1(i_data_bus[1018]), .A2(n4066), .B1(
        i_data_bus[922]), .B2(n4073), .ZN(n4623) );
  AOI22D1BWP30P140LVT U4993 ( .A1(i_data_bus[538]), .A2(n4722), .B1(
        i_data_bus[666]), .B2(n4730), .ZN(n4622) );
  AOI22D1BWP30P140LVT U4994 ( .A1(i_data_bus[698]), .A2(n4075), .B1(
        i_data_bus[378]), .B2(n4739), .ZN(n4621) );
  ND4D1BWP30P140LVT U4995 ( .A1(n4624), .A2(n4623), .A3(n4622), .A4(n4621), 
        .ZN(n4640) );
  AOI22D1BWP30P140LVT U4996 ( .A1(i_data_bus[602]), .A2(n4742), .B1(
        i_data_bus[730]), .B2(n4753), .ZN(n4628) );
  AOI22D1BWP30P140LVT U4997 ( .A1(i_data_bus[570]), .A2(n4723), .B1(
        i_data_bus[506]), .B2(n4111), .ZN(n4627) );
  AOI22D1BWP30P140LVT U4998 ( .A1(i_data_bus[218]), .A2(n4744), .B1(
        i_data_bus[346]), .B2(n4729), .ZN(n4626) );
  AOI22D1BWP30P140LVT U4999 ( .A1(i_data_bus[442]), .A2(n4732), .B1(
        i_data_bus[762]), .B2(n4088), .ZN(n4625) );
  ND4D1BWP30P140LVT U5000 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), 
        .ZN(n4639) );
  AOI22D1BWP30P140LVT U5001 ( .A1(i_data_bus[634]), .A2(n4733), .B1(
        i_data_bus[282]), .B2(n4731), .ZN(n4632) );
  AOI22D1BWP30P140LVT U5002 ( .A1(i_data_bus[58]), .A2(n4740), .B1(
        i_data_bus[314]), .B2(n4741), .ZN(n4631) );
  AOI22D1BWP30P140LVT U5003 ( .A1(i_data_bus[26]), .A2(n4097), .B1(
        i_data_bus[794]), .B2(n4721), .ZN(n4630) );
  AOI22D1BWP30P140LVT U5004 ( .A1(i_data_bus[826]), .A2(n4076), .B1(
        i_data_bus[474]), .B2(n4751), .ZN(n4629) );
  ND4D1BWP30P140LVT U5005 ( .A1(n4632), .A2(n4631), .A3(n4630), .A4(n4629), 
        .ZN(n4638) );
  AOI22D1BWP30P140LVT U5006 ( .A1(i_data_bus[858]), .A2(n4096), .B1(
        i_data_bus[250]), .B2(n4749), .ZN(n4636) );
  AOI22D1BWP30P140LVT U5007 ( .A1(i_data_bus[90]), .A2(n4724), .B1(
        i_data_bus[186]), .B2(n4738), .ZN(n4635) );
  AOI22D1BWP30P140LVT U5008 ( .A1(i_data_bus[890]), .A2(n4743), .B1(
        i_data_bus[154]), .B2(n4108), .ZN(n4634) );
  AOI22D1BWP30P140LVT U5009 ( .A1(i_data_bus[122]), .A2(n4750), .B1(
        i_data_bus[410]), .B2(n4752), .ZN(n4633) );
  ND4D1BWP30P140LVT U5010 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), 
        .ZN(n4637) );
  OR4D1BWP30P140LVT U5011 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), 
        .Z(o_data_bus[218]) );
  AOI22D1BWP30P140LVT U5012 ( .A1(i_data_bus[987]), .A2(n4068), .B1(
        i_data_bus[923]), .B2(n4073), .ZN(n4644) );
  AOI22D1BWP30P140LVT U5013 ( .A1(i_data_bus[1019]), .A2(n4066), .B1(
        i_data_bus[955]), .B2(n4070), .ZN(n4643) );
  AOI22D1BWP30P140LVT U5014 ( .A1(i_data_bus[91]), .A2(n4724), .B1(
        i_data_bus[891]), .B2(n4743), .ZN(n4642) );
  AOI22D1BWP30P140LVT U5015 ( .A1(i_data_bus[539]), .A2(n4722), .B1(
        i_data_bus[27]), .B2(n4097), .ZN(n4641) );
  ND4D1BWP30P140LVT U5016 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), 
        .ZN(n4660) );
  AOI22D1BWP30P140LVT U5017 ( .A1(i_data_bus[123]), .A2(n4750), .B1(
        i_data_bus[251]), .B2(n4749), .ZN(n4648) );
  AOI22D1BWP30P140LVT U5018 ( .A1(i_data_bus[603]), .A2(n4742), .B1(
        i_data_bus[219]), .B2(n4744), .ZN(n4647) );
  AOI22D1BWP30P140LVT U5019 ( .A1(i_data_bus[763]), .A2(n4088), .B1(
        i_data_bus[187]), .B2(n4738), .ZN(n4646) );
  AOI22D1BWP30P140LVT U5020 ( .A1(i_data_bus[571]), .A2(n4723), .B1(
        i_data_bus[635]), .B2(n4733), .ZN(n4645) );
  ND4D1BWP30P140LVT U5021 ( .A1(n4648), .A2(n4647), .A3(n4646), .A4(n4645), 
        .ZN(n4659) );
  AOI22D1BWP30P140LVT U5022 ( .A1(i_data_bus[443]), .A2(n4732), .B1(
        i_data_bus[315]), .B2(n4741), .ZN(n4652) );
  AOI22D1BWP30P140LVT U5023 ( .A1(i_data_bus[59]), .A2(n4740), .B1(
        i_data_bus[379]), .B2(n4739), .ZN(n4651) );
  AOI22D1BWP30P140LVT U5024 ( .A1(i_data_bus[411]), .A2(n4752), .B1(
        i_data_bus[795]), .B2(n4721), .ZN(n4650) );
  AOI22D1BWP30P140LVT U5025 ( .A1(i_data_bus[155]), .A2(n4108), .B1(
        i_data_bus[667]), .B2(n4730), .ZN(n4649) );
  ND4D1BWP30P140LVT U5026 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), 
        .ZN(n4658) );
  AOI22D1BWP30P140LVT U5027 ( .A1(i_data_bus[731]), .A2(n4753), .B1(
        i_data_bus[859]), .B2(n4096), .ZN(n4656) );
  AOI22D1BWP30P140LVT U5028 ( .A1(i_data_bus[283]), .A2(n4731), .B1(
        i_data_bus[475]), .B2(n4751), .ZN(n4655) );
  AOI22D1BWP30P140LVT U5029 ( .A1(i_data_bus[827]), .A2(n4076), .B1(
        i_data_bus[699]), .B2(n4075), .ZN(n4654) );
  AOI22D1BWP30P140LVT U5030 ( .A1(i_data_bus[507]), .A2(n4111), .B1(
        i_data_bus[347]), .B2(n4729), .ZN(n4653) );
  ND4D1BWP30P140LVT U5031 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), 
        .ZN(n4657) );
  OR4D1BWP30P140LVT U5032 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), 
        .Z(o_data_bus[219]) );
  AOI22D1BWP30P140LVT U5033 ( .A1(i_data_bus[988]), .A2(n4068), .B1(
        i_data_bus[956]), .B2(n4070), .ZN(n4664) );
  AOI22D1BWP30P140LVT U5034 ( .A1(i_data_bus[924]), .A2(n4073), .B1(
        i_data_bus[1020]), .B2(n4066), .ZN(n4663) );
  AOI22D1BWP30P140LVT U5035 ( .A1(i_data_bus[764]), .A2(n4088), .B1(
        i_data_bus[316]), .B2(n4741), .ZN(n4662) );
  AOI22D1BWP30P140LVT U5036 ( .A1(i_data_bus[188]), .A2(n4738), .B1(
        i_data_bus[860]), .B2(n4096), .ZN(n4661) );
  ND4D1BWP30P140LVT U5037 ( .A1(n4664), .A2(n4663), .A3(n4662), .A4(n4661), 
        .ZN(n4680) );
  AOI22D1BWP30P140LVT U5038 ( .A1(i_data_bus[348]), .A2(n4729), .B1(
        i_data_bus[796]), .B2(n4721), .ZN(n4668) );
  AOI22D1BWP30P140LVT U5039 ( .A1(i_data_bus[28]), .A2(n4097), .B1(
        i_data_bus[444]), .B2(n4732), .ZN(n4667) );
  AOI22D1BWP30P140LVT U5040 ( .A1(i_data_bus[636]), .A2(n4733), .B1(
        i_data_bus[572]), .B2(n4723), .ZN(n4666) );
  AOI22D1BWP30P140LVT U5041 ( .A1(i_data_bus[604]), .A2(n4742), .B1(
        i_data_bus[380]), .B2(n4739), .ZN(n4665) );
  ND4D1BWP30P140LVT U5042 ( .A1(n4668), .A2(n4667), .A3(n4666), .A4(n4665), 
        .ZN(n4679) );
  AOI22D1BWP30P140LVT U5043 ( .A1(i_data_bus[732]), .A2(n4753), .B1(
        i_data_bus[412]), .B2(n4752), .ZN(n4672) );
  AOI22D1BWP30P140LVT U5044 ( .A1(i_data_bus[124]), .A2(n4750), .B1(
        i_data_bus[284]), .B2(n4731), .ZN(n4671) );
  AOI22D1BWP30P140LVT U5045 ( .A1(i_data_bus[252]), .A2(n4749), .B1(
        i_data_bus[700]), .B2(n4075), .ZN(n4670) );
  AOI22D1BWP30P140LVT U5046 ( .A1(i_data_bus[60]), .A2(n4740), .B1(
        i_data_bus[892]), .B2(n4743), .ZN(n4669) );
  ND4D1BWP30P140LVT U5047 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), 
        .ZN(n4678) );
  AOI22D1BWP30P140LVT U5048 ( .A1(i_data_bus[828]), .A2(n4076), .B1(
        i_data_bus[156]), .B2(n4108), .ZN(n4676) );
  AOI22D1BWP30P140LVT U5049 ( .A1(i_data_bus[540]), .A2(n4722), .B1(
        i_data_bus[92]), .B2(n4724), .ZN(n4675) );
  AOI22D1BWP30P140LVT U5050 ( .A1(i_data_bus[220]), .A2(n4744), .B1(
        i_data_bus[476]), .B2(n4751), .ZN(n4674) );
  AOI22D1BWP30P140LVT U5051 ( .A1(i_data_bus[508]), .A2(n4111), .B1(
        i_data_bus[668]), .B2(n4730), .ZN(n4673) );
  ND4D1BWP30P140LVT U5052 ( .A1(n4676), .A2(n4675), .A3(n4674), .A4(n4673), 
        .ZN(n4677) );
  OR4D1BWP30P140LVT U5053 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), 
        .Z(o_data_bus[220]) );
  AOI22D1BWP30P140LVT U5054 ( .A1(i_data_bus[957]), .A2(n4070), .B1(
        i_data_bus[989]), .B2(n4068), .ZN(n4684) );
  AOI22D1BWP30P140LVT U5055 ( .A1(i_data_bus[925]), .A2(n4073), .B1(
        i_data_bus[1021]), .B2(n4066), .ZN(n4683) );
  AOI22D1BWP30P140LVT U5056 ( .A1(i_data_bus[93]), .A2(n4724), .B1(
        i_data_bus[893]), .B2(n4743), .ZN(n4682) );
  AOI22D1BWP30P140LVT U5057 ( .A1(i_data_bus[797]), .A2(n4721), .B1(
        i_data_bus[381]), .B2(n4739), .ZN(n4681) );
  ND4D1BWP30P140LVT U5058 ( .A1(n4684), .A2(n4683), .A3(n4682), .A4(n4681), 
        .ZN(n4700) );
  AOI22D1BWP30P140LVT U5059 ( .A1(i_data_bus[445]), .A2(n4732), .B1(
        i_data_bus[189]), .B2(n4738), .ZN(n4688) );
  AOI22D1BWP30P140LVT U5060 ( .A1(i_data_bus[637]), .A2(n4733), .B1(
        i_data_bus[669]), .B2(n4730), .ZN(n4687) );
  AOI22D1BWP30P140LVT U5061 ( .A1(i_data_bus[701]), .A2(n4075), .B1(
        i_data_bus[509]), .B2(n4111), .ZN(n4686) );
  AOI22D1BWP30P140LVT U5062 ( .A1(i_data_bus[573]), .A2(n4723), .B1(
        i_data_bus[829]), .B2(n4076), .ZN(n4685) );
  ND4D1BWP30P140LVT U5063 ( .A1(n4688), .A2(n4687), .A3(n4686), .A4(n4685), 
        .ZN(n4699) );
  AOI22D1BWP30P140LVT U5064 ( .A1(i_data_bus[157]), .A2(n4108), .B1(
        i_data_bus[349]), .B2(n4729), .ZN(n4692) );
  AOI22D1BWP30P140LVT U5065 ( .A1(i_data_bus[61]), .A2(n4740), .B1(
        i_data_bus[317]), .B2(n4741), .ZN(n4691) );
  AOI22D1BWP30P140LVT U5066 ( .A1(i_data_bus[765]), .A2(n4088), .B1(
        i_data_bus[733]), .B2(n4753), .ZN(n4690) );
  AOI22D1BWP30P140LVT U5067 ( .A1(i_data_bus[29]), .A2(n4097), .B1(
        i_data_bus[477]), .B2(n4751), .ZN(n4689) );
  ND4D1BWP30P140LVT U5068 ( .A1(n4692), .A2(n4691), .A3(n4690), .A4(n4689), 
        .ZN(n4698) );
  AOI22D1BWP30P140LVT U5069 ( .A1(i_data_bus[413]), .A2(n4752), .B1(
        i_data_bus[253]), .B2(n4749), .ZN(n4696) );
  AOI22D1BWP30P140LVT U5070 ( .A1(i_data_bus[605]), .A2(n4742), .B1(
        i_data_bus[221]), .B2(n4744), .ZN(n4695) );
  AOI22D1BWP30P140LVT U5071 ( .A1(i_data_bus[541]), .A2(n4722), .B1(
        i_data_bus[285]), .B2(n4731), .ZN(n4694) );
  AOI22D1BWP30P140LVT U5072 ( .A1(i_data_bus[125]), .A2(n4750), .B1(
        i_data_bus[861]), .B2(n4096), .ZN(n4693) );
  ND4D1BWP30P140LVT U5073 ( .A1(n4696), .A2(n4695), .A3(n4694), .A4(n4693), 
        .ZN(n4697) );
  OR4D1BWP30P140LVT U5074 ( .A1(n4700), .A2(n4699), .A3(n4698), .A4(n4697), 
        .Z(o_data_bus[221]) );
  AOI22D1BWP30P140LVT U5075 ( .A1(i_data_bus[958]), .A2(n4070), .B1(
        i_data_bus[990]), .B2(n4068), .ZN(n4704) );
  AOI22D1BWP30P140LVT U5076 ( .A1(i_data_bus[926]), .A2(n4073), .B1(
        i_data_bus[1022]), .B2(n4066), .ZN(n4703) );
  AOI22D1BWP30P140LVT U5077 ( .A1(i_data_bus[574]), .A2(n4723), .B1(
        i_data_bus[222]), .B2(n4744), .ZN(n4702) );
  AOI22D1BWP30P140LVT U5078 ( .A1(i_data_bus[542]), .A2(n4722), .B1(
        i_data_bus[318]), .B2(n4741), .ZN(n4701) );
  ND4D1BWP30P140LVT U5079 ( .A1(n4704), .A2(n4703), .A3(n4702), .A4(n4701), 
        .ZN(n4720) );
  AOI22D1BWP30P140LVT U5080 ( .A1(i_data_bus[62]), .A2(n4740), .B1(
        i_data_bus[350]), .B2(n4729), .ZN(n4708) );
  AOI22D1BWP30P140LVT U5081 ( .A1(i_data_bus[446]), .A2(n4732), .B1(
        i_data_bus[510]), .B2(n4111), .ZN(n4707) );
  AOI22D1BWP30P140LVT U5082 ( .A1(i_data_bus[830]), .A2(n4076), .B1(
        i_data_bus[414]), .B2(n4752), .ZN(n4706) );
  AOI22D1BWP30P140LVT U5083 ( .A1(i_data_bus[286]), .A2(n4731), .B1(
        i_data_bus[702]), .B2(n4075), .ZN(n4705) );
  ND4D1BWP30P140LVT U5084 ( .A1(n4708), .A2(n4707), .A3(n4706), .A4(n4705), 
        .ZN(n4719) );
  AOI22D1BWP30P140LVT U5085 ( .A1(i_data_bus[126]), .A2(n4750), .B1(
        i_data_bus[158]), .B2(n4108), .ZN(n4712) );
  AOI22D1BWP30P140LVT U5086 ( .A1(i_data_bus[254]), .A2(n4749), .B1(
        i_data_bus[478]), .B2(n4751), .ZN(n4711) );
  AOI22D1BWP30P140LVT U5087 ( .A1(i_data_bus[670]), .A2(n4730), .B1(
        i_data_bus[734]), .B2(n4753), .ZN(n4710) );
  AOI22D1BWP30P140LVT U5088 ( .A1(i_data_bus[94]), .A2(n4724), .B1(
        i_data_bus[862]), .B2(n4096), .ZN(n4709) );
  ND4D1BWP30P140LVT U5089 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), 
        .ZN(n4718) );
  AOI22D1BWP30P140LVT U5090 ( .A1(i_data_bus[798]), .A2(n4721), .B1(
        i_data_bus[382]), .B2(n4739), .ZN(n4716) );
  AOI22D1BWP30P140LVT U5091 ( .A1(i_data_bus[190]), .A2(n4738), .B1(
        i_data_bus[766]), .B2(n4088), .ZN(n4715) );
  AOI22D1BWP30P140LVT U5092 ( .A1(i_data_bus[30]), .A2(n4097), .B1(
        i_data_bus[606]), .B2(n4742), .ZN(n4714) );
  AOI22D1BWP30P140LVT U5093 ( .A1(i_data_bus[638]), .A2(n4733), .B1(
        i_data_bus[894]), .B2(n4743), .ZN(n4713) );
  ND4D1BWP30P140LVT U5094 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), 
        .ZN(n4717) );
  OR4D1BWP30P140LVT U5095 ( .A1(n4720), .A2(n4719), .A3(n4718), .A4(n4717), 
        .Z(o_data_bus[222]) );
  AOI22D1BWP30P140LVT U5096 ( .A1(i_data_bus[991]), .A2(n4068), .B1(
        i_data_bus[927]), .B2(n4073), .ZN(n4728) );
  AOI22D1BWP30P140LVT U5097 ( .A1(i_data_bus[1023]), .A2(n4066), .B1(
        i_data_bus[959]), .B2(n4070), .ZN(n4727) );
  AOI22D1BWP30P140LVT U5098 ( .A1(i_data_bus[543]), .A2(n4722), .B1(
        i_data_bus[799]), .B2(n4721), .ZN(n4726) );
  AOI22D1BWP30P140LVT U5099 ( .A1(i_data_bus[95]), .A2(n4724), .B1(
        i_data_bus[575]), .B2(n4723), .ZN(n4725) );
  ND4D1BWP30P140LVT U5100 ( .A1(n4728), .A2(n4727), .A3(n4726), .A4(n4725), 
        .ZN(n4761) );
  AOI22D1BWP30P140LVT U5101 ( .A1(i_data_bus[671]), .A2(n4730), .B1(
        i_data_bus[351]), .B2(n4729), .ZN(n4737) );
  AOI22D1BWP30P140LVT U5102 ( .A1(i_data_bus[31]), .A2(n4097), .B1(
        i_data_bus[159]), .B2(n4108), .ZN(n4736) );
  AOI22D1BWP30P140LVT U5103 ( .A1(i_data_bus[447]), .A2(n4732), .B1(
        i_data_bus[287]), .B2(n4731), .ZN(n4735) );
  AOI22D1BWP30P140LVT U5104 ( .A1(i_data_bus[639]), .A2(n4733), .B1(
        i_data_bus[831]), .B2(n4076), .ZN(n4734) );
  ND4D1BWP30P140LVT U5105 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), 
        .ZN(n4760) );
  AOI22D1BWP30P140LVT U5106 ( .A1(i_data_bus[703]), .A2(n4075), .B1(
        i_data_bus[191]), .B2(n4738), .ZN(n4748) );
  AOI22D1BWP30P140LVT U5107 ( .A1(i_data_bus[63]), .A2(n4740), .B1(
        i_data_bus[383]), .B2(n4739), .ZN(n4747) );
  AOI22D1BWP30P140LVT U5108 ( .A1(i_data_bus[607]), .A2(n4742), .B1(
        i_data_bus[319]), .B2(n4741), .ZN(n4746) );
  AOI22D1BWP30P140LVT U5109 ( .A1(i_data_bus[223]), .A2(n4744), .B1(
        i_data_bus[895]), .B2(n4743), .ZN(n4745) );
  ND4D1BWP30P140LVT U5110 ( .A1(n4748), .A2(n4747), .A3(n4746), .A4(n4745), 
        .ZN(n4759) );
  AOI22D1BWP30P140LVT U5111 ( .A1(i_data_bus[511]), .A2(n4111), .B1(
        i_data_bus[767]), .B2(n4088), .ZN(n4757) );
  AOI22D1BWP30P140LVT U5112 ( .A1(i_data_bus[127]), .A2(n4750), .B1(
        i_data_bus[255]), .B2(n4749), .ZN(n4756) );
  AOI22D1BWP30P140LVT U5113 ( .A1(i_data_bus[863]), .A2(n4096), .B1(
        i_data_bus[479]), .B2(n4751), .ZN(n4755) );
  AOI22D1BWP30P140LVT U5114 ( .A1(i_data_bus[735]), .A2(n4753), .B1(
        i_data_bus[415]), .B2(n4752), .ZN(n4754) );
  ND4D1BWP30P140LVT U5115 ( .A1(n4757), .A2(n4756), .A3(n4755), .A4(n4754), 
        .ZN(n4758) );
  OR4D1BWP30P140LVT U5116 ( .A1(n4761), .A2(n4760), .A3(n4759), .A4(n4758), 
        .Z(o_data_bus[223]) );
  AOI22D1BWP30P140LVT U5117 ( .A1(i_data_bus[992]), .A2(n5396), .B1(
        i_data_bus[32]), .B2(n5395), .ZN(n4782) );
  AOI22D1BWP30P140LVT U5118 ( .A1(i_data_bus[160]), .A2(n5391), .B1(
        i_data_bus[128]), .B2(n5399), .ZN(n4781) );
  AOI22D1BWP30P140LVT U5119 ( .A1(i_data_bus[480]), .A2(n223), .B1(
        i_data_bus[448]), .B2(n222), .ZN(n4780) );
  AOI22D1BWP30P140LVT U5120 ( .A1(i_data_bus[960]), .A2(n5392), .B1(
        i_data_bus[192]), .B2(n5400), .ZN(n4765) );
  AOI22D1BWP30P140LVT U5121 ( .A1(i_data_bus[96]), .A2(n5402), .B1(
        i_data_bus[224]), .B2(n5401), .ZN(n4764) );
  AOI22D1BWP30P140LVT U5122 ( .A1(i_data_bus[64]), .A2(n5390), .B1(
        i_data_bus[896]), .B2(n5389), .ZN(n4763) );
  AOI22D1BWP30P140LVT U5123 ( .A1(i_data_bus[928]), .A2(n5397), .B1(
        i_data_bus[0]), .B2(n5398), .ZN(n4762) );
  ND4D1BWP30P140LVT U5124 ( .A1(n4765), .A2(n4764), .A3(n4763), .A4(n4762), 
        .ZN(n4778) );
  MOAI22D1BWP30P140LVT U5125 ( .A1(n4766), .A2(n5351), .B1(i_data_bus[640]), 
        .B2(n5426), .ZN(n4777) );
  AOI22D1BWP30P140LVT U5126 ( .A1(i_data_bus[800]), .A2(n5427), .B1(
        i_data_bus[320]), .B2(n5422), .ZN(n4770) );
  AOI22D1BWP30P140LVT U5127 ( .A1(i_data_bus[384]), .A2(n5411), .B1(
        i_data_bus[768]), .B2(n5407), .ZN(n4769) );
  AOI22D1BWP30P140LVT U5128 ( .A1(i_data_bus[512]), .A2(n5414), .B1(
        i_data_bus[608]), .B2(n5416), .ZN(n4768) );
  AOI22D1BWP30P140LVT U5129 ( .A1(i_data_bus[544]), .A2(n5417), .B1(
        i_data_bus[576]), .B2(n5415), .ZN(n4767) );
  ND4D1BWP30P140LVT U5130 ( .A1(n4770), .A2(n4769), .A3(n4768), .A4(n4767), 
        .ZN(n4776) );
  AOI22D1BWP30P140LVT U5131 ( .A1(i_data_bus[352]), .A2(n5423), .B1(
        i_data_bus[672]), .B2(n5393), .ZN(n4774) );
  AOI22D1BWP30P140LVT U5132 ( .A1(i_data_bus[704]), .A2(n5424), .B1(
        i_data_bus[864]), .B2(n5410), .ZN(n4773) );
  AOI22D1BWP30P140LVT U5133 ( .A1(i_data_bus[416]), .A2(n5413), .B1(
        i_data_bus[288]), .B2(n5428), .ZN(n4772) );
  AOI22D1BWP30P140LVT U5134 ( .A1(i_data_bus[832]), .A2(n5425), .B1(
        i_data_bus[736]), .B2(n5412), .ZN(n4771) );
  ND4D1BWP30P140LVT U5135 ( .A1(n4774), .A2(n4773), .A3(n4772), .A4(n4771), 
        .ZN(n4775) );
  NR4D0BWP30P140LVT U5136 ( .A1(n4778), .A2(n4777), .A3(n4776), .A4(n4775), 
        .ZN(n4779) );
  ND4D1BWP30P140LVT U5137 ( .A1(n4782), .A2(n4781), .A3(n4780), .A4(n4779), 
        .ZN(o_data_bus[0]) );
  AOI22D1BWP30P140LVT U5138 ( .A1(i_data_bus[97]), .A2(n5402), .B1(
        i_data_bus[225]), .B2(n5401), .ZN(n4803) );
  AOI22D1BWP30P140LVT U5139 ( .A1(i_data_bus[65]), .A2(n5390), .B1(
        i_data_bus[193]), .B2(n5400), .ZN(n4802) );
  AOI22D1BWP30P140LVT U5140 ( .A1(i_data_bus[769]), .A2(n5407), .B1(
        i_data_bus[801]), .B2(n5427), .ZN(n4801) );
  AOI22D1BWP30P140LVT U5141 ( .A1(i_data_bus[961]), .A2(n5392), .B1(
        i_data_bus[993]), .B2(n5396), .ZN(n4786) );
  AOI22D1BWP30P140LVT U5142 ( .A1(i_data_bus[33]), .A2(n5395), .B1(
        i_data_bus[1]), .B2(n5398), .ZN(n4785) );
  AOI22D1BWP30P140LVT U5143 ( .A1(i_data_bus[897]), .A2(n5389), .B1(
        i_data_bus[929]), .B2(n5397), .ZN(n4784) );
  AOI22D1BWP30P140LVT U5144 ( .A1(i_data_bus[161]), .A2(n5391), .B1(
        i_data_bus[129]), .B2(n5399), .ZN(n4783) );
  ND4D1BWP30P140LVT U5145 ( .A1(n4786), .A2(n4785), .A3(n4784), .A4(n4783), 
        .ZN(n4799) );
  MOAI22D1BWP30P140LVT U5146 ( .A1(n4787), .A2(n5351), .B1(i_data_bus[865]), 
        .B2(n5410), .ZN(n4798) );
  AOI22D1BWP30P140LVT U5147 ( .A1(i_data_bus[705]), .A2(n5424), .B1(
        i_data_bus[321]), .B2(n5422), .ZN(n4791) );
  AOI22D1BWP30P140LVT U5148 ( .A1(i_data_bus[353]), .A2(n5423), .B1(
        i_data_bus[833]), .B2(n5425), .ZN(n4790) );
  AOI22D1BWP30P140LVT U5149 ( .A1(i_data_bus[577]), .A2(n5415), .B1(
        i_data_bus[545]), .B2(n5417), .ZN(n4789) );
  AOI22D1BWP30P140LVT U5150 ( .A1(i_data_bus[609]), .A2(n5416), .B1(
        i_data_bus[513]), .B2(n5414), .ZN(n4788) );
  ND4D1BWP30P140LVT U5151 ( .A1(n4791), .A2(n4790), .A3(n4789), .A4(n4788), 
        .ZN(n4797) );
  AOI22D1BWP30P140LVT U5152 ( .A1(i_data_bus[673]), .A2(n5393), .B1(
        i_data_bus[417]), .B2(n5413), .ZN(n4795) );
  AOI22D1BWP30P140LVT U5153 ( .A1(i_data_bus[449]), .A2(n222), .B1(
        i_data_bus[289]), .B2(n5428), .ZN(n4794) );
  AOI22D1BWP30P140LVT U5154 ( .A1(i_data_bus[481]), .A2(n223), .B1(
        i_data_bus[737]), .B2(n5412), .ZN(n4793) );
  AOI22D1BWP30P140LVT U5155 ( .A1(i_data_bus[385]), .A2(n5411), .B1(
        i_data_bus[641]), .B2(n5426), .ZN(n4792) );
  ND4D1BWP30P140LVT U5156 ( .A1(n4795), .A2(n4794), .A3(n4793), .A4(n4792), 
        .ZN(n4796) );
  NR4D0BWP30P140LVT U5157 ( .A1(n4799), .A2(n4798), .A3(n4797), .A4(n4796), 
        .ZN(n4800) );
  ND4D1BWP30P140LVT U5158 ( .A1(n4803), .A2(n4802), .A3(n4801), .A4(n4800), 
        .ZN(o_data_bus[1]) );
  AOI22D1BWP30P140LVT U5159 ( .A1(i_data_bus[962]), .A2(n5392), .B1(
        i_data_bus[994]), .B2(n5396), .ZN(n4824) );
  AOI22D1BWP30P140LVT U5160 ( .A1(i_data_bus[2]), .A2(n5398), .B1(
        i_data_bus[930]), .B2(n5397), .ZN(n4823) );
  AOI22D1BWP30P140LVT U5161 ( .A1(i_data_bus[450]), .A2(n222), .B1(
        i_data_bus[770]), .B2(n5407), .ZN(n4822) );
  AOI22D1BWP30P140LVT U5162 ( .A1(i_data_bus[98]), .A2(n5402), .B1(
        i_data_bus[130]), .B2(n5399), .ZN(n4807) );
  AOI22D1BWP30P140LVT U5163 ( .A1(i_data_bus[66]), .A2(n5390), .B1(
        i_data_bus[898]), .B2(n5389), .ZN(n4806) );
  AOI22D1BWP30P140LVT U5164 ( .A1(i_data_bus[34]), .A2(n5395), .B1(
        i_data_bus[194]), .B2(n5400), .ZN(n4805) );
  AOI22D1BWP30P140LVT U5165 ( .A1(i_data_bus[162]), .A2(n5391), .B1(
        i_data_bus[226]), .B2(n5401), .ZN(n4804) );
  ND4D1BWP30P140LVT U5166 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), 
        .ZN(n4820) );
  OAI22D1BWP30P140LVT U5167 ( .A1(n5535), .A2(n5351), .B1(n4808), .B2(n5220), 
        .ZN(n4819) );
  AOI22D1BWP30P140LVT U5168 ( .A1(i_data_bus[802]), .A2(n5427), .B1(
        i_data_bus[738]), .B2(n5412), .ZN(n4812) );
  AOI22D1BWP30P140LVT U5169 ( .A1(i_data_bus[482]), .A2(n223), .B1(
        i_data_bus[706]), .B2(n5424), .ZN(n4811) );
  AOI22D1BWP30P140LVT U5170 ( .A1(i_data_bus[578]), .A2(n5415), .B1(
        i_data_bus[546]), .B2(n5417), .ZN(n4810) );
  AOI22D1BWP30P140LVT U5171 ( .A1(i_data_bus[514]), .A2(n5414), .B1(
        i_data_bus[610]), .B2(n5416), .ZN(n4809) );
  ND4D1BWP30P140LVT U5172 ( .A1(n4812), .A2(n4811), .A3(n4810), .A4(n4809), 
        .ZN(n4818) );
  AOI22D1BWP30P140LVT U5173 ( .A1(i_data_bus[418]), .A2(n5413), .B1(
        i_data_bus[354]), .B2(n5423), .ZN(n4816) );
  AOI22D1BWP30P140LVT U5174 ( .A1(i_data_bus[674]), .A2(n5393), .B1(
        i_data_bus[834]), .B2(n5425), .ZN(n4815) );
  AOI22D1BWP30P140LVT U5175 ( .A1(i_data_bus[866]), .A2(n5410), .B1(
        i_data_bus[386]), .B2(n5411), .ZN(n4814) );
  AOI22D1BWP30P140LVT U5176 ( .A1(i_data_bus[290]), .A2(n5428), .B1(
        i_data_bus[642]), .B2(n5426), .ZN(n4813) );
  ND4D1BWP30P140LVT U5177 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), 
        .ZN(n4817) );
  NR4D0BWP30P140LVT U5178 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), 
        .ZN(n4821) );
  ND4D1BWP30P140LVT U5179 ( .A1(n4824), .A2(n4823), .A3(n4822), .A4(n4821), 
        .ZN(o_data_bus[2]) );
  AOI22D1BWP30P140LVT U5180 ( .A1(i_data_bus[99]), .A2(n5402), .B1(
        i_data_bus[963]), .B2(n5392), .ZN(n4844) );
  AOI22D1BWP30P140LVT U5181 ( .A1(i_data_bus[899]), .A2(n5389), .B1(
        i_data_bus[35]), .B2(n5395), .ZN(n4843) );
  AOI22D1BWP30P140LVT U5182 ( .A1(i_data_bus[771]), .A2(n5407), .B1(
        i_data_bus[739]), .B2(n5412), .ZN(n4842) );
  AOI22D1BWP30P140LVT U5183 ( .A1(i_data_bus[643]), .A2(n5426), .B1(
        i_data_bus[867]), .B2(n5410), .ZN(n4840) );
  AOI22D1BWP30P140LVT U5184 ( .A1(i_data_bus[931]), .A2(n5397), .B1(
        i_data_bus[227]), .B2(n5401), .ZN(n4828) );
  AOI22D1BWP30P140LVT U5185 ( .A1(i_data_bus[995]), .A2(n5396), .B1(
        i_data_bus[163]), .B2(n5391), .ZN(n4827) );
  AOI22D1BWP30P140LVT U5186 ( .A1(i_data_bus[67]), .A2(n5390), .B1(
        i_data_bus[3]), .B2(n5398), .ZN(n4826) );
  AOI22D1BWP30P140LVT U5187 ( .A1(i_data_bus[131]), .A2(n5399), .B1(
        i_data_bus[195]), .B2(n5400), .ZN(n4825) );
  ND4D1BWP30P140LVT U5188 ( .A1(n4828), .A2(n4827), .A3(n4826), .A4(n4825), 
        .ZN(n4839) );
  AOI22D1BWP30P140LVT U5189 ( .A1(i_data_bus[835]), .A2(n5425), .B1(
        i_data_bus[323]), .B2(n5422), .ZN(n4832) );
  AOI22D1BWP30P140LVT U5190 ( .A1(i_data_bus[387]), .A2(n5411), .B1(
        i_data_bus[675]), .B2(n5393), .ZN(n4831) );
  AOI22D1BWP30P140LVT U5191 ( .A1(i_data_bus[547]), .A2(n5417), .B1(
        i_data_bus[611]), .B2(n5416), .ZN(n4830) );
  AOI22D1BWP30P140LVT U5192 ( .A1(i_data_bus[515]), .A2(n5414), .B1(
        i_data_bus[579]), .B2(n5415), .ZN(n4829) );
  ND4D1BWP30P140LVT U5193 ( .A1(n4832), .A2(n4831), .A3(n4830), .A4(n4829), 
        .ZN(n4838) );
  AOI22D1BWP30P140LVT U5194 ( .A1(i_data_bus[419]), .A2(n5413), .B1(
        i_data_bus[291]), .B2(n5428), .ZN(n4836) );
  AOI22D1BWP30P140LVT U5195 ( .A1(i_data_bus[707]), .A2(n5424), .B1(
        i_data_bus[451]), .B2(n222), .ZN(n4835) );
  AOI22D1BWP30P140LVT U5196 ( .A1(i_data_bus[355]), .A2(n5423), .B1(
        i_data_bus[259]), .B2(n5394), .ZN(n4834) );
  AOI22D1BWP30P140LVT U5197 ( .A1(i_data_bus[483]), .A2(n223), .B1(
        i_data_bus[803]), .B2(n5427), .ZN(n4833) );
  ND4D1BWP30P140LVT U5198 ( .A1(n4836), .A2(n4835), .A3(n4834), .A4(n4833), 
        .ZN(n4837) );
  INR4D0BWP30P140LVT U5199 ( .A1(n4840), .B1(n4839), .B2(n4838), .B3(n4837), 
        .ZN(n4841) );
  ND4D1BWP30P140LVT U5200 ( .A1(n4844), .A2(n4843), .A3(n4842), .A4(n4841), 
        .ZN(o_data_bus[3]) );
  AOI22D1BWP30P140LVT U5201 ( .A1(i_data_bus[932]), .A2(n5397), .B1(
        i_data_bus[132]), .B2(n5399), .ZN(n4865) );
  AOI22D1BWP30P140LVT U5202 ( .A1(i_data_bus[36]), .A2(n5395), .B1(
        i_data_bus[196]), .B2(n5400), .ZN(n4864) );
  AOI22D1BWP30P140LVT U5203 ( .A1(i_data_bus[452]), .A2(n222), .B1(
        i_data_bus[484]), .B2(n223), .ZN(n4863) );
  AOI22D1BWP30P140LVT U5204 ( .A1(i_data_bus[964]), .A2(n5392), .B1(
        i_data_bus[996]), .B2(n5396), .ZN(n4848) );
  AOI22D1BWP30P140LVT U5205 ( .A1(i_data_bus[4]), .A2(n5398), .B1(
        i_data_bus[228]), .B2(n5401), .ZN(n4847) );
  AOI22D1BWP30P140LVT U5206 ( .A1(i_data_bus[100]), .A2(n5402), .B1(
        i_data_bus[164]), .B2(n5391), .ZN(n4846) );
  AOI22D1BWP30P140LVT U5207 ( .A1(i_data_bus[900]), .A2(n5389), .B1(
        i_data_bus[68]), .B2(n5390), .ZN(n4845) );
  ND4D1BWP30P140LVT U5208 ( .A1(n4848), .A2(n4847), .A3(n4846), .A4(n4845), 
        .ZN(n4861) );
  MOAI22D1BWP30P140LVT U5209 ( .A1(n4849), .A2(n5220), .B1(i_data_bus[676]), 
        .B2(n5393), .ZN(n4860) );
  AOI22D1BWP30P140LVT U5210 ( .A1(i_data_bus[708]), .A2(n5424), .B1(
        i_data_bus[420]), .B2(n5413), .ZN(n4853) );
  AOI22D1BWP30P140LVT U5211 ( .A1(i_data_bus[740]), .A2(n5412), .B1(
        i_data_bus[772]), .B2(n5407), .ZN(n4852) );
  AOI22D1BWP30P140LVT U5212 ( .A1(i_data_bus[548]), .A2(n5417), .B1(
        i_data_bus[516]), .B2(n5414), .ZN(n4851) );
  AOI22D1BWP30P140LVT U5213 ( .A1(i_data_bus[612]), .A2(n5416), .B1(
        i_data_bus[580]), .B2(n5415), .ZN(n4850) );
  ND4D1BWP30P140LVT U5214 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), 
        .ZN(n4859) );
  AOI22D1BWP30P140LVT U5215 ( .A1(i_data_bus[868]), .A2(n5410), .B1(
        i_data_bus[292]), .B2(n5428), .ZN(n4857) );
  AOI22D1BWP30P140LVT U5216 ( .A1(i_data_bus[260]), .A2(n5394), .B1(
        i_data_bus[388]), .B2(n5411), .ZN(n4856) );
  AOI22D1BWP30P140LVT U5217 ( .A1(i_data_bus[836]), .A2(n5425), .B1(
        i_data_bus[804]), .B2(n5427), .ZN(n4855) );
  AOI22D1BWP30P140LVT U5218 ( .A1(i_data_bus[644]), .A2(n5426), .B1(
        i_data_bus[356]), .B2(n5423), .ZN(n4854) );
  ND4D1BWP30P140LVT U5219 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), 
        .ZN(n4858) );
  NR4D0BWP30P140LVT U5220 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), 
        .ZN(n4862) );
  ND4D1BWP30P140LVT U5221 ( .A1(n4865), .A2(n4864), .A3(n4863), .A4(n4862), 
        .ZN(o_data_bus[4]) );
  AOI22D1BWP30P140LVT U5222 ( .A1(i_data_bus[37]), .A2(n5395), .B1(
        i_data_bus[997]), .B2(n5396), .ZN(n4885) );
  AOI22D1BWP30P140LVT U5223 ( .A1(i_data_bus[901]), .A2(n5389), .B1(
        i_data_bus[229]), .B2(n5401), .ZN(n4884) );
  AOI22D1BWP30P140LVT U5224 ( .A1(i_data_bus[485]), .A2(n223), .B1(
        i_data_bus[261]), .B2(n5394), .ZN(n4883) );
  AOI22D1BWP30P140LVT U5225 ( .A1(i_data_bus[101]), .A2(n5402), .B1(
        i_data_bus[69]), .B2(n5390), .ZN(n4869) );
  AOI22D1BWP30P140LVT U5226 ( .A1(i_data_bus[5]), .A2(n5398), .B1(
        i_data_bus[133]), .B2(n5399), .ZN(n4868) );
  AOI22D1BWP30P140LVT U5227 ( .A1(i_data_bus[933]), .A2(n5397), .B1(
        i_data_bus[965]), .B2(n5392), .ZN(n4867) );
  AOI22D1BWP30P140LVT U5228 ( .A1(i_data_bus[197]), .A2(n5400), .B1(
        i_data_bus[165]), .B2(n5391), .ZN(n4866) );
  ND4D1BWP30P140LVT U5229 ( .A1(n4869), .A2(n4868), .A3(n4867), .A4(n4866), 
        .ZN(n4881) );
  MOAI22D1BWP30P140LVT U5230 ( .A1(n5600), .A2(n5264), .B1(i_data_bus[741]), 
        .B2(n5412), .ZN(n4880) );
  AOI22D1BWP30P140LVT U5231 ( .A1(i_data_bus[645]), .A2(n5426), .B1(
        i_data_bus[325]), .B2(n5422), .ZN(n4873) );
  AOI22D1BWP30P140LVT U5232 ( .A1(i_data_bus[773]), .A2(n5407), .B1(
        i_data_bus[421]), .B2(n5413), .ZN(n4872) );
  AOI22D1BWP30P140LVT U5233 ( .A1(i_data_bus[549]), .A2(n5417), .B1(
        i_data_bus[581]), .B2(n5415), .ZN(n4871) );
  AOI22D1BWP30P140LVT U5234 ( .A1(i_data_bus[517]), .A2(n5414), .B1(
        i_data_bus[613]), .B2(n5416), .ZN(n4870) );
  ND4D1BWP30P140LVT U5235 ( .A1(n4873), .A2(n4872), .A3(n4871), .A4(n4870), 
        .ZN(n4879) );
  AOI22D1BWP30P140LVT U5236 ( .A1(i_data_bus[453]), .A2(n222), .B1(
        i_data_bus[357]), .B2(n5423), .ZN(n4877) );
  AOI22D1BWP30P140LVT U5237 ( .A1(i_data_bus[837]), .A2(n5425), .B1(
        i_data_bus[869]), .B2(n5410), .ZN(n4876) );
  AOI22D1BWP30P140LVT U5238 ( .A1(i_data_bus[677]), .A2(n5393), .B1(
        i_data_bus[805]), .B2(n5427), .ZN(n4875) );
  AOI22D1BWP30P140LVT U5239 ( .A1(i_data_bus[709]), .A2(n5424), .B1(
        i_data_bus[389]), .B2(n5411), .ZN(n4874) );
  ND4D1BWP30P140LVT U5240 ( .A1(n4877), .A2(n4876), .A3(n4875), .A4(n4874), 
        .ZN(n4878) );
  NR4D0BWP30P140LVT U5241 ( .A1(n4881), .A2(n4880), .A3(n4879), .A4(n4878), 
        .ZN(n4882) );
  ND4D1BWP30P140LVT U5242 ( .A1(n4885), .A2(n4884), .A3(n4883), .A4(n4882), 
        .ZN(o_data_bus[5]) );
  AOI22D1BWP30P140LVT U5243 ( .A1(i_data_bus[966]), .A2(n5392), .B1(
        i_data_bus[198]), .B2(n5400), .ZN(n4906) );
  AOI22D1BWP30P140LVT U5244 ( .A1(i_data_bus[934]), .A2(n5397), .B1(
        i_data_bus[166]), .B2(n5391), .ZN(n4905) );
  AOI22D1BWP30P140LVT U5245 ( .A1(i_data_bus[774]), .A2(n5407), .B1(
        i_data_bus[294]), .B2(n5428), .ZN(n4904) );
  AOI22D1BWP30P140LVT U5246 ( .A1(i_data_bus[998]), .A2(n5396), .B1(
        i_data_bus[230]), .B2(n5401), .ZN(n4889) );
  AOI22D1BWP30P140LVT U5247 ( .A1(i_data_bus[102]), .A2(n5402), .B1(
        i_data_bus[134]), .B2(n5399), .ZN(n4888) );
  AOI22D1BWP30P140LVT U5248 ( .A1(i_data_bus[6]), .A2(n5398), .B1(
        i_data_bus[70]), .B2(n5390), .ZN(n4887) );
  AOI22D1BWP30P140LVT U5249 ( .A1(i_data_bus[38]), .A2(n5395), .B1(
        i_data_bus[902]), .B2(n5389), .ZN(n4886) );
  ND4D1BWP30P140LVT U5250 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), 
        .ZN(n4902) );
  MOAI22D1BWP30P140LVT U5251 ( .A1(n4890), .A2(n228), .B1(i_data_bus[422]), 
        .B2(n5413), .ZN(n4901) );
  AOI22D1BWP30P140LVT U5252 ( .A1(i_data_bus[646]), .A2(n5426), .B1(
        i_data_bus[454]), .B2(n222), .ZN(n4894) );
  AOI22D1BWP30P140LVT U5253 ( .A1(i_data_bus[806]), .A2(n5427), .B1(
        i_data_bus[870]), .B2(n5410), .ZN(n4893) );
  AOI22D1BWP30P140LVT U5254 ( .A1(i_data_bus[550]), .A2(n5417), .B1(
        i_data_bus[518]), .B2(n5414), .ZN(n4892) );
  AOI22D1BWP30P140LVT U5255 ( .A1(i_data_bus[582]), .A2(n5415), .B1(
        i_data_bus[614]), .B2(n5416), .ZN(n4891) );
  ND4D1BWP30P140LVT U5256 ( .A1(n4894), .A2(n4893), .A3(n4892), .A4(n4891), 
        .ZN(n4900) );
  AOI22D1BWP30P140LVT U5257 ( .A1(i_data_bus[838]), .A2(n5425), .B1(
        i_data_bus[710]), .B2(n5424), .ZN(n4898) );
  AOI22D1BWP30P140LVT U5258 ( .A1(i_data_bus[486]), .A2(n223), .B1(
        i_data_bus[678]), .B2(n5393), .ZN(n4897) );
  AOI22D1BWP30P140LVT U5259 ( .A1(i_data_bus[742]), .A2(n5412), .B1(
        i_data_bus[262]), .B2(n5394), .ZN(n4896) );
  AOI22D1BWP30P140LVT U5260 ( .A1(i_data_bus[358]), .A2(n5423), .B1(
        i_data_bus[326]), .B2(n5422), .ZN(n4895) );
  ND4D1BWP30P140LVT U5261 ( .A1(n4898), .A2(n4897), .A3(n4896), .A4(n4895), 
        .ZN(n4899) );
  NR4D0BWP30P140LVT U5262 ( .A1(n4902), .A2(n4901), .A3(n4900), .A4(n4899), 
        .ZN(n4903) );
  ND4D1BWP30P140LVT U5263 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), 
        .ZN(o_data_bus[6]) );
  AOI22D1BWP30P140LVT U5264 ( .A1(i_data_bus[71]), .A2(n5390), .B1(
        i_data_bus[231]), .B2(n5401), .ZN(n4928) );
  AOI22D1BWP30P140LVT U5265 ( .A1(i_data_bus[967]), .A2(n5392), .B1(
        i_data_bus[999]), .B2(n5396), .ZN(n4927) );
  AOI22D1BWP30P140LVT U5266 ( .A1(i_data_bus[391]), .A2(n5411), .B1(
        i_data_bus[711]), .B2(n5424), .ZN(n4926) );
  AOI22D1BWP30P140LVT U5267 ( .A1(i_data_bus[7]), .A2(n5398), .B1(
        i_data_bus[199]), .B2(n5400), .ZN(n4910) );
  AOI22D1BWP30P140LVT U5268 ( .A1(i_data_bus[39]), .A2(n5395), .B1(
        i_data_bus[135]), .B2(n5399), .ZN(n4909) );
  AOI22D1BWP30P140LVT U5269 ( .A1(i_data_bus[103]), .A2(n5402), .B1(
        i_data_bus[935]), .B2(n5397), .ZN(n4908) );
  AOI22D1BWP30P140LVT U5270 ( .A1(i_data_bus[903]), .A2(n5389), .B1(
        i_data_bus[167]), .B2(n5391), .ZN(n4907) );
  ND4D1BWP30P140LVT U5271 ( .A1(n4910), .A2(n4909), .A3(n4908), .A4(n4907), 
        .ZN(n4924) );
  MOAI22D1BWP30P140LVT U5272 ( .A1(n4912), .A2(n4911), .B1(i_data_bus[423]), 
        .B2(n5413), .ZN(n4923) );
  AOI22D1BWP30P140LVT U5273 ( .A1(i_data_bus[871]), .A2(n5410), .B1(
        i_data_bus[647]), .B2(n5426), .ZN(n4916) );
  AOI22D1BWP30P140LVT U5274 ( .A1(i_data_bus[807]), .A2(n5427), .B1(
        i_data_bus[295]), .B2(n5428), .ZN(n4915) );
  AOI22D1BWP30P140LVT U5275 ( .A1(i_data_bus[519]), .A2(n5414), .B1(
        i_data_bus[583]), .B2(n5415), .ZN(n4914) );
  AOI22D1BWP30P140LVT U5276 ( .A1(i_data_bus[615]), .A2(n5416), .B1(
        i_data_bus[551]), .B2(n5417), .ZN(n4913) );
  ND4D1BWP30P140LVT U5277 ( .A1(n4916), .A2(n4915), .A3(n4914), .A4(n4913), 
        .ZN(n4922) );
  AOI22D1BWP30P140LVT U5278 ( .A1(i_data_bus[455]), .A2(n222), .B1(
        i_data_bus[775]), .B2(n5407), .ZN(n4920) );
  AOI22D1BWP30P140LVT U5279 ( .A1(i_data_bus[263]), .A2(n5394), .B1(
        i_data_bus[743]), .B2(n5412), .ZN(n4919) );
  AOI22D1BWP30P140LVT U5280 ( .A1(i_data_bus[679]), .A2(n5393), .B1(
        i_data_bus[839]), .B2(n5425), .ZN(n4918) );
  AOI22D1BWP30P140LVT U5281 ( .A1(i_data_bus[487]), .A2(n223), .B1(
        i_data_bus[327]), .B2(n5422), .ZN(n4917) );
  ND4D1BWP30P140LVT U5282 ( .A1(n4920), .A2(n4919), .A3(n4918), .A4(n4917), 
        .ZN(n4921) );
  NR4D0BWP30P140LVT U5283 ( .A1(n4924), .A2(n4923), .A3(n4922), .A4(n4921), 
        .ZN(n4925) );
  ND4D1BWP30P140LVT U5284 ( .A1(n4928), .A2(n4927), .A3(n4926), .A4(n4925), 
        .ZN(o_data_bus[7]) );
  AOI22D1BWP30P140LVT U5285 ( .A1(i_data_bus[904]), .A2(n5389), .B1(
        i_data_bus[232]), .B2(n5401), .ZN(n4948) );
  AOI22D1BWP30P140LVT U5286 ( .A1(i_data_bus[936]), .A2(n5397), .B1(
        i_data_bus[40]), .B2(n5395), .ZN(n4947) );
  AOI22D1BWP30P140LVT U5287 ( .A1(i_data_bus[680]), .A2(n5393), .B1(
        i_data_bus[488]), .B2(n223), .ZN(n4946) );
  AOI22D1BWP30P140LVT U5288 ( .A1(i_data_bus[72]), .A2(n5390), .B1(
        i_data_bus[200]), .B2(n5400), .ZN(n4932) );
  AOI22D1BWP30P140LVT U5289 ( .A1(i_data_bus[168]), .A2(n5391), .B1(
        i_data_bus[136]), .B2(n5399), .ZN(n4931) );
  AOI22D1BWP30P140LVT U5290 ( .A1(i_data_bus[8]), .A2(n5398), .B1(
        i_data_bus[1000]), .B2(n5396), .ZN(n4930) );
  AOI22D1BWP30P140LVT U5291 ( .A1(i_data_bus[968]), .A2(n5392), .B1(
        i_data_bus[104]), .B2(n5402), .ZN(n4929) );
  ND4D1BWP30P140LVT U5292 ( .A1(n4932), .A2(n4931), .A3(n4930), .A4(n4929), 
        .ZN(n4944) );
  MOAI22D1BWP30P140LVT U5293 ( .A1(n5663), .A2(n5264), .B1(i_data_bus[712]), 
        .B2(n5424), .ZN(n4943) );
  AOI22D1BWP30P140LVT U5294 ( .A1(i_data_bus[456]), .A2(n222), .B1(
        i_data_bus[360]), .B2(n5423), .ZN(n4936) );
  AOI22D1BWP30P140LVT U5295 ( .A1(i_data_bus[424]), .A2(n5413), .B1(
        i_data_bus[648]), .B2(n5426), .ZN(n4935) );
  AOI22D1BWP30P140LVT U5296 ( .A1(i_data_bus[552]), .A2(n5417), .B1(
        i_data_bus[520]), .B2(n5414), .ZN(n4934) );
  AOI22D1BWP30P140LVT U5297 ( .A1(i_data_bus[616]), .A2(n5416), .B1(
        i_data_bus[584]), .B2(n5415), .ZN(n4933) );
  ND4D1BWP30P140LVT U5298 ( .A1(n4936), .A2(n4935), .A3(n4934), .A4(n4933), 
        .ZN(n4942) );
  AOI22D1BWP30P140LVT U5299 ( .A1(i_data_bus[328]), .A2(n5422), .B1(
        i_data_bus[776]), .B2(n5407), .ZN(n4940) );
  AOI22D1BWP30P140LVT U5300 ( .A1(i_data_bus[264]), .A2(n5394), .B1(
        i_data_bus[808]), .B2(n5427), .ZN(n4939) );
  AOI22D1BWP30P140LVT U5301 ( .A1(i_data_bus[840]), .A2(n5425), .B1(
        i_data_bus[872]), .B2(n5410), .ZN(n4938) );
  AOI22D1BWP30P140LVT U5302 ( .A1(i_data_bus[744]), .A2(n5412), .B1(
        i_data_bus[392]), .B2(n5411), .ZN(n4937) );
  ND4D1BWP30P140LVT U5303 ( .A1(n4940), .A2(n4939), .A3(n4938), .A4(n4937), 
        .ZN(n4941) );
  NR4D0BWP30P140LVT U5304 ( .A1(n4944), .A2(n4943), .A3(n4942), .A4(n4941), 
        .ZN(n4945) );
  ND4D1BWP30P140LVT U5305 ( .A1(n4948), .A2(n4947), .A3(n4946), .A4(n4945), 
        .ZN(o_data_bus[8]) );
  AOI22D1BWP30P140LVT U5306 ( .A1(i_data_bus[41]), .A2(n5395), .B1(
        i_data_bus[937]), .B2(n5397), .ZN(n4969) );
  AOI22D1BWP30P140LVT U5307 ( .A1(i_data_bus[73]), .A2(n5390), .B1(
        i_data_bus[233]), .B2(n5401), .ZN(n4968) );
  AOI22D1BWP30P140LVT U5308 ( .A1(i_data_bus[809]), .A2(n5427), .B1(
        i_data_bus[777]), .B2(n5407), .ZN(n4967) );
  AOI22D1BWP30P140LVT U5309 ( .A1(i_data_bus[9]), .A2(n5398), .B1(
        i_data_bus[169]), .B2(n5391), .ZN(n4952) );
  AOI22D1BWP30P140LVT U5310 ( .A1(i_data_bus[969]), .A2(n5392), .B1(
        i_data_bus[1001]), .B2(n5396), .ZN(n4951) );
  AOI22D1BWP30P140LVT U5311 ( .A1(i_data_bus[105]), .A2(n5402), .B1(
        i_data_bus[201]), .B2(n5400), .ZN(n4950) );
  AOI22D1BWP30P140LVT U5312 ( .A1(i_data_bus[905]), .A2(n5389), .B1(
        i_data_bus[137]), .B2(n5399), .ZN(n4949) );
  ND4D1BWP30P140LVT U5313 ( .A1(n4952), .A2(n4951), .A3(n4950), .A4(n4949), 
        .ZN(n4965) );
  OAI22D1BWP30P140LVT U5314 ( .A1(n4953), .A2(n5308), .B1(n5684), .B2(n5264), 
        .ZN(n4964) );
  AOI22D1BWP30P140LVT U5315 ( .A1(i_data_bus[329]), .A2(n5422), .B1(
        i_data_bus[361]), .B2(n5423), .ZN(n4957) );
  AOI22D1BWP30P140LVT U5316 ( .A1(i_data_bus[265]), .A2(n5394), .B1(
        i_data_bus[841]), .B2(n5425), .ZN(n4956) );
  AOI22D1BWP30P140LVT U5317 ( .A1(i_data_bus[617]), .A2(n5416), .B1(
        i_data_bus[553]), .B2(n5417), .ZN(n4955) );
  AOI22D1BWP30P140LVT U5318 ( .A1(i_data_bus[521]), .A2(n5414), .B1(
        i_data_bus[585]), .B2(n5415), .ZN(n4954) );
  ND4D1BWP30P140LVT U5319 ( .A1(n4957), .A2(n4956), .A3(n4955), .A4(n4954), 
        .ZN(n4963) );
  AOI22D1BWP30P140LVT U5320 ( .A1(i_data_bus[713]), .A2(n5424), .B1(
        i_data_bus[457]), .B2(n222), .ZN(n4961) );
  AOI22D1BWP30P140LVT U5321 ( .A1(i_data_bus[745]), .A2(n5412), .B1(
        i_data_bus[681]), .B2(n5393), .ZN(n4960) );
  AOI22D1BWP30P140LVT U5322 ( .A1(i_data_bus[393]), .A2(n5411), .B1(
        i_data_bus[649]), .B2(n5426), .ZN(n4959) );
  AOI22D1BWP30P140LVT U5323 ( .A1(i_data_bus[873]), .A2(n5410), .B1(
        i_data_bus[425]), .B2(n5413), .ZN(n4958) );
  ND4D1BWP30P140LVT U5324 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), 
        .ZN(n4962) );
  NR4D0BWP30P140LVT U5325 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), 
        .ZN(n4966) );
  ND4D1BWP30P140LVT U5326 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), 
        .ZN(o_data_bus[9]) );
  AOI22D1BWP30P140LVT U5327 ( .A1(i_data_bus[74]), .A2(n5390), .B1(
        i_data_bus[170]), .B2(n5391), .ZN(n4989) );
  AOI22D1BWP30P140LVT U5328 ( .A1(i_data_bus[1002]), .A2(n5396), .B1(
        i_data_bus[202]), .B2(n5400), .ZN(n4988) );
  AOI22D1BWP30P140LVT U5329 ( .A1(i_data_bus[298]), .A2(n5428), .B1(
        i_data_bus[426]), .B2(n5413), .ZN(n4987) );
  AOI22D1BWP30P140LVT U5330 ( .A1(i_data_bus[42]), .A2(n5395), .B1(
        i_data_bus[906]), .B2(n5389), .ZN(n4973) );
  AOI22D1BWP30P140LVT U5331 ( .A1(i_data_bus[10]), .A2(n5398), .B1(
        i_data_bus[138]), .B2(n5399), .ZN(n4972) );
  AOI22D1BWP30P140LVT U5332 ( .A1(i_data_bus[106]), .A2(n5402), .B1(
        i_data_bus[938]), .B2(n5397), .ZN(n4971) );
  AOI22D1BWP30P140LVT U5333 ( .A1(i_data_bus[970]), .A2(n5392), .B1(
        i_data_bus[234]), .B2(n5401), .ZN(n4970) );
  ND4D1BWP30P140LVT U5334 ( .A1(n4973), .A2(n4972), .A3(n4971), .A4(n4970), 
        .ZN(n4985) );
  MOAI22D1BWP30P140LVT U5335 ( .A1(n5706), .A2(n5308), .B1(i_data_bus[458]), 
        .B2(n222), .ZN(n4984) );
  AOI22D1BWP30P140LVT U5336 ( .A1(i_data_bus[778]), .A2(n5407), .B1(
        i_data_bus[842]), .B2(n5425), .ZN(n4977) );
  AOI22D1BWP30P140LVT U5337 ( .A1(i_data_bus[874]), .A2(n5410), .B1(
        i_data_bus[746]), .B2(n5412), .ZN(n4976) );
  AOI22D1BWP30P140LVT U5338 ( .A1(i_data_bus[618]), .A2(n5416), .B1(
        i_data_bus[586]), .B2(n5415), .ZN(n4975) );
  AOI22D1BWP30P140LVT U5339 ( .A1(i_data_bus[554]), .A2(n5417), .B1(
        i_data_bus[522]), .B2(n5414), .ZN(n4974) );
  ND4D1BWP30P140LVT U5340 ( .A1(n4977), .A2(n4976), .A3(n4975), .A4(n4974), 
        .ZN(n4983) );
  AOI22D1BWP30P140LVT U5341 ( .A1(i_data_bus[362]), .A2(n5423), .B1(
        i_data_bus[266]), .B2(n5394), .ZN(n4981) );
  AOI22D1BWP30P140LVT U5342 ( .A1(i_data_bus[810]), .A2(n5427), .B1(
        i_data_bus[682]), .B2(n5393), .ZN(n4980) );
  AOI22D1BWP30P140LVT U5343 ( .A1(i_data_bus[330]), .A2(n5422), .B1(
        i_data_bus[714]), .B2(n5424), .ZN(n4979) );
  AOI22D1BWP30P140LVT U5344 ( .A1(i_data_bus[650]), .A2(n5426), .B1(
        i_data_bus[394]), .B2(n5411), .ZN(n4978) );
  ND4D1BWP30P140LVT U5345 ( .A1(n4981), .A2(n4980), .A3(n4979), .A4(n4978), 
        .ZN(n4982) );
  NR4D0BWP30P140LVT U5346 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), 
        .ZN(n4986) );
  ND4D1BWP30P140LVT U5347 ( .A1(n4989), .A2(n4988), .A3(n4987), .A4(n4986), 
        .ZN(o_data_bus[10]) );
  AOI22D1BWP30P140LVT U5348 ( .A1(i_data_bus[907]), .A2(n5389), .B1(
        i_data_bus[971]), .B2(n5392), .ZN(n5009) );
  AOI22D1BWP30P140LVT U5349 ( .A1(i_data_bus[1003]), .A2(n5396), .B1(
        i_data_bus[75]), .B2(n5390), .ZN(n5008) );
  AOI22D1BWP30P140LVT U5350 ( .A1(i_data_bus[875]), .A2(n5410), .B1(
        i_data_bus[843]), .B2(n5425), .ZN(n5007) );
  AOI22D1BWP30P140LVT U5351 ( .A1(i_data_bus[107]), .A2(n5402), .B1(
        i_data_bus[203]), .B2(n5400), .ZN(n4993) );
  AOI22D1BWP30P140LVT U5352 ( .A1(i_data_bus[939]), .A2(n5397), .B1(
        i_data_bus[11]), .B2(n5398), .ZN(n4992) );
  AOI22D1BWP30P140LVT U5353 ( .A1(i_data_bus[171]), .A2(n5391), .B1(
        i_data_bus[235]), .B2(n5401), .ZN(n4991) );
  AOI22D1BWP30P140LVT U5354 ( .A1(i_data_bus[43]), .A2(n5395), .B1(
        i_data_bus[139]), .B2(n5399), .ZN(n4990) );
  ND4D1BWP30P140LVT U5355 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), 
        .ZN(n5005) );
  MOAI22D1BWP30P140LVT U5356 ( .A1(n5729), .A2(n5408), .B1(i_data_bus[747]), 
        .B2(n5412), .ZN(n5004) );
  AOI22D1BWP30P140LVT U5357 ( .A1(i_data_bus[651]), .A2(n5426), .B1(
        i_data_bus[683]), .B2(n5393), .ZN(n4997) );
  AOI22D1BWP30P140LVT U5358 ( .A1(i_data_bus[427]), .A2(n5413), .B1(
        i_data_bus[715]), .B2(n5424), .ZN(n4996) );
  AOI22D1BWP30P140LVT U5359 ( .A1(i_data_bus[619]), .A2(n5416), .B1(
        i_data_bus[587]), .B2(n5415), .ZN(n4995) );
  AOI22D1BWP30P140LVT U5360 ( .A1(i_data_bus[523]), .A2(n5414), .B1(
        i_data_bus[555]), .B2(n5417), .ZN(n4994) );
  ND4D1BWP30P140LVT U5361 ( .A1(n4997), .A2(n4996), .A3(n4995), .A4(n4994), 
        .ZN(n5003) );
  AOI22D1BWP30P140LVT U5362 ( .A1(i_data_bus[395]), .A2(n5411), .B1(
        i_data_bus[811]), .B2(n5427), .ZN(n5001) );
  AOI22D1BWP30P140LVT U5363 ( .A1(i_data_bus[363]), .A2(n5423), .B1(
        i_data_bus[267]), .B2(n5394), .ZN(n5000) );
  AOI22D1BWP30P140LVT U5364 ( .A1(i_data_bus[779]), .A2(n5407), .B1(
        i_data_bus[299]), .B2(n5428), .ZN(n4999) );
  AOI22D1BWP30P140LVT U5365 ( .A1(i_data_bus[491]), .A2(n223), .B1(
        i_data_bus[331]), .B2(n5422), .ZN(n4998) );
  ND4D1BWP30P140LVT U5366 ( .A1(n5001), .A2(n5000), .A3(n4999), .A4(n4998), 
        .ZN(n5002) );
  NR4D0BWP30P140LVT U5367 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5002), 
        .ZN(n5006) );
  ND4D1BWP30P140LVT U5368 ( .A1(n5009), .A2(n5008), .A3(n5007), .A4(n5006), 
        .ZN(o_data_bus[11]) );
  AOI22D1BWP30P140LVT U5369 ( .A1(i_data_bus[12]), .A2(n5398), .B1(
        i_data_bus[140]), .B2(n5399), .ZN(n5031) );
  AOI22D1BWP30P140LVT U5370 ( .A1(i_data_bus[1004]), .A2(n5396), .B1(
        i_data_bus[108]), .B2(n5402), .ZN(n5030) );
  AOI22D1BWP30P140LVT U5371 ( .A1(i_data_bus[780]), .A2(n5407), .B1(
        i_data_bus[332]), .B2(n5422), .ZN(n5029) );
  AOI22D1BWP30P140LVT U5372 ( .A1(i_data_bus[76]), .A2(n5390), .B1(
        i_data_bus[204]), .B2(n5400), .ZN(n5013) );
  AOI22D1BWP30P140LVT U5373 ( .A1(i_data_bus[908]), .A2(n5389), .B1(
        i_data_bus[972]), .B2(n5392), .ZN(n5012) );
  AOI22D1BWP30P140LVT U5374 ( .A1(i_data_bus[940]), .A2(n5397), .B1(
        i_data_bus[172]), .B2(n5391), .ZN(n5011) );
  AOI22D1BWP30P140LVT U5375 ( .A1(i_data_bus[44]), .A2(n5395), .B1(
        i_data_bus[236]), .B2(n5401), .ZN(n5010) );
  ND4D1BWP30P140LVT U5376 ( .A1(n5013), .A2(n5012), .A3(n5011), .A4(n5010), 
        .ZN(n5027) );
  OAI22D1BWP30P140LVT U5377 ( .A1(n5015), .A2(n5408), .B1(n5014), .B2(n5308), 
        .ZN(n5026) );
  AOI22D1BWP30P140LVT U5378 ( .A1(i_data_bus[652]), .A2(n5426), .B1(
        i_data_bus[876]), .B2(n5410), .ZN(n5019) );
  AOI22D1BWP30P140LVT U5379 ( .A1(i_data_bus[684]), .A2(n5393), .B1(
        i_data_bus[812]), .B2(n5427), .ZN(n5018) );
  AOI22D1BWP30P140LVT U5380 ( .A1(i_data_bus[556]), .A2(n5417), .B1(
        i_data_bus[524]), .B2(n5414), .ZN(n5017) );
  AOI22D1BWP30P140LVT U5381 ( .A1(i_data_bus[620]), .A2(n5416), .B1(
        i_data_bus[588]), .B2(n5415), .ZN(n5016) );
  ND4D1BWP30P140LVT U5382 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), 
        .ZN(n5025) );
  AOI22D1BWP30P140LVT U5383 ( .A1(i_data_bus[300]), .A2(n5428), .B1(
        i_data_bus[364]), .B2(n5423), .ZN(n5023) );
  AOI22D1BWP30P140LVT U5384 ( .A1(i_data_bus[428]), .A2(n5413), .B1(
        i_data_bus[268]), .B2(n5394), .ZN(n5022) );
  AOI22D1BWP30P140LVT U5385 ( .A1(i_data_bus[748]), .A2(n5412), .B1(
        i_data_bus[396]), .B2(n5411), .ZN(n5021) );
  AOI22D1BWP30P140LVT U5386 ( .A1(i_data_bus[716]), .A2(n5424), .B1(
        i_data_bus[844]), .B2(n5425), .ZN(n5020) );
  ND4D1BWP30P140LVT U5387 ( .A1(n5023), .A2(n5022), .A3(n5021), .A4(n5020), 
        .ZN(n5024) );
  NR4D0BWP30P140LVT U5388 ( .A1(n5027), .A2(n5026), .A3(n5025), .A4(n5024), 
        .ZN(n5028) );
  ND4D1BWP30P140LVT U5389 ( .A1(n5031), .A2(n5030), .A3(n5029), .A4(n5028), 
        .ZN(o_data_bus[12]) );
  AOI22D1BWP30P140LVT U5390 ( .A1(i_data_bus[109]), .A2(n5402), .B1(
        i_data_bus[173]), .B2(n5391), .ZN(n5052) );
  AOI22D1BWP30P140LVT U5391 ( .A1(i_data_bus[237]), .A2(n5401), .B1(
        i_data_bus[141]), .B2(n5399), .ZN(n5051) );
  AOI22D1BWP30P140LVT U5392 ( .A1(i_data_bus[333]), .A2(n5422), .B1(
        i_data_bus[813]), .B2(n5427), .ZN(n5050) );
  AOI22D1BWP30P140LVT U5393 ( .A1(i_data_bus[45]), .A2(n5395), .B1(
        i_data_bus[77]), .B2(n5390), .ZN(n5035) );
  AOI22D1BWP30P140LVT U5394 ( .A1(i_data_bus[909]), .A2(n5389), .B1(
        i_data_bus[941]), .B2(n5397), .ZN(n5034) );
  AOI22D1BWP30P140LVT U5395 ( .A1(i_data_bus[1005]), .A2(n5396), .B1(
        i_data_bus[13]), .B2(n5398), .ZN(n5033) );
  AOI22D1BWP30P140LVT U5396 ( .A1(i_data_bus[973]), .A2(n5392), .B1(
        i_data_bus[205]), .B2(n5400), .ZN(n5032) );
  ND4D1BWP30P140LVT U5397 ( .A1(n5035), .A2(n5034), .A3(n5033), .A4(n5032), 
        .ZN(n5048) );
  MOAI22D1BWP30P140LVT U5398 ( .A1(n5036), .A2(n5308), .B1(i_data_bus[877]), 
        .B2(n5410), .ZN(n5047) );
  AOI22D1BWP30P140LVT U5399 ( .A1(i_data_bus[429]), .A2(n5413), .B1(
        i_data_bus[845]), .B2(n5425), .ZN(n5040) );
  AOI22D1BWP30P140LVT U5400 ( .A1(i_data_bus[653]), .A2(n5426), .B1(
        i_data_bus[461]), .B2(n222), .ZN(n5039) );
  AOI22D1BWP30P140LVT U5401 ( .A1(i_data_bus[621]), .A2(n5416), .B1(
        i_data_bus[589]), .B2(n5415), .ZN(n5038) );
  AOI22D1BWP30P140LVT U5402 ( .A1(i_data_bus[525]), .A2(n5414), .B1(
        i_data_bus[557]), .B2(n5417), .ZN(n5037) );
  ND4D1BWP30P140LVT U5403 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n5037), 
        .ZN(n5046) );
  AOI22D1BWP30P140LVT U5404 ( .A1(i_data_bus[397]), .A2(n5411), .B1(
        i_data_bus[717]), .B2(n5424), .ZN(n5044) );
  AOI22D1BWP30P140LVT U5405 ( .A1(i_data_bus[269]), .A2(n5394), .B1(
        i_data_bus[781]), .B2(n5407), .ZN(n5043) );
  AOI22D1BWP30P140LVT U5406 ( .A1(i_data_bus[365]), .A2(n5423), .B1(
        i_data_bus[301]), .B2(n5428), .ZN(n5042) );
  AOI22D1BWP30P140LVT U5407 ( .A1(i_data_bus[749]), .A2(n5412), .B1(
        i_data_bus[685]), .B2(n5393), .ZN(n5041) );
  ND4D1BWP30P140LVT U5408 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), 
        .ZN(n5045) );
  NR4D0BWP30P140LVT U5409 ( .A1(n5048), .A2(n5047), .A3(n5046), .A4(n5045), 
        .ZN(n5049) );
  ND4D1BWP30P140LVT U5410 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), 
        .ZN(o_data_bus[13]) );
  AOI22D1BWP30P140LVT U5411 ( .A1(i_data_bus[910]), .A2(n5389), .B1(
        i_data_bus[14]), .B2(n5398), .ZN(n5072) );
  AOI22D1BWP30P140LVT U5412 ( .A1(i_data_bus[974]), .A2(n5392), .B1(
        i_data_bus[142]), .B2(n5399), .ZN(n5071) );
  AOI22D1BWP30P140LVT U5413 ( .A1(i_data_bus[462]), .A2(n222), .B1(
        i_data_bus[398]), .B2(n5411), .ZN(n5070) );
  AOI22D1BWP30P140LVT U5414 ( .A1(i_data_bus[334]), .A2(n5422), .B1(
        i_data_bus[878]), .B2(n5410), .ZN(n5068) );
  AOI22D1BWP30P140LVT U5415 ( .A1(i_data_bus[1006]), .A2(n5396), .B1(
        i_data_bus[942]), .B2(n5397), .ZN(n5056) );
  AOI22D1BWP30P140LVT U5416 ( .A1(i_data_bus[46]), .A2(n5395), .B1(
        i_data_bus[206]), .B2(n5400), .ZN(n5055) );
  AOI22D1BWP30P140LVT U5417 ( .A1(i_data_bus[78]), .A2(n5390), .B1(
        i_data_bus[174]), .B2(n5391), .ZN(n5054) );
  AOI22D1BWP30P140LVT U5418 ( .A1(i_data_bus[110]), .A2(n5402), .B1(
        i_data_bus[238]), .B2(n5401), .ZN(n5053) );
  ND4D1BWP30P140LVT U5419 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), 
        .ZN(n5067) );
  AOI22D1BWP30P140LVT U5420 ( .A1(i_data_bus[846]), .A2(n5425), .B1(
        i_data_bus[302]), .B2(n5428), .ZN(n5060) );
  AOI22D1BWP30P140LVT U5421 ( .A1(i_data_bus[270]), .A2(n5394), .B1(
        i_data_bus[814]), .B2(n5427), .ZN(n5059) );
  AOI22D1BWP30P140LVT U5422 ( .A1(i_data_bus[558]), .A2(n5417), .B1(
        i_data_bus[622]), .B2(n5416), .ZN(n5058) );
  AOI22D1BWP30P140LVT U5423 ( .A1(i_data_bus[590]), .A2(n5415), .B1(
        i_data_bus[526]), .B2(n5414), .ZN(n5057) );
  ND4D1BWP30P140LVT U5424 ( .A1(n5060), .A2(n5059), .A3(n5058), .A4(n5057), 
        .ZN(n5066) );
  AOI22D1BWP30P140LVT U5425 ( .A1(i_data_bus[686]), .A2(n5393), .B1(
        i_data_bus[718]), .B2(n5424), .ZN(n5064) );
  AOI22D1BWP30P140LVT U5426 ( .A1(i_data_bus[782]), .A2(n5407), .B1(
        i_data_bus[430]), .B2(n5413), .ZN(n5063) );
  AOI22D1BWP30P140LVT U5427 ( .A1(i_data_bus[366]), .A2(n5423), .B1(
        i_data_bus[494]), .B2(n223), .ZN(n5062) );
  AOI22D1BWP30P140LVT U5428 ( .A1(i_data_bus[750]), .A2(n5412), .B1(
        i_data_bus[654]), .B2(n5426), .ZN(n5061) );
  ND4D1BWP30P140LVT U5429 ( .A1(n5064), .A2(n5063), .A3(n5062), .A4(n5061), 
        .ZN(n5065) );
  INR4D0BWP30P140LVT U5430 ( .A1(n5068), .B1(n5067), .B2(n5066), .B3(n5065), 
        .ZN(n5069) );
  ND4D1BWP30P140LVT U5431 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), 
        .ZN(o_data_bus[14]) );
  AOI22D1BWP30P140LVT U5432 ( .A1(i_data_bus[943]), .A2(n5397), .B1(
        i_data_bus[207]), .B2(n5400), .ZN(n5093) );
  AOI22D1BWP30P140LVT U5433 ( .A1(i_data_bus[975]), .A2(n5392), .B1(
        i_data_bus[175]), .B2(n5391), .ZN(n5092) );
  AOI22D1BWP30P140LVT U5434 ( .A1(i_data_bus[783]), .A2(n5407), .B1(
        i_data_bus[335]), .B2(n5422), .ZN(n5091) );
  AOI22D1BWP30P140LVT U5435 ( .A1(i_data_bus[111]), .A2(n5402), .B1(
        i_data_bus[1007]), .B2(n5396), .ZN(n5076) );
  AOI22D1BWP30P140LVT U5436 ( .A1(i_data_bus[911]), .A2(n5389), .B1(
        i_data_bus[15]), .B2(n5398), .ZN(n5075) );
  AOI22D1BWP30P140LVT U5437 ( .A1(i_data_bus[239]), .A2(n5401), .B1(
        i_data_bus[143]), .B2(n5399), .ZN(n5074) );
  AOI22D1BWP30P140LVT U5438 ( .A1(i_data_bus[79]), .A2(n5390), .B1(
        i_data_bus[47]), .B2(n5395), .ZN(n5073) );
  ND4D1BWP30P140LVT U5439 ( .A1(n5076), .A2(n5075), .A3(n5074), .A4(n5073), 
        .ZN(n5089) );
  MOAI22D1BWP30P140LVT U5440 ( .A1(n5077), .A2(n228), .B1(i_data_bus[655]), 
        .B2(n5426), .ZN(n5088) );
  AOI22D1BWP30P140LVT U5441 ( .A1(i_data_bus[719]), .A2(n5424), .B1(
        i_data_bus[687]), .B2(n5393), .ZN(n5081) );
  AOI22D1BWP30P140LVT U5442 ( .A1(i_data_bus[847]), .A2(n5425), .B1(
        i_data_bus[303]), .B2(n5428), .ZN(n5080) );
  AOI22D1BWP30P140LVT U5443 ( .A1(i_data_bus[527]), .A2(n5414), .B1(
        i_data_bus[623]), .B2(n5416), .ZN(n5079) );
  AOI22D1BWP30P140LVT U5444 ( .A1(i_data_bus[591]), .A2(n5415), .B1(
        i_data_bus[559]), .B2(n5417), .ZN(n5078) );
  ND4D1BWP30P140LVT U5445 ( .A1(n5081), .A2(n5080), .A3(n5079), .A4(n5078), 
        .ZN(n5087) );
  AOI22D1BWP30P140LVT U5446 ( .A1(i_data_bus[495]), .A2(n223), .B1(
        i_data_bus[879]), .B2(n5410), .ZN(n5085) );
  AOI22D1BWP30P140LVT U5447 ( .A1(i_data_bus[815]), .A2(n5427), .B1(
        i_data_bus[367]), .B2(n5423), .ZN(n5084) );
  AOI22D1BWP30P140LVT U5448 ( .A1(i_data_bus[271]), .A2(n5394), .B1(
        i_data_bus[463]), .B2(n222), .ZN(n5083) );
  AOI22D1BWP30P140LVT U5449 ( .A1(i_data_bus[751]), .A2(n5412), .B1(
        i_data_bus[431]), .B2(n5413), .ZN(n5082) );
  ND4D1BWP30P140LVT U5450 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), 
        .ZN(n5086) );
  NR4D0BWP30P140LVT U5451 ( .A1(n5089), .A2(n5088), .A3(n5087), .A4(n5086), 
        .ZN(n5090) );
  ND4D1BWP30P140LVT U5452 ( .A1(n5093), .A2(n5092), .A3(n5091), .A4(n5090), 
        .ZN(o_data_bus[15]) );
  AOI22D1BWP30P140LVT U5453 ( .A1(i_data_bus[976]), .A2(n5392), .B1(
        i_data_bus[16]), .B2(n5398), .ZN(n5113) );
  AOI22D1BWP30P140LVT U5454 ( .A1(i_data_bus[912]), .A2(n5389), .B1(
        i_data_bus[1008]), .B2(n5396), .ZN(n5112) );
  AOI22D1BWP30P140LVT U5455 ( .A1(i_data_bus[304]), .A2(n5428), .B1(
        i_data_bus[656]), .B2(n5426), .ZN(n5111) );
  AOI22D1BWP30P140LVT U5456 ( .A1(i_data_bus[144]), .A2(n5399), .B1(
        i_data_bus[176]), .B2(n5391), .ZN(n5097) );
  AOI22D1BWP30P140LVT U5457 ( .A1(i_data_bus[48]), .A2(n5395), .B1(
        i_data_bus[240]), .B2(n5401), .ZN(n5096) );
  AOI22D1BWP30P140LVT U5458 ( .A1(i_data_bus[80]), .A2(n5390), .B1(
        i_data_bus[112]), .B2(n5402), .ZN(n5095) );
  AOI22D1BWP30P140LVT U5459 ( .A1(i_data_bus[944]), .A2(n5397), .B1(
        i_data_bus[208]), .B2(n5400), .ZN(n5094) );
  ND4D1BWP30P140LVT U5460 ( .A1(n5097), .A2(n5096), .A3(n5095), .A4(n5094), 
        .ZN(n5109) );
  MOAI22D1BWP30P140LVT U5461 ( .A1(n5834), .A2(n228), .B1(i_data_bus[880]), 
        .B2(n5410), .ZN(n5108) );
  AOI22D1BWP30P140LVT U5462 ( .A1(i_data_bus[464]), .A2(n222), .B1(
        i_data_bus[688]), .B2(n5393), .ZN(n5101) );
  AOI22D1BWP30P140LVT U5463 ( .A1(i_data_bus[336]), .A2(n5422), .B1(
        i_data_bus[720]), .B2(n5424), .ZN(n5100) );
  AOI22D1BWP30P140LVT U5464 ( .A1(i_data_bus[560]), .A2(n5417), .B1(
        i_data_bus[624]), .B2(n5416), .ZN(n5099) );
  AOI22D1BWP30P140LVT U5465 ( .A1(i_data_bus[528]), .A2(n5414), .B1(
        i_data_bus[592]), .B2(n5415), .ZN(n5098) );
  ND4D1BWP30P140LVT U5466 ( .A1(n5101), .A2(n5100), .A3(n5099), .A4(n5098), 
        .ZN(n5107) );
  AOI22D1BWP30P140LVT U5467 ( .A1(i_data_bus[784]), .A2(n5407), .B1(
        i_data_bus[272]), .B2(n5394), .ZN(n5105) );
  AOI22D1BWP30P140LVT U5468 ( .A1(i_data_bus[816]), .A2(n5427), .B1(
        i_data_bus[848]), .B2(n5425), .ZN(n5104) );
  AOI22D1BWP30P140LVT U5469 ( .A1(i_data_bus[496]), .A2(n223), .B1(
        i_data_bus[368]), .B2(n5423), .ZN(n5103) );
  AOI22D1BWP30P140LVT U5470 ( .A1(i_data_bus[432]), .A2(n5413), .B1(
        i_data_bus[752]), .B2(n5412), .ZN(n5102) );
  ND4D1BWP30P140LVT U5471 ( .A1(n5105), .A2(n5104), .A3(n5103), .A4(n5102), 
        .ZN(n5106) );
  NR4D0BWP30P140LVT U5472 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), 
        .ZN(n5110) );
  ND4D1BWP30P140LVT U5473 ( .A1(n5113), .A2(n5112), .A3(n5111), .A4(n5110), 
        .ZN(o_data_bus[16]) );
  AOI22D1BWP30P140LVT U5474 ( .A1(i_data_bus[913]), .A2(n5389), .B1(
        i_data_bus[145]), .B2(n5399), .ZN(n5133) );
  AOI22D1BWP30P140LVT U5475 ( .A1(i_data_bus[1009]), .A2(n5396), .B1(
        i_data_bus[209]), .B2(n5400), .ZN(n5132) );
  AOI22D1BWP30P140LVT U5476 ( .A1(i_data_bus[721]), .A2(n5424), .B1(
        i_data_bus[273]), .B2(n5394), .ZN(n5131) );
  AOI22D1BWP30P140LVT U5477 ( .A1(i_data_bus[689]), .A2(n5393), .B1(
        i_data_bus[465]), .B2(n222), .ZN(n5129) );
  AOI22D1BWP30P140LVT U5478 ( .A1(i_data_bus[17]), .A2(n5398), .B1(
        i_data_bus[177]), .B2(n5391), .ZN(n5117) );
  AOI22D1BWP30P140LVT U5479 ( .A1(i_data_bus[49]), .A2(n5395), .B1(
        i_data_bus[945]), .B2(n5397), .ZN(n5116) );
  AOI22D1BWP30P140LVT U5480 ( .A1(i_data_bus[977]), .A2(n5392), .B1(
        i_data_bus[241]), .B2(n5401), .ZN(n5115) );
  AOI22D1BWP30P140LVT U5481 ( .A1(i_data_bus[81]), .A2(n5390), .B1(
        i_data_bus[113]), .B2(n5402), .ZN(n5114) );
  ND4D1BWP30P140LVT U5482 ( .A1(n5117), .A2(n5116), .A3(n5115), .A4(n5114), 
        .ZN(n5128) );
  AOI22D1BWP30P140LVT U5483 ( .A1(i_data_bus[753]), .A2(n5412), .B1(
        i_data_bus[497]), .B2(n223), .ZN(n5121) );
  AOI22D1BWP30P140LVT U5484 ( .A1(i_data_bus[433]), .A2(n5413), .B1(
        i_data_bus[401]), .B2(n5411), .ZN(n5120) );
  AOI22D1BWP30P140LVT U5485 ( .A1(i_data_bus[625]), .A2(n5416), .B1(
        i_data_bus[561]), .B2(n5417), .ZN(n5119) );
  AOI22D1BWP30P140LVT U5486 ( .A1(i_data_bus[593]), .A2(n5415), .B1(
        i_data_bus[529]), .B2(n5414), .ZN(n5118) );
  ND4D1BWP30P140LVT U5487 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), 
        .ZN(n5127) );
  AOI22D1BWP30P140LVT U5488 ( .A1(i_data_bus[305]), .A2(n5428), .B1(
        i_data_bus[369]), .B2(n5423), .ZN(n5125) );
  AOI22D1BWP30P140LVT U5489 ( .A1(i_data_bus[337]), .A2(n5422), .B1(
        i_data_bus[785]), .B2(n5407), .ZN(n5124) );
  AOI22D1BWP30P140LVT U5490 ( .A1(i_data_bus[849]), .A2(n5425), .B1(
        i_data_bus[817]), .B2(n5427), .ZN(n5123) );
  AOI22D1BWP30P140LVT U5491 ( .A1(i_data_bus[881]), .A2(n5410), .B1(
        i_data_bus[657]), .B2(n5426), .ZN(n5122) );
  ND4D1BWP30P140LVT U5492 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), 
        .ZN(n5126) );
  INR4D0BWP30P140LVT U5493 ( .A1(n5129), .B1(n5128), .B2(n5127), .B3(n5126), 
        .ZN(n5130) );
  ND4D1BWP30P140LVT U5494 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), 
        .ZN(o_data_bus[17]) );
  AOI22D1BWP30P140LVT U5495 ( .A1(i_data_bus[82]), .A2(n5390), .B1(
        i_data_bus[914]), .B2(n5389), .ZN(n5153) );
  AOI22D1BWP30P140LVT U5496 ( .A1(i_data_bus[946]), .A2(n5397), .B1(
        i_data_bus[210]), .B2(n5400), .ZN(n5152) );
  AOI22D1BWP30P140LVT U5497 ( .A1(i_data_bus[370]), .A2(n5423), .B1(
        i_data_bus[306]), .B2(n5428), .ZN(n5151) );
  AOI22D1BWP30P140LVT U5498 ( .A1(i_data_bus[882]), .A2(n5410), .B1(
        i_data_bus[722]), .B2(n5424), .ZN(n5149) );
  AOI22D1BWP30P140LVT U5499 ( .A1(i_data_bus[978]), .A2(n5392), .B1(
        i_data_bus[114]), .B2(n5402), .ZN(n5137) );
  AOI22D1BWP30P140LVT U5500 ( .A1(i_data_bus[1010]), .A2(n5396), .B1(
        i_data_bus[146]), .B2(n5399), .ZN(n5136) );
  AOI22D1BWP30P140LVT U5501 ( .A1(i_data_bus[50]), .A2(n5395), .B1(
        i_data_bus[18]), .B2(n5398), .ZN(n5135) );
  AOI22D1BWP30P140LVT U5502 ( .A1(i_data_bus[242]), .A2(n5401), .B1(
        i_data_bus[178]), .B2(n5391), .ZN(n5134) );
  ND4D1BWP30P140LVT U5503 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), 
        .ZN(n5148) );
  AOI22D1BWP30P140LVT U5504 ( .A1(i_data_bus[818]), .A2(n5427), .B1(
        i_data_bus[498]), .B2(n223), .ZN(n5141) );
  AOI22D1BWP30P140LVT U5505 ( .A1(i_data_bus[690]), .A2(n5393), .B1(
        i_data_bus[274]), .B2(n5394), .ZN(n5140) );
  AOI22D1BWP30P140LVT U5506 ( .A1(i_data_bus[530]), .A2(n5414), .B1(
        i_data_bus[562]), .B2(n5417), .ZN(n5139) );
  AOI22D1BWP30P140LVT U5507 ( .A1(i_data_bus[626]), .A2(n5416), .B1(
        i_data_bus[594]), .B2(n5415), .ZN(n5138) );
  ND4D1BWP30P140LVT U5508 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), 
        .ZN(n5147) );
  AOI22D1BWP30P140LVT U5509 ( .A1(i_data_bus[466]), .A2(n222), .B1(
        i_data_bus[754]), .B2(n5412), .ZN(n5145) );
  AOI22D1BWP30P140LVT U5510 ( .A1(i_data_bus[402]), .A2(n5411), .B1(
        i_data_bus[850]), .B2(n5425), .ZN(n5144) );
  AOI22D1BWP30P140LVT U5511 ( .A1(i_data_bus[658]), .A2(n5426), .B1(
        i_data_bus[786]), .B2(n5407), .ZN(n5143) );
  AOI22D1BWP30P140LVT U5512 ( .A1(i_data_bus[434]), .A2(n5413), .B1(
        i_data_bus[338]), .B2(n5422), .ZN(n5142) );
  ND4D1BWP30P140LVT U5513 ( .A1(n5145), .A2(n5144), .A3(n5143), .A4(n5142), 
        .ZN(n5146) );
  INR4D0BWP30P140LVT U5514 ( .A1(n5149), .B1(n5148), .B2(n5147), .B3(n5146), 
        .ZN(n5150) );
  ND4D1BWP30P140LVT U5515 ( .A1(n5153), .A2(n5152), .A3(n5151), .A4(n5150), 
        .ZN(o_data_bus[18]) );
  AOI22D1BWP30P140LVT U5516 ( .A1(i_data_bus[947]), .A2(n5397), .B1(
        i_data_bus[915]), .B2(n5389), .ZN(n5174) );
  AOI22D1BWP30P140LVT U5517 ( .A1(i_data_bus[51]), .A2(n5395), .B1(
        i_data_bus[243]), .B2(n5401), .ZN(n5173) );
  AOI22D1BWP30P140LVT U5518 ( .A1(i_data_bus[275]), .A2(n5394), .B1(
        i_data_bus[467]), .B2(n222), .ZN(n5172) );
  AOI22D1BWP30P140LVT U5519 ( .A1(i_data_bus[115]), .A2(n5402), .B1(
        i_data_bus[83]), .B2(n5390), .ZN(n5157) );
  AOI22D1BWP30P140LVT U5520 ( .A1(i_data_bus[1011]), .A2(n5396), .B1(
        i_data_bus[19]), .B2(n5398), .ZN(n5156) );
  AOI22D1BWP30P140LVT U5521 ( .A1(i_data_bus[979]), .A2(n5392), .B1(
        i_data_bus[211]), .B2(n5400), .ZN(n5155) );
  AOI22D1BWP30P140LVT U5522 ( .A1(i_data_bus[179]), .A2(n5391), .B1(
        i_data_bus[147]), .B2(n5399), .ZN(n5154) );
  ND4D1BWP30P140LVT U5523 ( .A1(n5157), .A2(n5156), .A3(n5155), .A4(n5154), 
        .ZN(n5170) );
  MOAI22D1BWP30P140LVT U5524 ( .A1(n5158), .A2(n5264), .B1(i_data_bus[371]), 
        .B2(n5423), .ZN(n5169) );
  AOI22D1BWP30P140LVT U5525 ( .A1(i_data_bus[403]), .A2(n5411), .B1(
        i_data_bus[691]), .B2(n5393), .ZN(n5162) );
  AOI22D1BWP30P140LVT U5526 ( .A1(i_data_bus[819]), .A2(n5427), .B1(
        i_data_bus[723]), .B2(n5424), .ZN(n5161) );
  AOI22D1BWP30P140LVT U5527 ( .A1(i_data_bus[563]), .A2(n5417), .B1(
        i_data_bus[627]), .B2(n5416), .ZN(n5160) );
  AOI22D1BWP30P140LVT U5528 ( .A1(i_data_bus[531]), .A2(n5414), .B1(
        i_data_bus[595]), .B2(n5415), .ZN(n5159) );
  ND4D1BWP30P140LVT U5529 ( .A1(n5162), .A2(n5161), .A3(n5160), .A4(n5159), 
        .ZN(n5168) );
  AOI22D1BWP30P140LVT U5530 ( .A1(i_data_bus[787]), .A2(n5407), .B1(
        i_data_bus[883]), .B2(n5410), .ZN(n5166) );
  AOI22D1BWP30P140LVT U5531 ( .A1(i_data_bus[755]), .A2(n5412), .B1(
        i_data_bus[659]), .B2(n5426), .ZN(n5165) );
  AOI22D1BWP30P140LVT U5532 ( .A1(i_data_bus[851]), .A2(n5425), .B1(
        i_data_bus[435]), .B2(n5413), .ZN(n5164) );
  AOI22D1BWP30P140LVT U5533 ( .A1(i_data_bus[339]), .A2(n5422), .B1(
        i_data_bus[499]), .B2(n223), .ZN(n5163) );
  ND4D1BWP30P140LVT U5534 ( .A1(n5166), .A2(n5165), .A3(n5164), .A4(n5163), 
        .ZN(n5167) );
  NR4D0BWP30P140LVT U5535 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), 
        .ZN(n5171) );
  ND4D1BWP30P140LVT U5536 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), 
        .ZN(o_data_bus[19]) );
  AOI22D1BWP30P140LVT U5537 ( .A1(i_data_bus[84]), .A2(n5390), .B1(
        i_data_bus[180]), .B2(n5391), .ZN(n5194) );
  AOI22D1BWP30P140LVT U5538 ( .A1(i_data_bus[948]), .A2(n5397), .B1(
        i_data_bus[244]), .B2(n5401), .ZN(n5193) );
  AOI22D1BWP30P140LVT U5539 ( .A1(i_data_bus[724]), .A2(n5424), .B1(
        i_data_bus[436]), .B2(n5413), .ZN(n5192) );
  AOI22D1BWP30P140LVT U5540 ( .A1(i_data_bus[660]), .A2(n5426), .B1(
        i_data_bus[404]), .B2(n5411), .ZN(n5190) );
  AOI22D1BWP30P140LVT U5541 ( .A1(i_data_bus[20]), .A2(n5398), .B1(
        i_data_bus[212]), .B2(n5400), .ZN(n5178) );
  AOI22D1BWP30P140LVT U5542 ( .A1(i_data_bus[116]), .A2(n5402), .B1(
        i_data_bus[148]), .B2(n5399), .ZN(n5177) );
  AOI22D1BWP30P140LVT U5543 ( .A1(i_data_bus[980]), .A2(n5392), .B1(
        i_data_bus[1012]), .B2(n5396), .ZN(n5176) );
  AOI22D1BWP30P140LVT U5544 ( .A1(i_data_bus[52]), .A2(n5395), .B1(
        i_data_bus[916]), .B2(n5389), .ZN(n5175) );
  ND4D1BWP30P140LVT U5545 ( .A1(n5178), .A2(n5177), .A3(n5176), .A4(n5175), 
        .ZN(n5189) );
  AOI22D1BWP30P140LVT U5546 ( .A1(i_data_bus[852]), .A2(n5425), .B1(
        i_data_bus[276]), .B2(n5394), .ZN(n5182) );
  AOI22D1BWP30P140LVT U5547 ( .A1(i_data_bus[756]), .A2(n5412), .B1(
        i_data_bus[500]), .B2(n223), .ZN(n5181) );
  AOI22D1BWP30P140LVT U5548 ( .A1(i_data_bus[596]), .A2(n5415), .B1(
        i_data_bus[532]), .B2(n5414), .ZN(n5180) );
  AOI22D1BWP30P140LVT U5549 ( .A1(i_data_bus[564]), .A2(n5417), .B1(
        i_data_bus[628]), .B2(n5416), .ZN(n5179) );
  ND4D1BWP30P140LVT U5550 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), 
        .ZN(n5188) );
  AOI22D1BWP30P140LVT U5551 ( .A1(i_data_bus[692]), .A2(n5393), .B1(
        i_data_bus[468]), .B2(n222), .ZN(n5186) );
  AOI22D1BWP30P140LVT U5552 ( .A1(i_data_bus[340]), .A2(n5422), .B1(
        i_data_bus[788]), .B2(n5407), .ZN(n5185) );
  AOI22D1BWP30P140LVT U5553 ( .A1(i_data_bus[820]), .A2(n5427), .B1(
        i_data_bus[308]), .B2(n5428), .ZN(n5184) );
  AOI22D1BWP30P140LVT U5554 ( .A1(i_data_bus[884]), .A2(n5410), .B1(
        i_data_bus[372]), .B2(n5423), .ZN(n5183) );
  ND4D1BWP30P140LVT U5555 ( .A1(n5186), .A2(n5185), .A3(n5184), .A4(n5183), 
        .ZN(n5187) );
  INR4D0BWP30P140LVT U5556 ( .A1(n5190), .B1(n5189), .B2(n5188), .B3(n5187), 
        .ZN(n5191) );
  ND4D1BWP30P140LVT U5557 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), 
        .ZN(o_data_bus[20]) );
  AOI22D1BWP30P140LVT U5558 ( .A1(i_data_bus[53]), .A2(n5395), .B1(
        i_data_bus[181]), .B2(n5391), .ZN(n5215) );
  AOI22D1BWP30P140LVT U5559 ( .A1(i_data_bus[117]), .A2(n5402), .B1(
        i_data_bus[21]), .B2(n5398), .ZN(n5214) );
  AOI22D1BWP30P140LVT U5560 ( .A1(i_data_bus[757]), .A2(n5412), .B1(
        i_data_bus[501]), .B2(n223), .ZN(n5213) );
  AOI22D1BWP30P140LVT U5561 ( .A1(i_data_bus[85]), .A2(n5390), .B1(
        i_data_bus[149]), .B2(n5399), .ZN(n5198) );
  AOI22D1BWP30P140LVT U5562 ( .A1(i_data_bus[213]), .A2(n5400), .B1(
        i_data_bus[245]), .B2(n5401), .ZN(n5197) );
  AOI22D1BWP30P140LVT U5563 ( .A1(i_data_bus[917]), .A2(n5389), .B1(
        i_data_bus[1013]), .B2(n5396), .ZN(n5196) );
  AOI22D1BWP30P140LVT U5564 ( .A1(i_data_bus[949]), .A2(n5397), .B1(
        i_data_bus[981]), .B2(n5392), .ZN(n5195) );
  ND4D1BWP30P140LVT U5565 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), 
        .ZN(n5211) );
  MOAI22D1BWP30P140LVT U5566 ( .A1(n5199), .A2(n5264), .B1(i_data_bus[725]), 
        .B2(n5424), .ZN(n5210) );
  AOI22D1BWP30P140LVT U5567 ( .A1(i_data_bus[341]), .A2(n5422), .B1(
        i_data_bus[277]), .B2(n5394), .ZN(n5203) );
  AOI22D1BWP30P140LVT U5568 ( .A1(i_data_bus[853]), .A2(n5425), .B1(
        i_data_bus[405]), .B2(n5411), .ZN(n5202) );
  AOI22D1BWP30P140LVT U5569 ( .A1(i_data_bus[597]), .A2(n5415), .B1(
        i_data_bus[565]), .B2(n5417), .ZN(n5201) );
  AOI22D1BWP30P140LVT U5570 ( .A1(i_data_bus[629]), .A2(n5416), .B1(
        i_data_bus[533]), .B2(n5414), .ZN(n5200) );
  ND4D1BWP30P140LVT U5571 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), 
        .ZN(n5209) );
  AOI22D1BWP30P140LVT U5572 ( .A1(i_data_bus[789]), .A2(n5407), .B1(
        i_data_bus[373]), .B2(n5423), .ZN(n5207) );
  AOI22D1BWP30P140LVT U5573 ( .A1(i_data_bus[821]), .A2(n5427), .B1(
        i_data_bus[437]), .B2(n5413), .ZN(n5206) );
  AOI22D1BWP30P140LVT U5574 ( .A1(i_data_bus[661]), .A2(n5426), .B1(
        i_data_bus[885]), .B2(n5410), .ZN(n5205) );
  AOI22D1BWP30P140LVT U5575 ( .A1(i_data_bus[693]), .A2(n5393), .B1(
        i_data_bus[469]), .B2(n222), .ZN(n5204) );
  ND4D1BWP30P140LVT U5576 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), 
        .ZN(n5208) );
  NR4D0BWP30P140LVT U5577 ( .A1(n5211), .A2(n5210), .A3(n5209), .A4(n5208), 
        .ZN(n5212) );
  ND4D1BWP30P140LVT U5578 ( .A1(n5215), .A2(n5214), .A3(n5213), .A4(n5212), 
        .ZN(o_data_bus[21]) );
  AOI22D1BWP30P140LVT U5579 ( .A1(i_data_bus[182]), .A2(n5391), .B1(
        i_data_bus[214]), .B2(n5400), .ZN(n5238) );
  AOI22D1BWP30P140LVT U5580 ( .A1(i_data_bus[54]), .A2(n5395), .B1(
        i_data_bus[22]), .B2(n5398), .ZN(n5237) );
  AOI22D1BWP30P140LVT U5581 ( .A1(i_data_bus[310]), .A2(n5428), .B1(
        i_data_bus[854]), .B2(n5425), .ZN(n5236) );
  AOI22D1BWP30P140LVT U5582 ( .A1(i_data_bus[918]), .A2(n5389), .B1(
        i_data_bus[950]), .B2(n5397), .ZN(n5219) );
  AOI22D1BWP30P140LVT U5583 ( .A1(i_data_bus[246]), .A2(n5401), .B1(
        i_data_bus[150]), .B2(n5399), .ZN(n5218) );
  AOI22D1BWP30P140LVT U5584 ( .A1(i_data_bus[118]), .A2(n5402), .B1(
        i_data_bus[86]), .B2(n5390), .ZN(n5217) );
  AOI22D1BWP30P140LVT U5585 ( .A1(i_data_bus[1014]), .A2(n5396), .B1(
        i_data_bus[982]), .B2(n5392), .ZN(n5216) );
  ND4D1BWP30P140LVT U5586 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), 
        .ZN(n5234) );
  OAI22D1BWP30P140LVT U5587 ( .A1(n5222), .A2(n5408), .B1(n5221), .B2(n5220), 
        .ZN(n5233) );
  AOI22D1BWP30P140LVT U5588 ( .A1(i_data_bus[438]), .A2(n5413), .B1(
        i_data_bus[374]), .B2(n5423), .ZN(n5226) );
  AOI22D1BWP30P140LVT U5589 ( .A1(i_data_bus[822]), .A2(n5427), .B1(
        i_data_bus[758]), .B2(n5412), .ZN(n5225) );
  AOI22D1BWP30P140LVT U5590 ( .A1(i_data_bus[534]), .A2(n5414), .B1(
        i_data_bus[598]), .B2(n5415), .ZN(n5224) );
  AOI22D1BWP30P140LVT U5591 ( .A1(i_data_bus[566]), .A2(n5417), .B1(
        i_data_bus[630]), .B2(n5416), .ZN(n5223) );
  ND4D1BWP30P140LVT U5592 ( .A1(n5226), .A2(n5225), .A3(n5224), .A4(n5223), 
        .ZN(n5232) );
  AOI22D1BWP30P140LVT U5593 ( .A1(i_data_bus[406]), .A2(n5411), .B1(
        i_data_bus[278]), .B2(n5394), .ZN(n5230) );
  AOI22D1BWP30P140LVT U5594 ( .A1(i_data_bus[790]), .A2(n5407), .B1(
        i_data_bus[502]), .B2(n223), .ZN(n5229) );
  AOI22D1BWP30P140LVT U5595 ( .A1(i_data_bus[726]), .A2(n5424), .B1(
        i_data_bus[886]), .B2(n5410), .ZN(n5228) );
  AOI22D1BWP30P140LVT U5596 ( .A1(i_data_bus[694]), .A2(n5393), .B1(
        i_data_bus[662]), .B2(n5426), .ZN(n5227) );
  ND4D1BWP30P140LVT U5597 ( .A1(n5230), .A2(n5229), .A3(n5228), .A4(n5227), 
        .ZN(n5231) );
  NR4D0BWP30P140LVT U5598 ( .A1(n5234), .A2(n5233), .A3(n5232), .A4(n5231), 
        .ZN(n5235) );
  ND4D1BWP30P140LVT U5599 ( .A1(n5238), .A2(n5237), .A3(n5236), .A4(n5235), 
        .ZN(o_data_bus[22]) );
  AOI22D1BWP30P140LVT U5600 ( .A1(i_data_bus[1015]), .A2(n5396), .B1(
        i_data_bus[951]), .B2(n5397), .ZN(n5259) );
  AOI22D1BWP30P140LVT U5601 ( .A1(i_data_bus[119]), .A2(n5402), .B1(
        i_data_bus[215]), .B2(n5400), .ZN(n5258) );
  AOI22D1BWP30P140LVT U5602 ( .A1(i_data_bus[503]), .A2(n223), .B1(
        i_data_bus[343]), .B2(n5422), .ZN(n5257) );
  AOI22D1BWP30P140LVT U5603 ( .A1(i_data_bus[55]), .A2(n5395), .B1(
        i_data_bus[919]), .B2(n5389), .ZN(n5242) );
  AOI22D1BWP30P140LVT U5604 ( .A1(i_data_bus[983]), .A2(n5392), .B1(
        i_data_bus[151]), .B2(n5399), .ZN(n5241) );
  AOI22D1BWP30P140LVT U5605 ( .A1(i_data_bus[23]), .A2(n5398), .B1(
        i_data_bus[183]), .B2(n5391), .ZN(n5240) );
  AOI22D1BWP30P140LVT U5606 ( .A1(i_data_bus[87]), .A2(n5390), .B1(
        i_data_bus[247]), .B2(n5401), .ZN(n5239) );
  ND4D1BWP30P140LVT U5607 ( .A1(n5242), .A2(n5241), .A3(n5240), .A4(n5239), 
        .ZN(n5255) );
  MOAI22D1BWP30P140LVT U5608 ( .A1(n5243), .A2(n5408), .B1(i_data_bus[823]), 
        .B2(n5427), .ZN(n5254) );
  AOI22D1BWP30P140LVT U5609 ( .A1(i_data_bus[759]), .A2(n5412), .B1(
        i_data_bus[407]), .B2(n5411), .ZN(n5247) );
  AOI22D1BWP30P140LVT U5610 ( .A1(i_data_bus[695]), .A2(n5393), .B1(
        i_data_bus[311]), .B2(n5428), .ZN(n5246) );
  AOI22D1BWP30P140LVT U5611 ( .A1(i_data_bus[631]), .A2(n5416), .B1(
        i_data_bus[599]), .B2(n5415), .ZN(n5245) );
  AOI22D1BWP30P140LVT U5612 ( .A1(i_data_bus[535]), .A2(n5414), .B1(
        i_data_bus[567]), .B2(n5417), .ZN(n5244) );
  ND4D1BWP30P140LVT U5613 ( .A1(n5247), .A2(n5246), .A3(n5245), .A4(n5244), 
        .ZN(n5253) );
  AOI22D1BWP30P140LVT U5614 ( .A1(i_data_bus[439]), .A2(n5413), .B1(
        i_data_bus[727]), .B2(n5424), .ZN(n5251) );
  AOI22D1BWP30P140LVT U5615 ( .A1(i_data_bus[887]), .A2(n5410), .B1(
        i_data_bus[279]), .B2(n5394), .ZN(n5250) );
  AOI22D1BWP30P140LVT U5616 ( .A1(i_data_bus[663]), .A2(n5426), .B1(
        i_data_bus[375]), .B2(n5423), .ZN(n5249) );
  AOI22D1BWP30P140LVT U5617 ( .A1(i_data_bus[791]), .A2(n5407), .B1(
        i_data_bus[855]), .B2(n5425), .ZN(n5248) );
  ND4D1BWP30P140LVT U5618 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), 
        .ZN(n5252) );
  NR4D0BWP30P140LVT U5619 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), 
        .ZN(n5256) );
  ND4D1BWP30P140LVT U5620 ( .A1(n5259), .A2(n5258), .A3(n5257), .A4(n5256), 
        .ZN(o_data_bus[23]) );
  AOI22D1BWP30P140LVT U5621 ( .A1(i_data_bus[152]), .A2(n5399), .B1(
        i_data_bus[184]), .B2(n5391), .ZN(n5281) );
  AOI22D1BWP30P140LVT U5622 ( .A1(i_data_bus[120]), .A2(n5402), .B1(
        i_data_bus[248]), .B2(n5401), .ZN(n5280) );
  AOI22D1BWP30P140LVT U5623 ( .A1(i_data_bus[408]), .A2(n5411), .B1(
        i_data_bus[664]), .B2(n5426), .ZN(n5279) );
  AOI22D1BWP30P140LVT U5624 ( .A1(i_data_bus[1016]), .A2(n5396), .B1(
        i_data_bus[24]), .B2(n5398), .ZN(n5263) );
  AOI22D1BWP30P140LVT U5625 ( .A1(i_data_bus[56]), .A2(n5395), .B1(
        i_data_bus[920]), .B2(n5389), .ZN(n5262) );
  AOI22D1BWP30P140LVT U5626 ( .A1(i_data_bus[984]), .A2(n5392), .B1(
        i_data_bus[88]), .B2(n5390), .ZN(n5261) );
  AOI22D1BWP30P140LVT U5627 ( .A1(i_data_bus[952]), .A2(n5397), .B1(
        i_data_bus[216]), .B2(n5400), .ZN(n5260) );
  ND4D1BWP30P140LVT U5628 ( .A1(n5263), .A2(n5262), .A3(n5261), .A4(n5260), 
        .ZN(n5277) );
  MOAI22D1BWP30P140LVT U5629 ( .A1(n5265), .A2(n5264), .B1(i_data_bus[728]), 
        .B2(n5424), .ZN(n5276) );
  AOI22D1BWP30P140LVT U5630 ( .A1(i_data_bus[792]), .A2(n5407), .B1(
        i_data_bus[824]), .B2(n5427), .ZN(n5269) );
  AOI22D1BWP30P140LVT U5631 ( .A1(i_data_bus[344]), .A2(n5422), .B1(
        i_data_bus[376]), .B2(n5423), .ZN(n5268) );
  AOI22D1BWP30P140LVT U5632 ( .A1(i_data_bus[632]), .A2(n5416), .B1(
        i_data_bus[536]), .B2(n5414), .ZN(n5267) );
  AOI22D1BWP30P140LVT U5633 ( .A1(i_data_bus[600]), .A2(n5415), .B1(
        i_data_bus[568]), .B2(n5417), .ZN(n5266) );
  ND4D1BWP30P140LVT U5634 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), 
        .ZN(n5275) );
  AOI22D1BWP30P140LVT U5635 ( .A1(i_data_bus[280]), .A2(n5394), .B1(
        i_data_bus[472]), .B2(n222), .ZN(n5273) );
  AOI22D1BWP30P140LVT U5636 ( .A1(i_data_bus[856]), .A2(n5425), .B1(
        i_data_bus[504]), .B2(n223), .ZN(n5272) );
  AOI22D1BWP30P140LVT U5637 ( .A1(i_data_bus[696]), .A2(n5393), .B1(
        i_data_bus[888]), .B2(n5410), .ZN(n5271) );
  AOI22D1BWP30P140LVT U5638 ( .A1(i_data_bus[440]), .A2(n5413), .B1(
        i_data_bus[760]), .B2(n5412), .ZN(n5270) );
  ND4D1BWP30P140LVT U5639 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), 
        .ZN(n5274) );
  NR4D0BWP30P140LVT U5640 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), 
        .ZN(n5278) );
  ND4D1BWP30P140LVT U5641 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), 
        .ZN(o_data_bus[24]) );
  AOI22D1BWP30P140LVT U5642 ( .A1(i_data_bus[121]), .A2(n5402), .B1(
        i_data_bus[249]), .B2(n5401), .ZN(n5302) );
  AOI22D1BWP30P140LVT U5643 ( .A1(i_data_bus[1017]), .A2(n5396), .B1(
        i_data_bus[89]), .B2(n5390), .ZN(n5301) );
  AOI22D1BWP30P140LVT U5644 ( .A1(i_data_bus[665]), .A2(n5426), .B1(
        i_data_bus[857]), .B2(n5425), .ZN(n5300) );
  AOI22D1BWP30P140LVT U5645 ( .A1(i_data_bus[25]), .A2(n5398), .B1(
        i_data_bus[153]), .B2(n5399), .ZN(n5285) );
  AOI22D1BWP30P140LVT U5646 ( .A1(i_data_bus[57]), .A2(n5395), .B1(
        i_data_bus[921]), .B2(n5389), .ZN(n5284) );
  AOI22D1BWP30P140LVT U5647 ( .A1(i_data_bus[953]), .A2(n5397), .B1(
        i_data_bus[185]), .B2(n5391), .ZN(n5283) );
  AOI22D1BWP30P140LVT U5648 ( .A1(i_data_bus[985]), .A2(n5392), .B1(
        i_data_bus[217]), .B2(n5400), .ZN(n5282) );
  ND4D1BWP30P140LVT U5649 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), 
        .ZN(n5298) );
  MOAI22D1BWP30P140LVT U5650 ( .A1(n5286), .A2(n5308), .B1(i_data_bus[729]), 
        .B2(n5424), .ZN(n5297) );
  AOI22D1BWP30P140LVT U5651 ( .A1(i_data_bus[345]), .A2(n5422), .B1(
        i_data_bus[761]), .B2(n5412), .ZN(n5290) );
  AOI22D1BWP30P140LVT U5652 ( .A1(i_data_bus[793]), .A2(n5407), .B1(
        i_data_bus[281]), .B2(n5394), .ZN(n5289) );
  AOI22D1BWP30P140LVT U5653 ( .A1(i_data_bus[569]), .A2(n5417), .B1(
        i_data_bus[601]), .B2(n5415), .ZN(n5288) );
  AOI22D1BWP30P140LVT U5654 ( .A1(i_data_bus[633]), .A2(n5416), .B1(
        i_data_bus[537]), .B2(n5414), .ZN(n5287) );
  ND4D1BWP30P140LVT U5655 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), 
        .ZN(n5296) );
  AOI22D1BWP30P140LVT U5656 ( .A1(i_data_bus[825]), .A2(n5427), .B1(
        i_data_bus[409]), .B2(n5411), .ZN(n5294) );
  AOI22D1BWP30P140LVT U5657 ( .A1(i_data_bus[377]), .A2(n5423), .B1(
        i_data_bus[473]), .B2(n222), .ZN(n5293) );
  AOI22D1BWP30P140LVT U5658 ( .A1(i_data_bus[313]), .A2(n5428), .B1(
        i_data_bus[441]), .B2(n5413), .ZN(n5292) );
  AOI22D1BWP30P140LVT U5659 ( .A1(i_data_bus[697]), .A2(n5393), .B1(
        i_data_bus[889]), .B2(n5410), .ZN(n5291) );
  ND4D1BWP30P140LVT U5660 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), 
        .ZN(n5295) );
  NR4D0BWP30P140LVT U5661 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), 
        .ZN(n5299) );
  ND4D1BWP30P140LVT U5662 ( .A1(n5302), .A2(n5301), .A3(n5300), .A4(n5299), 
        .ZN(o_data_bus[25]) );
  AOI22D1BWP30P140LVT U5663 ( .A1(i_data_bus[90]), .A2(n5390), .B1(
        i_data_bus[986]), .B2(n5392), .ZN(n5325) );
  AOI22D1BWP30P140LVT U5664 ( .A1(i_data_bus[1018]), .A2(n5396), .B1(
        i_data_bus[154]), .B2(n5399), .ZN(n5324) );
  AOI22D1BWP30P140LVT U5665 ( .A1(i_data_bus[442]), .A2(n5413), .B1(
        i_data_bus[698]), .B2(n5393), .ZN(n5323) );
  AOI22D1BWP30P140LVT U5666 ( .A1(i_data_bus[922]), .A2(n5389), .B1(
        i_data_bus[250]), .B2(n5401), .ZN(n5306) );
  AOI22D1BWP30P140LVT U5667 ( .A1(i_data_bus[954]), .A2(n5397), .B1(
        i_data_bus[186]), .B2(n5391), .ZN(n5305) );
  AOI22D1BWP30P140LVT U5668 ( .A1(i_data_bus[26]), .A2(n5398), .B1(
        i_data_bus[58]), .B2(n5395), .ZN(n5304) );
  AOI22D1BWP30P140LVT U5669 ( .A1(i_data_bus[122]), .A2(n5402), .B1(
        i_data_bus[218]), .B2(n5400), .ZN(n5303) );
  ND4D1BWP30P140LVT U5670 ( .A1(n5306), .A2(n5305), .A3(n5304), .A4(n5303), 
        .ZN(n5321) );
  OAI22D1BWP30P140LVT U5671 ( .A1(n5309), .A2(n5308), .B1(n5307), .B2(n228), 
        .ZN(n5320) );
  AOI22D1BWP30P140LVT U5672 ( .A1(i_data_bus[826]), .A2(n5427), .B1(
        i_data_bus[890]), .B2(n5410), .ZN(n5313) );
  AOI22D1BWP30P140LVT U5673 ( .A1(i_data_bus[346]), .A2(n5422), .B1(
        i_data_bus[762]), .B2(n5412), .ZN(n5312) );
  AOI22D1BWP30P140LVT U5674 ( .A1(i_data_bus[538]), .A2(n5414), .B1(
        i_data_bus[570]), .B2(n5417), .ZN(n5311) );
  AOI22D1BWP30P140LVT U5675 ( .A1(i_data_bus[602]), .A2(n5415), .B1(
        i_data_bus[634]), .B2(n5416), .ZN(n5310) );
  ND4D1BWP30P140LVT U5676 ( .A1(n5313), .A2(n5312), .A3(n5311), .A4(n5310), 
        .ZN(n5319) );
  AOI22D1BWP30P140LVT U5677 ( .A1(i_data_bus[858]), .A2(n5425), .B1(
        i_data_bus[730]), .B2(n5424), .ZN(n5317) );
  AOI22D1BWP30P140LVT U5678 ( .A1(i_data_bus[666]), .A2(n5426), .B1(
        i_data_bus[474]), .B2(n222), .ZN(n5316) );
  AOI22D1BWP30P140LVT U5679 ( .A1(i_data_bus[314]), .A2(n5428), .B1(
        i_data_bus[378]), .B2(n5423), .ZN(n5315) );
  AOI22D1BWP30P140LVT U5680 ( .A1(i_data_bus[282]), .A2(n5394), .B1(
        i_data_bus[794]), .B2(n5407), .ZN(n5314) );
  ND4D1BWP30P140LVT U5681 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), 
        .ZN(n5318) );
  NR4D0BWP30P140LVT U5682 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), 
        .ZN(n5322) );
  ND4D1BWP30P140LVT U5683 ( .A1(n5325), .A2(n5324), .A3(n5323), .A4(n5322), 
        .ZN(o_data_bus[26]) );
  AOI22D1BWP30P140LVT U5684 ( .A1(i_data_bus[60]), .A2(n5395), .B1(
        i_data_bus[220]), .B2(n5400), .ZN(n5346) );
  AOI22D1BWP30P140LVT U5685 ( .A1(i_data_bus[92]), .A2(n5390), .B1(
        i_data_bus[156]), .B2(n5399), .ZN(n5345) );
  AOI22D1BWP30P140LVT U5686 ( .A1(i_data_bus[508]), .A2(n223), .B1(
        i_data_bus[700]), .B2(n5393), .ZN(n5344) );
  AOI22D1BWP30P140LVT U5687 ( .A1(i_data_bus[956]), .A2(n5397), .B1(
        i_data_bus[1020]), .B2(n5396), .ZN(n5329) );
  AOI22D1BWP30P140LVT U5688 ( .A1(i_data_bus[988]), .A2(n5392), .B1(
        i_data_bus[252]), .B2(n5401), .ZN(n5328) );
  AOI22D1BWP30P140LVT U5689 ( .A1(i_data_bus[28]), .A2(n5398), .B1(
        i_data_bus[188]), .B2(n5391), .ZN(n5327) );
  AOI22D1BWP30P140LVT U5690 ( .A1(i_data_bus[924]), .A2(n5389), .B1(
        i_data_bus[124]), .B2(n5402), .ZN(n5326) );
  ND4D1BWP30P140LVT U5691 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), 
        .ZN(n5342) );
  MOAI22D1BWP30P140LVT U5692 ( .A1(n5330), .A2(n5351), .B1(i_data_bus[316]), 
        .B2(n5428), .ZN(n5341) );
  AOI22D1BWP30P140LVT U5693 ( .A1(i_data_bus[764]), .A2(n5412), .B1(
        i_data_bus[668]), .B2(n5426), .ZN(n5334) );
  AOI22D1BWP30P140LVT U5694 ( .A1(i_data_bus[348]), .A2(n5422), .B1(
        i_data_bus[380]), .B2(n5423), .ZN(n5333) );
  AOI22D1BWP30P140LVT U5695 ( .A1(i_data_bus[636]), .A2(n5416), .B1(
        i_data_bus[572]), .B2(n5417), .ZN(n5332) );
  AOI22D1BWP30P140LVT U5696 ( .A1(i_data_bus[540]), .A2(n5414), .B1(
        i_data_bus[604]), .B2(n5415), .ZN(n5331) );
  ND4D1BWP30P140LVT U5697 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), 
        .ZN(n5340) );
  AOI22D1BWP30P140LVT U5698 ( .A1(i_data_bus[828]), .A2(n5427), .B1(
        i_data_bus[860]), .B2(n5425), .ZN(n5338) );
  AOI22D1BWP30P140LVT U5699 ( .A1(i_data_bus[892]), .A2(n5410), .B1(
        i_data_bus[412]), .B2(n5411), .ZN(n5337) );
  AOI22D1BWP30P140LVT U5700 ( .A1(i_data_bus[796]), .A2(n5407), .B1(
        i_data_bus[732]), .B2(n5424), .ZN(n5336) );
  AOI22D1BWP30P140LVT U5701 ( .A1(i_data_bus[444]), .A2(n5413), .B1(
        i_data_bus[476]), .B2(n222), .ZN(n5335) );
  ND4D1BWP30P140LVT U5702 ( .A1(n5338), .A2(n5337), .A3(n5336), .A4(n5335), 
        .ZN(n5339) );
  NR4D0BWP30P140LVT U5703 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), 
        .ZN(n5343) );
  ND4D1BWP30P140LVT U5704 ( .A1(n5346), .A2(n5345), .A3(n5344), .A4(n5343), 
        .ZN(o_data_bus[28]) );
  AOI22D1BWP30P140LVT U5705 ( .A1(i_data_bus[29]), .A2(n5398), .B1(
        i_data_bus[93]), .B2(n5390), .ZN(n5368) );
  AOI22D1BWP30P140LVT U5706 ( .A1(i_data_bus[957]), .A2(n5397), .B1(
        i_data_bus[1021]), .B2(n5396), .ZN(n5367) );
  AOI22D1BWP30P140LVT U5707 ( .A1(i_data_bus[765]), .A2(n5412), .B1(
        i_data_bus[829]), .B2(n5427), .ZN(n5366) );
  AOI22D1BWP30P140LVT U5708 ( .A1(i_data_bus[61]), .A2(n5395), .B1(
        i_data_bus[157]), .B2(n5399), .ZN(n5350) );
  AOI22D1BWP30P140LVT U5709 ( .A1(i_data_bus[925]), .A2(n5389), .B1(
        i_data_bus[189]), .B2(n5391), .ZN(n5349) );
  AOI22D1BWP30P140LVT U5710 ( .A1(i_data_bus[989]), .A2(n5392), .B1(
        i_data_bus[253]), .B2(n5401), .ZN(n5348) );
  AOI22D1BWP30P140LVT U5711 ( .A1(i_data_bus[125]), .A2(n5402), .B1(
        i_data_bus[221]), .B2(n5400), .ZN(n5347) );
  ND4D1BWP30P140LVT U5712 ( .A1(n5350), .A2(n5349), .A3(n5348), .A4(n5347), 
        .ZN(n5364) );
  MOAI22D1BWP30P140LVT U5713 ( .A1(n5352), .A2(n5351), .B1(i_data_bus[733]), 
        .B2(n5424), .ZN(n5363) );
  AOI22D1BWP30P140LVT U5714 ( .A1(i_data_bus[349]), .A2(n5422), .B1(
        i_data_bus[477]), .B2(n222), .ZN(n5356) );
  AOI22D1BWP30P140LVT U5715 ( .A1(i_data_bus[509]), .A2(n223), .B1(
        i_data_bus[797]), .B2(n5407), .ZN(n5355) );
  AOI22D1BWP30P140LVT U5716 ( .A1(i_data_bus[637]), .A2(n5416), .B1(
        i_data_bus[541]), .B2(n5414), .ZN(n5354) );
  AOI22D1BWP30P140LVT U5717 ( .A1(i_data_bus[573]), .A2(n5417), .B1(
        i_data_bus[605]), .B2(n5415), .ZN(n5353) );
  ND4D1BWP30P140LVT U5718 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), 
        .ZN(n5362) );
  AOI22D1BWP30P140LVT U5719 ( .A1(i_data_bus[445]), .A2(n5413), .B1(
        i_data_bus[381]), .B2(n5423), .ZN(n5360) );
  AOI22D1BWP30P140LVT U5720 ( .A1(i_data_bus[669]), .A2(n5426), .B1(
        i_data_bus[317]), .B2(n5428), .ZN(n5359) );
  AOI22D1BWP30P140LVT U5721 ( .A1(i_data_bus[701]), .A2(n5393), .B1(
        i_data_bus[413]), .B2(n5411), .ZN(n5358) );
  AOI22D1BWP30P140LVT U5722 ( .A1(i_data_bus[861]), .A2(n5425), .B1(
        i_data_bus[893]), .B2(n5410), .ZN(n5357) );
  ND4D1BWP30P140LVT U5723 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), 
        .ZN(n5361) );
  NR4D0BWP30P140LVT U5724 ( .A1(n5364), .A2(n5363), .A3(n5362), .A4(n5361), 
        .ZN(n5365) );
  ND4D1BWP30P140LVT U5725 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), 
        .ZN(o_data_bus[29]) );
  AOI22D1BWP30P140LVT U5726 ( .A1(i_data_bus[62]), .A2(n5395), .B1(
        i_data_bus[190]), .B2(n5391), .ZN(n5388) );
  AOI22D1BWP30P140LVT U5727 ( .A1(i_data_bus[126]), .A2(n5402), .B1(
        i_data_bus[1022]), .B2(n5396), .ZN(n5387) );
  AOI22D1BWP30P140LVT U5728 ( .A1(i_data_bus[318]), .A2(n5428), .B1(
        i_data_bus[414]), .B2(n5411), .ZN(n5386) );
  AOI22D1BWP30P140LVT U5729 ( .A1(i_data_bus[446]), .A2(n5413), .B1(
        i_data_bus[702]), .B2(n5393), .ZN(n5384) );
  AOI22D1BWP30P140LVT U5730 ( .A1(i_data_bus[926]), .A2(n5389), .B1(
        i_data_bus[990]), .B2(n5392), .ZN(n5372) );
  AOI22D1BWP30P140LVT U5731 ( .A1(i_data_bus[30]), .A2(n5398), .B1(
        i_data_bus[94]), .B2(n5390), .ZN(n5371) );
  AOI22D1BWP30P140LVT U5732 ( .A1(i_data_bus[958]), .A2(n5397), .B1(
        i_data_bus[222]), .B2(n5400), .ZN(n5370) );
  AOI22D1BWP30P140LVT U5733 ( .A1(i_data_bus[254]), .A2(n5401), .B1(
        i_data_bus[158]), .B2(n5399), .ZN(n5369) );
  ND4D1BWP30P140LVT U5734 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), 
        .ZN(n5383) );
  AOI22D1BWP30P140LVT U5735 ( .A1(i_data_bus[350]), .A2(n5422), .B1(
        i_data_bus[766]), .B2(n5412), .ZN(n5376) );
  AOI22D1BWP30P140LVT U5736 ( .A1(i_data_bus[862]), .A2(n5425), .B1(
        i_data_bus[798]), .B2(n5407), .ZN(n5375) );
  AOI22D1BWP30P140LVT U5737 ( .A1(i_data_bus[574]), .A2(n5417), .B1(
        i_data_bus[606]), .B2(n5415), .ZN(n5374) );
  AOI22D1BWP30P140LVT U5738 ( .A1(i_data_bus[542]), .A2(n5414), .B1(
        i_data_bus[638]), .B2(n5416), .ZN(n5373) );
  ND4D1BWP30P140LVT U5739 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), 
        .ZN(n5382) );
  AOI22D1BWP30P140LVT U5740 ( .A1(i_data_bus[382]), .A2(n5423), .B1(
        i_data_bus[894]), .B2(n5410), .ZN(n5380) );
  AOI22D1BWP30P140LVT U5741 ( .A1(i_data_bus[670]), .A2(n5426), .B1(
        i_data_bus[510]), .B2(n223), .ZN(n5379) );
  AOI22D1BWP30P140LVT U5742 ( .A1(i_data_bus[830]), .A2(n5427), .B1(
        i_data_bus[734]), .B2(n5424), .ZN(n5378) );
  AOI22D1BWP30P140LVT U5743 ( .A1(i_data_bus[286]), .A2(n5394), .B1(
        i_data_bus[478]), .B2(n222), .ZN(n5377) );
  ND4D1BWP30P140LVT U5744 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), 
        .ZN(n5381) );
  INR4D0BWP30P140LVT U5745 ( .A1(n5384), .B1(n5383), .B2(n5382), .B3(n5381), 
        .ZN(n5385) );
  ND4D1BWP30P140LVT U5746 ( .A1(n5388), .A2(n5387), .A3(n5386), .A4(n5385), 
        .ZN(o_data_bus[30]) );
  AOI22D1BWP30P140LVT U5747 ( .A1(i_data_bus[95]), .A2(n5390), .B1(
        i_data_bus[927]), .B2(n5389), .ZN(n5440) );
  AOI22D1BWP30P140LVT U5748 ( .A1(i_data_bus[991]), .A2(n5392), .B1(
        i_data_bus[191]), .B2(n5391), .ZN(n5439) );
  AOI22D1BWP30P140LVT U5749 ( .A1(i_data_bus[287]), .A2(n5394), .B1(
        i_data_bus[703]), .B2(n5393), .ZN(n5438) );
  AOI22D1BWP30P140LVT U5750 ( .A1(i_data_bus[1023]), .A2(n5396), .B1(
        i_data_bus[63]), .B2(n5395), .ZN(n5406) );
  AOI22D1BWP30P140LVT U5751 ( .A1(i_data_bus[31]), .A2(n5398), .B1(
        i_data_bus[959]), .B2(n5397), .ZN(n5405) );
  AOI22D1BWP30P140LVT U5752 ( .A1(i_data_bus[223]), .A2(n5400), .B1(
        i_data_bus[159]), .B2(n5399), .ZN(n5404) );
  AOI22D1BWP30P140LVT U5753 ( .A1(i_data_bus[127]), .A2(n5402), .B1(
        i_data_bus[255]), .B2(n5401), .ZN(n5403) );
  ND4D1BWP30P140LVT U5754 ( .A1(n5406), .A2(n5405), .A3(n5404), .A4(n5403), 
        .ZN(n5436) );
  MOAI22D1BWP30P140LVT U5755 ( .A1(n5409), .A2(n5408), .B1(i_data_bus[799]), 
        .B2(n5407), .ZN(n5435) );
  AOI22D1BWP30P140LVT U5756 ( .A1(i_data_bus[415]), .A2(n5411), .B1(
        i_data_bus[895]), .B2(n5410), .ZN(n5421) );
  AOI22D1BWP30P140LVT U5757 ( .A1(i_data_bus[447]), .A2(n5413), .B1(
        i_data_bus[767]), .B2(n5412), .ZN(n5420) );
  AOI22D1BWP30P140LVT U5758 ( .A1(i_data_bus[607]), .A2(n5415), .B1(
        i_data_bus[543]), .B2(n5414), .ZN(n5419) );
  AOI22D1BWP30P140LVT U5759 ( .A1(i_data_bus[575]), .A2(n5417), .B1(
        i_data_bus[639]), .B2(n5416), .ZN(n5418) );
  ND4D1BWP30P140LVT U5760 ( .A1(n5421), .A2(n5420), .A3(n5419), .A4(n5418), 
        .ZN(n5434) );
  AOI22D1BWP30P140LVT U5761 ( .A1(i_data_bus[511]), .A2(n223), .B1(
        i_data_bus[351]), .B2(n5422), .ZN(n5432) );
  AOI22D1BWP30P140LVT U5762 ( .A1(i_data_bus[735]), .A2(n5424), .B1(
        i_data_bus[383]), .B2(n5423), .ZN(n5431) );
  AOI22D1BWP30P140LVT U5763 ( .A1(i_data_bus[671]), .A2(n5426), .B1(
        i_data_bus[863]), .B2(n5425), .ZN(n5430) );
  AOI22D1BWP30P140LVT U5764 ( .A1(i_data_bus[319]), .A2(n5428), .B1(
        i_data_bus[831]), .B2(n5427), .ZN(n5429) );
  ND4D1BWP30P140LVT U5765 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), 
        .ZN(n5433) );
  NR4D0BWP30P140LVT U5766 ( .A1(n5436), .A2(n5435), .A3(n5434), .A4(n5433), 
        .ZN(n5437) );
  ND4D1BWP30P140LVT U5767 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(n5437), 
        .ZN(o_data_bus[31]) );
  NR3D0P7BWP30P140LVT U5768 ( .A1(n5453), .A2(n5442), .A3(n5441), .ZN(n6157)
         );
  INVD1BWP30P140LVT U5769 ( .I(i_cmd[199]), .ZN(n5443) );
  NR3D0P7BWP30P140LVT U5770 ( .A1(n5444), .A2(n5443), .A3(n5460), .ZN(n5445)
         );
  AOI22D1BWP30P140LVT U5771 ( .A1(i_data_bus[32]), .A2(n6157), .B1(
        i_data_bus[768]), .B2(n6165), .ZN(n5509) );
  NR3D0P7BWP30P140LVT U5772 ( .A1(n5453), .A2(n5447), .A3(n5446), .ZN(n6162)
         );
  INR3D2BWP30P140LVT U5773 ( .A1(i_cmd[183]), .B1(n5448), .B2(n5462), .ZN(
        n6167) );
  AOI22D1BWP30P140LVT U5774 ( .A1(i_data_bus[96]), .A2(n6162), .B1(
        i_data_bus[704]), .B2(n6167), .ZN(n5508) );
  ND3D1BWP30P140LVT U5775 ( .A1(i_valid[11]), .A2(i_cmd[95]), .A3(n5468), .ZN(
        n6116) );
  ND3D1BWP30P140LVT U5776 ( .A1(i_valid[10]), .A2(i_cmd[87]), .A3(n5468), .ZN(
        n6094) );
  AOI22D1BWP30P140LVT U5777 ( .A1(i_data_bus[352]), .A2(n6188), .B1(
        i_data_bus[320]), .B2(n6178), .ZN(n5507) );
  NR3D0P7BWP30P140LVT U5778 ( .A1(n5453), .A2(n5450), .A3(n5449), .ZN(n6169)
         );
  NR3D0P7BWP30P140LVT U5779 ( .A1(n5453), .A2(n5452), .A3(n5451), .ZN(n6163)
         );
  AOI22D1BWP30P140LVT U5780 ( .A1(i_data_bus[0]), .A2(n6169), .B1(
        i_data_bus[64]), .B2(n6163), .ZN(n5467) );
  INVD1BWP30P140LVT U5781 ( .I(i_cmd[167]), .ZN(n5454) );
  NR3D0P7BWP30P140LVT U5782 ( .A1(n5455), .A2(n5454), .A3(n5462), .ZN(n5456)
         );
  INR3D2BWP30P140LVT U5783 ( .A1(i_cmd[223]), .B1(n5457), .B2(n5460), .ZN(
        n6168) );
  AOI22D1BWP30P140LVT U5784 ( .A1(i_data_bus[640]), .A2(n6156), .B1(
        i_data_bus[864]), .B2(n6168), .ZN(n5466) );
  INR3D2BWP30P140LVT U5785 ( .A1(i_cmd[191]), .B1(n5458), .B2(n5462), .ZN(
        n6159) );
  INR3D2BWP30P140LVT U5786 ( .A1(i_cmd[207]), .B1(n5459), .B2(n5460), .ZN(
        n6166) );
  AOI22D1BWP30P140LVT U5787 ( .A1(i_data_bus[736]), .A2(n6159), .B1(
        i_data_bus[800]), .B2(n6166), .ZN(n5465) );
  INR3D2BWP30P140LVT U5788 ( .A1(i_cmd[215]), .B1(n5461), .B2(n5460), .ZN(
        n6164) );
  INR3D2BWP30P140LVT U5789 ( .A1(i_cmd[175]), .B1(n5463), .B2(n5462), .ZN(
        n6158) );
  AOI22D1BWP30P140LVT U5790 ( .A1(i_data_bus[832]), .A2(n6164), .B1(
        i_data_bus[672]), .B2(n6158), .ZN(n5464) );
  ND4D1BWP30P140LVT U5791 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), 
        .ZN(n5505) );
  ND3D1BWP30P140LVT U5792 ( .A1(i_valid[15]), .A2(i_cmd[127]), .A3(n5492), 
        .ZN(n5898) );
  ND3D1BWP30P140LVT U5793 ( .A1(i_valid[9]), .A2(i_cmd[79]), .A3(n5468), .ZN(
        n5920) );
  MOAI22D1BWP30P140LVT U5794 ( .A1(n5469), .A2(n5898), .B1(i_data_bus[288]), 
        .B2(n6193), .ZN(n5504) );
  INR3D2BWP30P140LVT U5795 ( .A1(i_cmd[255]), .B1(n5470), .B2(n5489), .ZN(
        n6177) );
  AOI22D1BWP30P140LVT U5796 ( .A1(i_data_bus[992]), .A2(n6177), .B1(
        i_data_bus[224]), .B2(n6160), .ZN(n5485) );
  INVD1BWP30P140LVT U5797 ( .I(i_cmd[231]), .ZN(n5472) );
  AOI22D1BWP30P140LVT U5798 ( .A1(i_data_bus[896]), .A2(n5474), .B1(
        i_data_bus[384]), .B2(n6192), .ZN(n5484) );
  INR3D2BWP30P140LVT U5799 ( .A1(i_cmd[159]), .B1(n5478), .B2(n5480), .ZN(
        n6182) );
  AOI22D1BWP30P140LVT U5800 ( .A1(i_data_bus[512]), .A2(n6181), .B1(
        i_data_bus[608]), .B2(n6182), .ZN(n5483) );
  INR3D2BWP30P140LVT U5801 ( .A1(i_cmd[143]), .B1(n5479), .B2(n5480), .ZN(
        n6180) );
  INR3D2BWP30P140LVT U5802 ( .A1(i_cmd[151]), .B1(n5481), .B2(n5480), .ZN(
        n6179) );
  AOI22D1BWP30P140LVT U5803 ( .A1(i_data_bus[544]), .A2(n6180), .B1(
        i_data_bus[576]), .B2(n6179), .ZN(n5482) );
  ND4D1BWP30P140LVT U5804 ( .A1(n5485), .A2(n5484), .A3(n5483), .A4(n5482), 
        .ZN(n5503) );
  INR3D2BWP30P140LVT U5805 ( .A1(i_cmd[239]), .B1(n5486), .B2(n5489), .ZN(
        n6191) );
  AOI22D1BWP30P140LVT U5806 ( .A1(i_data_bus[928]), .A2(n6191), .B1(
        i_data_bus[160]), .B2(n5488), .ZN(n5501) );
  INR3D2BWP30P140LVT U5807 ( .A1(i_cmd[247]), .B1(n5490), .B2(n5489), .ZN(
        n6161) );
  ND3D1BWP30P140LVT U5808 ( .A1(i_valid[13]), .A2(i_cmd[111]), .A3(n5492), 
        .ZN(n5986) );
  INVD1BWP30P140LVT U5809 ( .I(n5986), .ZN(n5491) );
  AOI22D1BWP30P140LVT U5810 ( .A1(i_data_bus[960]), .A2(n6161), .B1(
        i_data_bus[416]), .B2(n5491), .ZN(n5500) );
  ND3D1BWP30P140LVT U5811 ( .A1(i_valid[14]), .A2(i_cmd[119]), .A3(n5492), 
        .ZN(n5728) );
  AOI22D1BWP30P140LVT U5812 ( .A1(i_data_bus[448]), .A2(n6187), .B1(
        i_data_bus[128]), .B2(n6190), .ZN(n5499) );
  AOI22D1BWP30P140LVT U5813 ( .A1(i_data_bus[192]), .A2(n6189), .B1(
        i_data_bus[256]), .B2(n6143), .ZN(n5498) );
  ND4D1BWP30P140LVT U5814 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), 
        .ZN(n5502) );
  NR4D0BWP30P140LVT U5815 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), 
        .ZN(n5506) );
  ND4D1BWP30P140LVT U5816 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), 
        .ZN(o_data_bus[224]) );
  AOI22D1BWP30P140LVT U5817 ( .A1(i_data_bus[865]), .A2(n6168), .B1(
        i_data_bus[833]), .B2(n6164), .ZN(n5530) );
  AOI22D1BWP30P140LVT U5818 ( .A1(i_data_bus[1]), .A2(n6169), .B1(
        i_data_bus[641]), .B2(n6156), .ZN(n5529) );
  AOI22D1BWP30P140LVT U5819 ( .A1(i_data_bus[897]), .A2(n5474), .B1(
        i_data_bus[321]), .B2(n6178), .ZN(n5528) );
  AOI22D1BWP30P140LVT U5820 ( .A1(i_data_bus[33]), .A2(n6157), .B1(
        i_data_bus[705]), .B2(n6167), .ZN(n5513) );
  AOI22D1BWP30P140LVT U5821 ( .A1(i_data_bus[97]), .A2(n6162), .B1(
        i_data_bus[673]), .B2(n6158), .ZN(n5512) );
  AOI22D1BWP30P140LVT U5822 ( .A1(i_data_bus[65]), .A2(n6163), .B1(
        i_data_bus[769]), .B2(n6165), .ZN(n5511) );
  AOI22D1BWP30P140LVT U5823 ( .A1(i_data_bus[801]), .A2(n6166), .B1(
        i_data_bus[737]), .B2(n6159), .ZN(n5510) );
  ND4D1BWP30P140LVT U5824 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5510), 
        .ZN(n5526) );
  MOAI22D1BWP30P140LVT U5825 ( .A1(n5514), .A2(n5898), .B1(i_data_bus[193]), 
        .B2(n6189), .ZN(n5525) );
  AOI22D1BWP30P140LVT U5826 ( .A1(i_data_bus[961]), .A2(n6161), .B1(
        i_data_bus[385]), .B2(n6192), .ZN(n5518) );
  AOI22D1BWP30P140LVT U5827 ( .A1(i_data_bus[353]), .A2(n6188), .B1(
        i_data_bus[289]), .B2(n6193), .ZN(n5517) );
  AOI22D1BWP30P140LVT U5828 ( .A1(i_data_bus[545]), .A2(n6180), .B1(
        i_data_bus[513]), .B2(n6181), .ZN(n5516) );
  AOI22D1BWP30P140LVT U5829 ( .A1(i_data_bus[577]), .A2(n6179), .B1(
        i_data_bus[609]), .B2(n6182), .ZN(n5515) );
  ND4D1BWP30P140LVT U5830 ( .A1(n5518), .A2(n5517), .A3(n5516), .A4(n5515), 
        .ZN(n5524) );
  AOI22D1BWP30P140LVT U5831 ( .A1(i_data_bus[993]), .A2(n6177), .B1(
        i_data_bus[225]), .B2(n6160), .ZN(n5522) );
  AOI22D1BWP30P140LVT U5832 ( .A1(i_data_bus[161]), .A2(n5488), .B1(
        i_data_bus[417]), .B2(n5491), .ZN(n5521) );
  AOI22D1BWP30P140LVT U5833 ( .A1(i_data_bus[929]), .A2(n6191), .B1(
        i_data_bus[449]), .B2(n6187), .ZN(n5520) );
  AOI22D1BWP30P140LVT U5834 ( .A1(i_data_bus[257]), .A2(n6143), .B1(
        i_data_bus[129]), .B2(n6190), .ZN(n5519) );
  ND4D1BWP30P140LVT U5835 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), 
        .ZN(n5523) );
  NR4D0BWP30P140LVT U5836 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), 
        .ZN(n5527) );
  ND4D1BWP30P140LVT U5837 ( .A1(n5530), .A2(n5529), .A3(n5528), .A4(n5527), 
        .ZN(o_data_bus[225]) );
  AOI22D1BWP30P140LVT U5838 ( .A1(i_data_bus[66]), .A2(n6163), .B1(
        i_data_bus[34]), .B2(n6157), .ZN(n5552) );
  AOI22D1BWP30P140LVT U5839 ( .A1(i_data_bus[770]), .A2(n6165), .B1(
        i_data_bus[706]), .B2(n6167), .ZN(n5551) );
  AOI22D1BWP30P140LVT U5840 ( .A1(i_data_bus[386]), .A2(n6192), .B1(
        i_data_bus[130]), .B2(n6190), .ZN(n5550) );
  AOI22D1BWP30P140LVT U5841 ( .A1(i_data_bus[802]), .A2(n6166), .B1(
        i_data_bus[738]), .B2(n6159), .ZN(n5534) );
  AOI22D1BWP30P140LVT U5842 ( .A1(i_data_bus[98]), .A2(n6162), .B1(
        i_data_bus[642]), .B2(n6156), .ZN(n5533) );
  AOI22D1BWP30P140LVT U5843 ( .A1(i_data_bus[2]), .A2(n6169), .B1(
        i_data_bus[834]), .B2(n6164), .ZN(n5532) );
  AOI22D1BWP30P140LVT U5844 ( .A1(i_data_bus[866]), .A2(n6168), .B1(
        i_data_bus[674]), .B2(n6158), .ZN(n5531) );
  ND4D1BWP30P140LVT U5845 ( .A1(n5534), .A2(n5533), .A3(n5532), .A4(n5531), 
        .ZN(n5548) );
  INVD1BWP30P140LVT U5846 ( .I(n6189), .ZN(n5963) );
  OAI22D1BWP30P140LVT U5847 ( .A1(n5536), .A2(n5963), .B1(n5535), .B2(n120), 
        .ZN(n5547) );
  AOI22D1BWP30P140LVT U5848 ( .A1(i_data_bus[962]), .A2(n6161), .B1(
        i_data_bus[322]), .B2(n6178), .ZN(n5540) );
  AOI22D1BWP30P140LVT U5849 ( .A1(i_data_bus[290]), .A2(n6193), .B1(
        i_data_bus[482]), .B2(n6174), .ZN(n5539) );
  AOI22D1BWP30P140LVT U5850 ( .A1(i_data_bus[578]), .A2(n6179), .B1(
        i_data_bus[610]), .B2(n6182), .ZN(n5538) );
  AOI22D1BWP30P140LVT U5851 ( .A1(i_data_bus[546]), .A2(n6180), .B1(
        i_data_bus[514]), .B2(n6181), .ZN(n5537) );
  ND4D1BWP30P140LVT U5852 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), 
        .ZN(n5546) );
  AOI22D1BWP30P140LVT U5853 ( .A1(i_data_bus[930]), .A2(n6191), .B1(
        i_data_bus[418]), .B2(n5491), .ZN(n5544) );
  AOI22D1BWP30P140LVT U5854 ( .A1(i_data_bus[898]), .A2(n5474), .B1(
        i_data_bus[450]), .B2(n6187), .ZN(n5543) );
  AOI22D1BWP30P140LVT U5855 ( .A1(i_data_bus[994]), .A2(n6177), .B1(
        i_data_bus[354]), .B2(n6188), .ZN(n5542) );
  AOI22D1BWP30P140LVT U5856 ( .A1(i_data_bus[162]), .A2(n5488), .B1(
        i_data_bus[226]), .B2(n6160), .ZN(n5541) );
  ND4D1BWP30P140LVT U5857 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), 
        .ZN(n5545) );
  NR4D0BWP30P140LVT U5858 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), 
        .ZN(n5549) );
  ND4D1BWP30P140LVT U5859 ( .A1(n5552), .A2(n5551), .A3(n5550), .A4(n5549), 
        .ZN(o_data_bus[226]) );
  AOI22D1BWP30P140LVT U5860 ( .A1(i_data_bus[771]), .A2(n6165), .B1(
        i_data_bus[739]), .B2(n6159), .ZN(n5574) );
  AOI22D1BWP30P140LVT U5861 ( .A1(i_data_bus[67]), .A2(n6163), .B1(
        i_data_bus[35]), .B2(n6157), .ZN(n5573) );
  AOI22D1BWP30P140LVT U5862 ( .A1(i_data_bus[963]), .A2(n6161), .B1(
        i_data_bus[195]), .B2(n6189), .ZN(n5572) );
  AOI22D1BWP30P140LVT U5863 ( .A1(i_data_bus[3]), .A2(n6169), .B1(
        i_data_bus[803]), .B2(n6166), .ZN(n5556) );
  AOI22D1BWP30P140LVT U5864 ( .A1(i_data_bus[99]), .A2(n6162), .B1(
        i_data_bus[707]), .B2(n6167), .ZN(n5555) );
  AOI22D1BWP30P140LVT U5865 ( .A1(i_data_bus[835]), .A2(n6164), .B1(
        i_data_bus[867]), .B2(n6168), .ZN(n5554) );
  AOI22D1BWP30P140LVT U5866 ( .A1(i_data_bus[675]), .A2(n6158), .B1(
        i_data_bus[643]), .B2(n6156), .ZN(n5553) );
  ND4D1BWP30P140LVT U5867 ( .A1(n5556), .A2(n5555), .A3(n5554), .A4(n5553), 
        .ZN(n5570) );
  INVD1BWP30P140LVT U5868 ( .I(n6190), .ZN(n5876) );
  OAI22D1BWP30P140LVT U5869 ( .A1(n5558), .A2(n5986), .B1(n5557), .B2(n5876), 
        .ZN(n5569) );
  AOI22D1BWP30P140LVT U5870 ( .A1(i_data_bus[355]), .A2(n6188), .B1(
        i_data_bus[227]), .B2(n6160), .ZN(n5562) );
  AOI22D1BWP30P140LVT U5871 ( .A1(i_data_bus[995]), .A2(n6177), .B1(
        i_data_bus[323]), .B2(n6178), .ZN(n5561) );
  AOI22D1BWP30P140LVT U5872 ( .A1(i_data_bus[515]), .A2(n6181), .B1(
        i_data_bus[579]), .B2(n6179), .ZN(n5560) );
  AOI22D1BWP30P140LVT U5873 ( .A1(i_data_bus[547]), .A2(n6180), .B1(
        i_data_bus[611]), .B2(n6182), .ZN(n5559) );
  ND4D1BWP30P140LVT U5874 ( .A1(n5562), .A2(n5561), .A3(n5560), .A4(n5559), 
        .ZN(n5568) );
  AOI22D1BWP30P140LVT U5875 ( .A1(i_data_bus[899]), .A2(n5474), .B1(
        i_data_bus[483]), .B2(n6174), .ZN(n5566) );
  AOI22D1BWP30P140LVT U5876 ( .A1(i_data_bus[163]), .A2(n5488), .B1(
        i_data_bus[451]), .B2(n6187), .ZN(n5565) );
  AOI22D1BWP30P140LVT U5877 ( .A1(i_data_bus[387]), .A2(n6192), .B1(
        i_data_bus[291]), .B2(n6193), .ZN(n5564) );
  AOI22D1BWP30P140LVT U5878 ( .A1(i_data_bus[931]), .A2(n6191), .B1(
        i_data_bus[259]), .B2(n6143), .ZN(n5563) );
  ND4D1BWP30P140LVT U5879 ( .A1(n5566), .A2(n5565), .A3(n5564), .A4(n5563), 
        .ZN(n5567) );
  NR4D0BWP30P140LVT U5880 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), 
        .ZN(n5571) );
  ND4D1BWP30P140LVT U5881 ( .A1(n5574), .A2(n5573), .A3(n5572), .A4(n5571), 
        .ZN(o_data_bus[227]) );
  AOI22D1BWP30P140LVT U5882 ( .A1(i_data_bus[4]), .A2(n6169), .B1(
        i_data_bus[836]), .B2(n6164), .ZN(n5595) );
  AOI22D1BWP30P140LVT U5883 ( .A1(i_data_bus[740]), .A2(n6159), .B1(
        i_data_bus[868]), .B2(n6168), .ZN(n5594) );
  AOI22D1BWP30P140LVT U5884 ( .A1(i_data_bus[932]), .A2(n6191), .B1(
        i_data_bus[324]), .B2(n6178), .ZN(n5593) );
  AOI22D1BWP30P140LVT U5885 ( .A1(i_data_bus[708]), .A2(n6167), .B1(
        i_data_bus[676]), .B2(n6158), .ZN(n5578) );
  AOI22D1BWP30P140LVT U5886 ( .A1(i_data_bus[772]), .A2(n6165), .B1(
        i_data_bus[804]), .B2(n6166), .ZN(n5577) );
  AOI22D1BWP30P140LVT U5887 ( .A1(i_data_bus[68]), .A2(n6163), .B1(
        i_data_bus[36]), .B2(n6157), .ZN(n5576) );
  AOI22D1BWP30P140LVT U5888 ( .A1(i_data_bus[100]), .A2(n6162), .B1(
        i_data_bus[644]), .B2(n6156), .ZN(n5575) );
  ND4D1BWP30P140LVT U5889 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), 
        .ZN(n5591) );
  MOAI22D1BWP30P140LVT U5890 ( .A1(n5579), .A2(n5728), .B1(i_data_bus[196]), 
        .B2(n6189), .ZN(n5590) );
  AOI22D1BWP30P140LVT U5891 ( .A1(i_data_bus[228]), .A2(n6160), .B1(
        i_data_bus[164]), .B2(n5488), .ZN(n5583) );
  AOI22D1BWP30P140LVT U5892 ( .A1(i_data_bus[996]), .A2(n6177), .B1(
        i_data_bus[484]), .B2(n6174), .ZN(n5582) );
  AOI22D1BWP30P140LVT U5893 ( .A1(i_data_bus[548]), .A2(n6180), .B1(
        i_data_bus[580]), .B2(n6179), .ZN(n5581) );
  AOI22D1BWP30P140LVT U5894 ( .A1(i_data_bus[612]), .A2(n6182), .B1(
        i_data_bus[516]), .B2(n6181), .ZN(n5580) );
  ND4D1BWP30P140LVT U5895 ( .A1(n5583), .A2(n5582), .A3(n5581), .A4(n5580), 
        .ZN(n5589) );
  AOI22D1BWP30P140LVT U5896 ( .A1(i_data_bus[964]), .A2(n6161), .B1(
        i_data_bus[356]), .B2(n6188), .ZN(n5587) );
  AOI22D1BWP30P140LVT U5897 ( .A1(i_data_bus[900]), .A2(n5474), .B1(
        i_data_bus[420]), .B2(n5491), .ZN(n5586) );
  AOI22D1BWP30P140LVT U5898 ( .A1(i_data_bus[292]), .A2(n6193), .B1(
        i_data_bus[388]), .B2(n6192), .ZN(n5585) );
  AOI22D1BWP30P140LVT U5899 ( .A1(i_data_bus[132]), .A2(n6190), .B1(
        i_data_bus[260]), .B2(n6143), .ZN(n5584) );
  ND4D1BWP30P140LVT U5900 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), 
        .ZN(n5588) );
  NR4D0BWP30P140LVT U5901 ( .A1(n5591), .A2(n5590), .A3(n5589), .A4(n5588), 
        .ZN(n5592) );
  ND4D1BWP30P140LVT U5902 ( .A1(n5595), .A2(n5594), .A3(n5593), .A4(n5592), 
        .ZN(o_data_bus[228]) );
  AOI22D1BWP30P140LVT U5903 ( .A1(i_data_bus[37]), .A2(n6157), .B1(
        i_data_bus[645]), .B2(n6156), .ZN(n5616) );
  AOI22D1BWP30P140LVT U5904 ( .A1(i_data_bus[69]), .A2(n6163), .B1(
        i_data_bus[805]), .B2(n6166), .ZN(n5615) );
  AOI22D1BWP30P140LVT U5905 ( .A1(i_data_bus[165]), .A2(n5488), .B1(
        i_data_bus[389]), .B2(n6192), .ZN(n5614) );
  AOI22D1BWP30P140LVT U5906 ( .A1(i_data_bus[101]), .A2(n6162), .B1(
        i_data_bus[677]), .B2(n6158), .ZN(n5599) );
  AOI22D1BWP30P140LVT U5907 ( .A1(i_data_bus[837]), .A2(n6164), .B1(
        i_data_bus[869]), .B2(n6168), .ZN(n5598) );
  AOI22D1BWP30P140LVT U5908 ( .A1(i_data_bus[5]), .A2(n6169), .B1(
        i_data_bus[773]), .B2(n6165), .ZN(n5597) );
  AOI22D1BWP30P140LVT U5909 ( .A1(i_data_bus[709]), .A2(n6167), .B1(
        i_data_bus[741]), .B2(n6159), .ZN(n5596) );
  ND4D1BWP30P140LVT U5910 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), 
        .ZN(n5612) );
  MOAI22D1BWP30P140LVT U5911 ( .A1(n5600), .A2(n5920), .B1(i_data_bus[453]), 
        .B2(n6187), .ZN(n5611) );
  AOI22D1BWP30P140LVT U5912 ( .A1(i_data_bus[933]), .A2(n6191), .B1(
        i_data_bus[261]), .B2(n6143), .ZN(n5604) );
  AOI22D1BWP30P140LVT U5913 ( .A1(i_data_bus[901]), .A2(n5474), .B1(
        i_data_bus[197]), .B2(n6189), .ZN(n5603) );
  AOI22D1BWP30P140LVT U5914 ( .A1(i_data_bus[581]), .A2(n6179), .B1(
        i_data_bus[613]), .B2(n6182), .ZN(n5602) );
  AOI22D1BWP30P140LVT U5915 ( .A1(i_data_bus[517]), .A2(n6181), .B1(
        i_data_bus[549]), .B2(n6180), .ZN(n5601) );
  ND4D1BWP30P140LVT U5916 ( .A1(n5604), .A2(n5603), .A3(n5602), .A4(n5601), 
        .ZN(n5610) );
  AOI22D1BWP30P140LVT U5917 ( .A1(i_data_bus[965]), .A2(n6161), .B1(
        i_data_bus[485]), .B2(n6174), .ZN(n5608) );
  AOI22D1BWP30P140LVT U5918 ( .A1(i_data_bus[997]), .A2(n6177), .B1(
        i_data_bus[325]), .B2(n6178), .ZN(n5607) );
  AOI22D1BWP30P140LVT U5919 ( .A1(i_data_bus[133]), .A2(n6190), .B1(
        i_data_bus[229]), .B2(n6160), .ZN(n5606) );
  AOI22D1BWP30P140LVT U5920 ( .A1(i_data_bus[357]), .A2(n6188), .B1(
        i_data_bus[421]), .B2(n5491), .ZN(n5605) );
  ND4D1BWP30P140LVT U5921 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), 
        .ZN(n5609) );
  NR4D0BWP30P140LVT U5922 ( .A1(n5612), .A2(n5611), .A3(n5610), .A4(n5609), 
        .ZN(n5613) );
  ND4D1BWP30P140LVT U5923 ( .A1(n5616), .A2(n5615), .A3(n5614), .A4(n5613), 
        .ZN(o_data_bus[229]) );
  AOI22D1BWP30P140LVT U5924 ( .A1(i_data_bus[742]), .A2(n6159), .B1(
        i_data_bus[710]), .B2(n6167), .ZN(n5637) );
  AOI22D1BWP30P140LVT U5925 ( .A1(i_data_bus[6]), .A2(n6169), .B1(
        i_data_bus[678]), .B2(n6158), .ZN(n5636) );
  AOI22D1BWP30P140LVT U5926 ( .A1(i_data_bus[934]), .A2(n6191), .B1(
        i_data_bus[390]), .B2(n6192), .ZN(n5635) );
  AOI22D1BWP30P140LVT U5927 ( .A1(i_data_bus[70]), .A2(n6163), .B1(
        i_data_bus[870]), .B2(n6168), .ZN(n5620) );
  AOI22D1BWP30P140LVT U5928 ( .A1(i_data_bus[38]), .A2(n6157), .B1(
        i_data_bus[838]), .B2(n6164), .ZN(n5619) );
  AOI22D1BWP30P140LVT U5929 ( .A1(i_data_bus[806]), .A2(n6166), .B1(
        i_data_bus[646]), .B2(n6156), .ZN(n5618) );
  AOI22D1BWP30P140LVT U5930 ( .A1(i_data_bus[102]), .A2(n6162), .B1(
        i_data_bus[774]), .B2(n6165), .ZN(n5617) );
  ND4D1BWP30P140LVT U5931 ( .A1(n5620), .A2(n5619), .A3(n5618), .A4(n5617), 
        .ZN(n5633) );
  MOAI22D1BWP30P140LVT U5932 ( .A1(n5621), .A2(n5728), .B1(i_data_bus[262]), 
        .B2(n6143), .ZN(n5632) );
  AOI22D1BWP30P140LVT U5933 ( .A1(i_data_bus[230]), .A2(n6160), .B1(
        i_data_bus[358]), .B2(n6188), .ZN(n5625) );
  AOI22D1BWP30P140LVT U5934 ( .A1(i_data_bus[486]), .A2(n6174), .B1(
        i_data_bus[134]), .B2(n6190), .ZN(n5624) );
  AOI22D1BWP30P140LVT U5935 ( .A1(i_data_bus[582]), .A2(n6179), .B1(
        i_data_bus[550]), .B2(n6180), .ZN(n5623) );
  AOI22D1BWP30P140LVT U5936 ( .A1(i_data_bus[614]), .A2(n6182), .B1(
        i_data_bus[518]), .B2(n6181), .ZN(n5622) );
  ND4D1BWP30P140LVT U5937 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), 
        .ZN(n5631) );
  AOI22D1BWP30P140LVT U5938 ( .A1(i_data_bus[902]), .A2(n5474), .B1(
        i_data_bus[326]), .B2(n6178), .ZN(n5629) );
  AOI22D1BWP30P140LVT U5939 ( .A1(i_data_bus[998]), .A2(n6177), .B1(
        i_data_bus[198]), .B2(n6189), .ZN(n5628) );
  AOI22D1BWP30P140LVT U5940 ( .A1(i_data_bus[166]), .A2(n5488), .B1(
        i_data_bus[422]), .B2(n5491), .ZN(n5627) );
  AOI22D1BWP30P140LVT U5941 ( .A1(i_data_bus[966]), .A2(n6161), .B1(
        i_data_bus[294]), .B2(n6193), .ZN(n5626) );
  ND4D1BWP30P140LVT U5942 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), 
        .ZN(n5630) );
  NR4D0BWP30P140LVT U5943 ( .A1(n5633), .A2(n5632), .A3(n5631), .A4(n5630), 
        .ZN(n5634) );
  ND4D1BWP30P140LVT U5944 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), 
        .ZN(o_data_bus[230]) );
  AOI22D1BWP30P140LVT U5945 ( .A1(i_data_bus[839]), .A2(n6164), .B1(
        i_data_bus[647]), .B2(n6156), .ZN(n5658) );
  AOI22D1BWP30P140LVT U5946 ( .A1(i_data_bus[103]), .A2(n6162), .B1(
        i_data_bus[743]), .B2(n6159), .ZN(n5657) );
  AOI22D1BWP30P140LVT U5947 ( .A1(i_data_bus[967]), .A2(n6161), .B1(
        i_data_bus[295]), .B2(n6193), .ZN(n5656) );
  AOI22D1BWP30P140LVT U5948 ( .A1(i_data_bus[39]), .A2(n6157), .B1(
        i_data_bus[7]), .B2(n6169), .ZN(n5641) );
  AOI22D1BWP30P140LVT U5949 ( .A1(i_data_bus[807]), .A2(n6166), .B1(
        i_data_bus[711]), .B2(n6167), .ZN(n5640) );
  AOI22D1BWP30P140LVT U5950 ( .A1(i_data_bus[71]), .A2(n6163), .B1(
        i_data_bus[871]), .B2(n6168), .ZN(n5639) );
  AOI22D1BWP30P140LVT U5951 ( .A1(i_data_bus[679]), .A2(n6158), .B1(
        i_data_bus[775]), .B2(n6165), .ZN(n5638) );
  ND4D1BWP30P140LVT U5952 ( .A1(n5641), .A2(n5640), .A3(n5639), .A4(n5638), 
        .ZN(n5654) );
  MOAI22D1BWP30P140LVT U5953 ( .A1(n5642), .A2(n5963), .B1(i_data_bus[391]), 
        .B2(n6192), .ZN(n5653) );
  AOI22D1BWP30P140LVT U5954 ( .A1(i_data_bus[935]), .A2(n6191), .B1(
        i_data_bus[487]), .B2(n6174), .ZN(n5646) );
  AOI22D1BWP30P140LVT U5955 ( .A1(i_data_bus[455]), .A2(n6187), .B1(
        i_data_bus[327]), .B2(n6178), .ZN(n5645) );
  AOI22D1BWP30P140LVT U5956 ( .A1(i_data_bus[519]), .A2(n6181), .B1(
        i_data_bus[583]), .B2(n6179), .ZN(n5644) );
  AOI22D1BWP30P140LVT U5957 ( .A1(i_data_bus[615]), .A2(n6182), .B1(
        i_data_bus[551]), .B2(n6180), .ZN(n5643) );
  ND4D1BWP30P140LVT U5958 ( .A1(n5646), .A2(n5645), .A3(n5644), .A4(n5643), 
        .ZN(n5652) );
  AOI22D1BWP30P140LVT U5959 ( .A1(i_data_bus[263]), .A2(n6143), .B1(
        i_data_bus[135]), .B2(n6190), .ZN(n5650) );
  AOI22D1BWP30P140LVT U5960 ( .A1(i_data_bus[359]), .A2(n6188), .B1(
        i_data_bus[231]), .B2(n6160), .ZN(n5649) );
  AOI22D1BWP30P140LVT U5961 ( .A1(i_data_bus[903]), .A2(n5474), .B1(
        i_data_bus[999]), .B2(n6177), .ZN(n5648) );
  AOI22D1BWP30P140LVT U5962 ( .A1(i_data_bus[167]), .A2(n5488), .B1(
        i_data_bus[423]), .B2(n5491), .ZN(n5647) );
  ND4D1BWP30P140LVT U5963 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), 
        .ZN(n5651) );
  NR4D0BWP30P140LVT U5964 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), 
        .ZN(n5655) );
  ND4D1BWP30P140LVT U5965 ( .A1(n5658), .A2(n5657), .A3(n5656), .A4(n5655), 
        .ZN(o_data_bus[231]) );
  AOI22D1BWP30P140LVT U5966 ( .A1(i_data_bus[744]), .A2(n6159), .B1(
        i_data_bus[680]), .B2(n6158), .ZN(n5679) );
  AOI22D1BWP30P140LVT U5967 ( .A1(i_data_bus[104]), .A2(n6162), .B1(
        i_data_bus[72]), .B2(n6163), .ZN(n5678) );
  AOI22D1BWP30P140LVT U5968 ( .A1(i_data_bus[200]), .A2(n6189), .B1(
        i_data_bus[136]), .B2(n6190), .ZN(n5677) );
  AOI22D1BWP30P140LVT U5969 ( .A1(i_data_bus[808]), .A2(n6166), .B1(
        i_data_bus[776]), .B2(n6165), .ZN(n5662) );
  AOI22D1BWP30P140LVT U5970 ( .A1(i_data_bus[8]), .A2(n6169), .B1(
        i_data_bus[40]), .B2(n6157), .ZN(n5661) );
  AOI22D1BWP30P140LVT U5971 ( .A1(i_data_bus[872]), .A2(n6168), .B1(
        i_data_bus[648]), .B2(n6156), .ZN(n5660) );
  AOI22D1BWP30P140LVT U5972 ( .A1(i_data_bus[840]), .A2(n6164), .B1(
        i_data_bus[712]), .B2(n6167), .ZN(n5659) );
  ND4D1BWP30P140LVT U5973 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), 
        .ZN(n5675) );
  MOAI22D1BWP30P140LVT U5974 ( .A1(n5663), .A2(n5920), .B1(i_data_bus[424]), 
        .B2(n5491), .ZN(n5674) );
  AOI22D1BWP30P140LVT U5975 ( .A1(i_data_bus[168]), .A2(n5488), .B1(
        i_data_bus[392]), .B2(n6192), .ZN(n5667) );
  AOI22D1BWP30P140LVT U5976 ( .A1(i_data_bus[936]), .A2(n6191), .B1(
        i_data_bus[456]), .B2(n6187), .ZN(n5666) );
  AOI22D1BWP30P140LVT U5977 ( .A1(i_data_bus[584]), .A2(n6179), .B1(
        i_data_bus[520]), .B2(n6181), .ZN(n5665) );
  AOI22D1BWP30P140LVT U5978 ( .A1(i_data_bus[616]), .A2(n6182), .B1(
        i_data_bus[552]), .B2(n6180), .ZN(n5664) );
  ND4D1BWP30P140LVT U5979 ( .A1(n5667), .A2(n5666), .A3(n5665), .A4(n5664), 
        .ZN(n5673) );
  AOI22D1BWP30P140LVT U5980 ( .A1(i_data_bus[968]), .A2(n6161), .B1(
        i_data_bus[488]), .B2(n6174), .ZN(n5671) );
  AOI22D1BWP30P140LVT U5981 ( .A1(i_data_bus[1000]), .A2(n6177), .B1(
        i_data_bus[904]), .B2(n5474), .ZN(n5670) );
  AOI22D1BWP30P140LVT U5982 ( .A1(i_data_bus[264]), .A2(n6143), .B1(
        i_data_bus[360]), .B2(n6188), .ZN(n5669) );
  AOI22D1BWP30P140LVT U5983 ( .A1(i_data_bus[328]), .A2(n6178), .B1(
        i_data_bus[232]), .B2(n6160), .ZN(n5668) );
  ND4D1BWP30P140LVT U5984 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), 
        .ZN(n5672) );
  NR4D0BWP30P140LVT U5985 ( .A1(n5675), .A2(n5674), .A3(n5673), .A4(n5672), 
        .ZN(n5676) );
  ND4D1BWP30P140LVT U5986 ( .A1(n5679), .A2(n5678), .A3(n5677), .A4(n5676), 
        .ZN(o_data_bus[232]) );
  AOI22D1BWP30P140LVT U5987 ( .A1(i_data_bus[73]), .A2(n6163), .B1(
        i_data_bus[105]), .B2(n6162), .ZN(n5700) );
  AOI22D1BWP30P140LVT U5988 ( .A1(i_data_bus[777]), .A2(n6165), .B1(
        i_data_bus[649]), .B2(n6156), .ZN(n5699) );
  AOI22D1BWP30P140LVT U5989 ( .A1(i_data_bus[969]), .A2(n6161), .B1(
        i_data_bus[329]), .B2(n6178), .ZN(n5698) );
  AOI22D1BWP30P140LVT U5990 ( .A1(i_data_bus[873]), .A2(n6168), .B1(
        i_data_bus[841]), .B2(n6164), .ZN(n5683) );
  AOI22D1BWP30P140LVT U5991 ( .A1(i_data_bus[41]), .A2(n6157), .B1(
        i_data_bus[713]), .B2(n6167), .ZN(n5682) );
  AOI22D1BWP30P140LVT U5992 ( .A1(i_data_bus[9]), .A2(n6169), .B1(
        i_data_bus[809]), .B2(n6166), .ZN(n5681) );
  AOI22D1BWP30P140LVT U5993 ( .A1(i_data_bus[745]), .A2(n6159), .B1(
        i_data_bus[681]), .B2(n6158), .ZN(n5680) );
  ND4D1BWP30P140LVT U5994 ( .A1(n5683), .A2(n5682), .A3(n5681), .A4(n5680), 
        .ZN(n5696) );
  MOAI22D1BWP30P140LVT U5995 ( .A1(n5684), .A2(n5920), .B1(i_data_bus[137]), 
        .B2(n6190), .ZN(n5695) );
  AOI22D1BWP30P140LVT U5996 ( .A1(i_data_bus[905]), .A2(n5474), .B1(
        i_data_bus[937]), .B2(n6191), .ZN(n5688) );
  AOI22D1BWP30P140LVT U5997 ( .A1(i_data_bus[1001]), .A2(n6177), .B1(
        i_data_bus[489]), .B2(n6174), .ZN(n5687) );
  AOI22D1BWP30P140LVT U5998 ( .A1(i_data_bus[617]), .A2(n6182), .B1(
        i_data_bus[553]), .B2(n6180), .ZN(n5686) );
  AOI22D1BWP30P140LVT U5999 ( .A1(i_data_bus[521]), .A2(n6181), .B1(
        i_data_bus[585]), .B2(n6179), .ZN(n5685) );
  ND4D1BWP30P140LVT U6000 ( .A1(n5688), .A2(n5687), .A3(n5686), .A4(n5685), 
        .ZN(n5694) );
  AOI22D1BWP30P140LVT U6001 ( .A1(i_data_bus[233]), .A2(n6160), .B1(
        i_data_bus[265]), .B2(n6143), .ZN(n5692) );
  AOI22D1BWP30P140LVT U6002 ( .A1(i_data_bus[425]), .A2(n5491), .B1(
        i_data_bus[457]), .B2(n6187), .ZN(n5691) );
  AOI22D1BWP30P140LVT U6003 ( .A1(i_data_bus[201]), .A2(n6189), .B1(
        i_data_bus[169]), .B2(n5488), .ZN(n5690) );
  AOI22D1BWP30P140LVT U6004 ( .A1(i_data_bus[361]), .A2(n6188), .B1(
        i_data_bus[393]), .B2(n6192), .ZN(n5689) );
  ND4D1BWP30P140LVT U6005 ( .A1(n5692), .A2(n5691), .A3(n5690), .A4(n5689), 
        .ZN(n5693) );
  NR4D0BWP30P140LVT U6006 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), 
        .ZN(n5697) );
  ND4D1BWP30P140LVT U6007 ( .A1(n5700), .A2(n5699), .A3(n5698), .A4(n5697), 
        .ZN(o_data_bus[233]) );
  AOI22D1BWP30P140LVT U6008 ( .A1(i_data_bus[810]), .A2(n6166), .B1(
        i_data_bus[682]), .B2(n6158), .ZN(n5722) );
  AOI22D1BWP30P140LVT U6009 ( .A1(i_data_bus[10]), .A2(n6169), .B1(
        i_data_bus[874]), .B2(n6168), .ZN(n5721) );
  AOI22D1BWP30P140LVT U6010 ( .A1(i_data_bus[266]), .A2(n6143), .B1(
        i_data_bus[138]), .B2(n6190), .ZN(n5720) );
  AOI22D1BWP30P140LVT U6011 ( .A1(i_data_bus[106]), .A2(n6162), .B1(
        i_data_bus[842]), .B2(n6164), .ZN(n5704) );
  AOI22D1BWP30P140LVT U6012 ( .A1(i_data_bus[650]), .A2(n6156), .B1(
        i_data_bus[746]), .B2(n6159), .ZN(n5703) );
  AOI22D1BWP30P140LVT U6013 ( .A1(i_data_bus[778]), .A2(n6165), .B1(
        i_data_bus[714]), .B2(n6167), .ZN(n5702) );
  AOI22D1BWP30P140LVT U6014 ( .A1(i_data_bus[42]), .A2(n6157), .B1(
        i_data_bus[74]), .B2(n6163), .ZN(n5701) );
  ND4D1BWP30P140LVT U6015 ( .A1(n5704), .A2(n5703), .A3(n5702), .A4(n5701), 
        .ZN(n5718) );
  OAI22D1BWP30P140LVT U6016 ( .A1(n5706), .A2(n5898), .B1(n5705), .B2(n119), 
        .ZN(n5717) );
  AOI22D1BWP30P140LVT U6017 ( .A1(i_data_bus[234]), .A2(n6160), .B1(
        i_data_bus[458]), .B2(n6187), .ZN(n5710) );
  AOI22D1BWP30P140LVT U6018 ( .A1(i_data_bus[1002]), .A2(n6177), .B1(
        i_data_bus[330]), .B2(n6178), .ZN(n5709) );
  AOI22D1BWP30P140LVT U6019 ( .A1(i_data_bus[618]), .A2(n6182), .B1(
        i_data_bus[586]), .B2(n6179), .ZN(n5708) );
  AOI22D1BWP30P140LVT U6020 ( .A1(i_data_bus[554]), .A2(n6180), .B1(
        i_data_bus[522]), .B2(n6181), .ZN(n5707) );
  ND4D1BWP30P140LVT U6021 ( .A1(n5710), .A2(n5709), .A3(n5708), .A4(n5707), 
        .ZN(n5716) );
  AOI22D1BWP30P140LVT U6022 ( .A1(i_data_bus[938]), .A2(n6191), .B1(
        i_data_bus[298]), .B2(n6193), .ZN(n5714) );
  AOI22D1BWP30P140LVT U6023 ( .A1(i_data_bus[906]), .A2(n5474), .B1(
        i_data_bus[202]), .B2(n6189), .ZN(n5713) );
  AOI22D1BWP30P140LVT U6024 ( .A1(i_data_bus[170]), .A2(n5488), .B1(
        i_data_bus[426]), .B2(n5491), .ZN(n5712) );
  AOI22D1BWP30P140LVT U6025 ( .A1(i_data_bus[970]), .A2(n6161), .B1(
        i_data_bus[362]), .B2(n6188), .ZN(n5711) );
  ND4D1BWP30P140LVT U6026 ( .A1(n5714), .A2(n5713), .A3(n5712), .A4(n5711), 
        .ZN(n5715) );
  NR4D0BWP30P140LVT U6027 ( .A1(n5718), .A2(n5717), .A3(n5716), .A4(n5715), 
        .ZN(n5719) );
  ND4D1BWP30P140LVT U6028 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), 
        .ZN(o_data_bus[234]) );
  AOI22D1BWP30P140LVT U6029 ( .A1(i_data_bus[651]), .A2(n6156), .B1(
        i_data_bus[715]), .B2(n6167), .ZN(n5745) );
  AOI22D1BWP30P140LVT U6030 ( .A1(i_data_bus[107]), .A2(n6162), .B1(
        i_data_bus[683]), .B2(n6158), .ZN(n5744) );
  AOI22D1BWP30P140LVT U6031 ( .A1(i_data_bus[907]), .A2(n5474), .B1(
        i_data_bus[203]), .B2(n6189), .ZN(n5743) );
  AOI22D1BWP30P140LVT U6032 ( .A1(i_data_bus[843]), .A2(n6164), .B1(
        i_data_bus[811]), .B2(n6166), .ZN(n5726) );
  AOI22D1BWP30P140LVT U6033 ( .A1(i_data_bus[43]), .A2(n6157), .B1(
        i_data_bus[779]), .B2(n6165), .ZN(n5725) );
  AOI22D1BWP30P140LVT U6034 ( .A1(i_data_bus[11]), .A2(n6169), .B1(
        i_data_bus[875]), .B2(n6168), .ZN(n5724) );
  AOI22D1BWP30P140LVT U6035 ( .A1(i_data_bus[75]), .A2(n6163), .B1(
        i_data_bus[747]), .B2(n6159), .ZN(n5723) );
  ND4D1BWP30P140LVT U6036 ( .A1(n5726), .A2(n5725), .A3(n5724), .A4(n5723), 
        .ZN(n5741) );
  OAI22D1BWP30P140LVT U6037 ( .A1(n5729), .A2(n5728), .B1(n5727), .B2(n6094), 
        .ZN(n5740) );
  AOI22D1BWP30P140LVT U6038 ( .A1(i_data_bus[1003]), .A2(n6177), .B1(
        i_data_bus[139]), .B2(n6190), .ZN(n5733) );
  AOI22D1BWP30P140LVT U6039 ( .A1(i_data_bus[491]), .A2(n6174), .B1(
        i_data_bus[235]), .B2(n6160), .ZN(n5732) );
  AOI22D1BWP30P140LVT U6040 ( .A1(i_data_bus[619]), .A2(n6182), .B1(
        i_data_bus[555]), .B2(n6180), .ZN(n5731) );
  AOI22D1BWP30P140LVT U6041 ( .A1(i_data_bus[523]), .A2(n6181), .B1(
        i_data_bus[587]), .B2(n6179), .ZN(n5730) );
  ND4D1BWP30P140LVT U6042 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), 
        .ZN(n5739) );
  AOI22D1BWP30P140LVT U6043 ( .A1(i_data_bus[939]), .A2(n6191), .B1(
        i_data_bus[395]), .B2(n6192), .ZN(n5737) );
  AOI22D1BWP30P140LVT U6044 ( .A1(i_data_bus[971]), .A2(n6161), .B1(
        i_data_bus[363]), .B2(n6188), .ZN(n5736) );
  AOI22D1BWP30P140LVT U6045 ( .A1(i_data_bus[427]), .A2(n5491), .B1(
        i_data_bus[299]), .B2(n6193), .ZN(n5735) );
  AOI22D1BWP30P140LVT U6046 ( .A1(i_data_bus[171]), .A2(n5488), .B1(
        i_data_bus[267]), .B2(n6143), .ZN(n5734) );
  ND4D1BWP30P140LVT U6047 ( .A1(n5737), .A2(n5736), .A3(n5735), .A4(n5734), 
        .ZN(n5738) );
  NR4D0BWP30P140LVT U6048 ( .A1(n5741), .A2(n5740), .A3(n5739), .A4(n5738), 
        .ZN(n5742) );
  ND4D1BWP30P140LVT U6049 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), 
        .ZN(o_data_bus[235]) );
  AOI22D1BWP30P140LVT U6050 ( .A1(i_data_bus[12]), .A2(n6169), .B1(
        i_data_bus[108]), .B2(n6162), .ZN(n5766) );
  AOI22D1BWP30P140LVT U6051 ( .A1(i_data_bus[44]), .A2(n6157), .B1(
        i_data_bus[684]), .B2(n6158), .ZN(n5765) );
  AOI22D1BWP30P140LVT U6052 ( .A1(i_data_bus[460]), .A2(n6187), .B1(
        i_data_bus[492]), .B2(n6174), .ZN(n5764) );
  AOI22D1BWP30P140LVT U6053 ( .A1(i_data_bus[748]), .A2(n6159), .B1(
        i_data_bus[844]), .B2(n6164), .ZN(n5749) );
  AOI22D1BWP30P140LVT U6054 ( .A1(i_data_bus[780]), .A2(n6165), .B1(
        i_data_bus[876]), .B2(n6168), .ZN(n5748) );
  AOI22D1BWP30P140LVT U6055 ( .A1(i_data_bus[812]), .A2(n6166), .B1(
        i_data_bus[652]), .B2(n6156), .ZN(n5747) );
  AOI22D1BWP30P140LVT U6056 ( .A1(i_data_bus[76]), .A2(n6163), .B1(
        i_data_bus[716]), .B2(n6167), .ZN(n5746) );
  ND4D1BWP30P140LVT U6057 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), 
        .ZN(n5762) );
  MOAI22D1BWP30P140LVT U6058 ( .A1(n5750), .A2(n6175), .B1(i_data_bus[236]), 
        .B2(n6160), .ZN(n5761) );
  AOI22D1BWP30P140LVT U6059 ( .A1(i_data_bus[1004]), .A2(n6177), .B1(
        i_data_bus[300]), .B2(n6193), .ZN(n5754) );
  AOI22D1BWP30P140LVT U6060 ( .A1(i_data_bus[908]), .A2(n5474), .B1(
        i_data_bus[972]), .B2(n6161), .ZN(n5753) );
  AOI22D1BWP30P140LVT U6061 ( .A1(i_data_bus[524]), .A2(n6181), .B1(
        i_data_bus[588]), .B2(n6179), .ZN(n5752) );
  AOI22D1BWP30P140LVT U6062 ( .A1(i_data_bus[620]), .A2(n6182), .B1(
        i_data_bus[556]), .B2(n6180), .ZN(n5751) );
  ND4D1BWP30P140LVT U6063 ( .A1(n5754), .A2(n5753), .A3(n5752), .A4(n5751), 
        .ZN(n5760) );
  AOI22D1BWP30P140LVT U6064 ( .A1(i_data_bus[940]), .A2(n6191), .B1(
        i_data_bus[140]), .B2(n6190), .ZN(n5758) );
  AOI22D1BWP30P140LVT U6065 ( .A1(i_data_bus[268]), .A2(n6143), .B1(
        i_data_bus[204]), .B2(n6189), .ZN(n5757) );
  AOI22D1BWP30P140LVT U6066 ( .A1(i_data_bus[364]), .A2(n6188), .B1(
        i_data_bus[396]), .B2(n6192), .ZN(n5756) );
  AOI22D1BWP30P140LVT U6067 ( .A1(i_data_bus[428]), .A2(n5491), .B1(
        i_data_bus[332]), .B2(n6178), .ZN(n5755) );
  ND4D1BWP30P140LVT U6068 ( .A1(n5758), .A2(n5757), .A3(n5756), .A4(n5755), 
        .ZN(n5759) );
  NR4D0BWP30P140LVT U6069 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), 
        .ZN(n5763) );
  ND4D1BWP30P140LVT U6070 ( .A1(n5766), .A2(n5765), .A3(n5764), .A4(n5763), 
        .ZN(o_data_bus[236]) );
  AOI22D1BWP30P140LVT U6071 ( .A1(i_data_bus[45]), .A2(n6157), .B1(
        i_data_bus[717]), .B2(n6167), .ZN(n5787) );
  AOI22D1BWP30P140LVT U6072 ( .A1(i_data_bus[845]), .A2(n6164), .B1(
        i_data_bus[813]), .B2(n6166), .ZN(n5786) );
  AOI22D1BWP30P140LVT U6073 ( .A1(i_data_bus[237]), .A2(n6160), .B1(
        i_data_bus[141]), .B2(n6190), .ZN(n5785) );
  AOI22D1BWP30P140LVT U6074 ( .A1(i_data_bus[781]), .A2(n6165), .B1(
        i_data_bus[749]), .B2(n6159), .ZN(n5770) );
  AOI22D1BWP30P140LVT U6075 ( .A1(i_data_bus[77]), .A2(n6163), .B1(
        i_data_bus[685]), .B2(n6158), .ZN(n5769) );
  AOI22D1BWP30P140LVT U6076 ( .A1(i_data_bus[109]), .A2(n6162), .B1(
        i_data_bus[877]), .B2(n6168), .ZN(n5768) );
  AOI22D1BWP30P140LVT U6077 ( .A1(i_data_bus[13]), .A2(n6169), .B1(
        i_data_bus[653]), .B2(n6156), .ZN(n5767) );
  ND4D1BWP30P140LVT U6078 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), 
        .ZN(n5783) );
  MOAI22D1BWP30P140LVT U6079 ( .A1(n5771), .A2(n6175), .B1(i_data_bus[365]), 
        .B2(n6188), .ZN(n5782) );
  AOI22D1BWP30P140LVT U6080 ( .A1(i_data_bus[909]), .A2(n5474), .B1(
        i_data_bus[461]), .B2(n6187), .ZN(n5775) );
  AOI22D1BWP30P140LVT U6081 ( .A1(i_data_bus[973]), .A2(n6161), .B1(
        i_data_bus[1005]), .B2(n6177), .ZN(n5774) );
  AOI22D1BWP30P140LVT U6082 ( .A1(i_data_bus[621]), .A2(n6182), .B1(
        i_data_bus[557]), .B2(n6180), .ZN(n5773) );
  AOI22D1BWP30P140LVT U6083 ( .A1(i_data_bus[525]), .A2(n6181), .B1(
        i_data_bus[589]), .B2(n6179), .ZN(n5772) );
  ND4D1BWP30P140LVT U6084 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), 
        .ZN(n5781) );
  AOI22D1BWP30P140LVT U6085 ( .A1(i_data_bus[269]), .A2(n6143), .B1(
        i_data_bus[429]), .B2(n5491), .ZN(n5779) );
  AOI22D1BWP30P140LVT U6086 ( .A1(i_data_bus[397]), .A2(n6192), .B1(
        i_data_bus[493]), .B2(n6174), .ZN(n5778) );
  AOI22D1BWP30P140LVT U6087 ( .A1(i_data_bus[941]), .A2(n6191), .B1(
        i_data_bus[333]), .B2(n6178), .ZN(n5777) );
  AOI22D1BWP30P140LVT U6088 ( .A1(i_data_bus[205]), .A2(n6189), .B1(
        i_data_bus[301]), .B2(n6193), .ZN(n5776) );
  ND4D1BWP30P140LVT U6089 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), 
        .ZN(n5780) );
  NR4D0BWP30P140LVT U6090 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), 
        .ZN(n5784) );
  ND4D1BWP30P140LVT U6091 ( .A1(n5787), .A2(n5786), .A3(n5785), .A4(n5784), 
        .ZN(o_data_bus[237]) );
  AOI22D1BWP30P140LVT U6092 ( .A1(i_data_bus[46]), .A2(n6157), .B1(
        i_data_bus[654]), .B2(n6156), .ZN(n5808) );
  AOI22D1BWP30P140LVT U6093 ( .A1(i_data_bus[110]), .A2(n6162), .B1(
        i_data_bus[78]), .B2(n6163), .ZN(n5807) );
  AOI22D1BWP30P140LVT U6094 ( .A1(i_data_bus[942]), .A2(n6191), .B1(
        i_data_bus[174]), .B2(n5488), .ZN(n5806) );
  AOI22D1BWP30P140LVT U6095 ( .A1(i_data_bus[814]), .A2(n6166), .B1(
        i_data_bus[846]), .B2(n6164), .ZN(n5791) );
  AOI22D1BWP30P140LVT U6096 ( .A1(i_data_bus[14]), .A2(n6169), .B1(
        i_data_bus[878]), .B2(n6168), .ZN(n5790) );
  AOI22D1BWP30P140LVT U6097 ( .A1(i_data_bus[782]), .A2(n6165), .B1(
        i_data_bus[686]), .B2(n6158), .ZN(n5789) );
  AOI22D1BWP30P140LVT U6098 ( .A1(i_data_bus[750]), .A2(n6159), .B1(
        i_data_bus[718]), .B2(n6167), .ZN(n5788) );
  ND4D1BWP30P140LVT U6099 ( .A1(n5791), .A2(n5790), .A3(n5789), .A4(n5788), 
        .ZN(n5804) );
  MOAI22D1BWP30P140LVT U6100 ( .A1(n5792), .A2(n5898), .B1(i_data_bus[302]), 
        .B2(n6193), .ZN(n5803) );
  AOI22D1BWP30P140LVT U6101 ( .A1(i_data_bus[270]), .A2(n6143), .B1(
        i_data_bus[206]), .B2(n6189), .ZN(n5796) );
  AOI22D1BWP30P140LVT U6102 ( .A1(i_data_bus[910]), .A2(n5474), .B1(
        i_data_bus[334]), .B2(n6178), .ZN(n5795) );
  AOI22D1BWP30P140LVT U6103 ( .A1(i_data_bus[558]), .A2(n6180), .B1(
        i_data_bus[526]), .B2(n6181), .ZN(n5794) );
  AOI22D1BWP30P140LVT U6104 ( .A1(i_data_bus[590]), .A2(n6179), .B1(
        i_data_bus[622]), .B2(n6182), .ZN(n5793) );
  ND4D1BWP30P140LVT U6105 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), 
        .ZN(n5802) );
  AOI22D1BWP30P140LVT U6106 ( .A1(i_data_bus[366]), .A2(n6188), .B1(
        i_data_bus[462]), .B2(n6187), .ZN(n5800) );
  AOI22D1BWP30P140LVT U6107 ( .A1(i_data_bus[142]), .A2(n6190), .B1(
        i_data_bus[398]), .B2(n6192), .ZN(n5799) );
  AOI22D1BWP30P140LVT U6108 ( .A1(i_data_bus[1006]), .A2(n6177), .B1(
        i_data_bus[430]), .B2(n5491), .ZN(n5798) );
  AOI22D1BWP30P140LVT U6109 ( .A1(i_data_bus[974]), .A2(n6161), .B1(
        i_data_bus[238]), .B2(n6160), .ZN(n5797) );
  ND4D1BWP30P140LVT U6110 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), 
        .ZN(n5801) );
  NR4D0BWP30P140LVT U6111 ( .A1(n5804), .A2(n5803), .A3(n5802), .A4(n5801), 
        .ZN(n5805) );
  ND4D1BWP30P140LVT U6112 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), 
        .ZN(o_data_bus[238]) );
  AOI22D1BWP30P140LVT U6113 ( .A1(i_data_bus[111]), .A2(n6162), .B1(
        i_data_bus[687]), .B2(n6158), .ZN(n5829) );
  AOI22D1BWP30P140LVT U6114 ( .A1(i_data_bus[47]), .A2(n6157), .B1(
        i_data_bus[783]), .B2(n6165), .ZN(n5828) );
  AOI22D1BWP30P140LVT U6115 ( .A1(i_data_bus[431]), .A2(n5491), .B1(
        i_data_bus[463]), .B2(n6187), .ZN(n5827) );
  AOI22D1BWP30P140LVT U6116 ( .A1(i_data_bus[719]), .A2(n6167), .B1(
        i_data_bus[655]), .B2(n6156), .ZN(n5812) );
  AOI22D1BWP30P140LVT U6117 ( .A1(i_data_bus[15]), .A2(n6169), .B1(
        i_data_bus[751]), .B2(n6159), .ZN(n5811) );
  AOI22D1BWP30P140LVT U6118 ( .A1(i_data_bus[879]), .A2(n6168), .B1(
        i_data_bus[815]), .B2(n6166), .ZN(n5810) );
  AOI22D1BWP30P140LVT U6119 ( .A1(i_data_bus[79]), .A2(n6163), .B1(
        i_data_bus[847]), .B2(n6164), .ZN(n5809) );
  ND4D1BWP30P140LVT U6120 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), 
        .ZN(n5825) );
  MOAI22D1BWP30P140LVT U6121 ( .A1(n5813), .A2(n6116), .B1(i_data_bus[335]), 
        .B2(n6178), .ZN(n5824) );
  AOI22D1BWP30P140LVT U6122 ( .A1(i_data_bus[911]), .A2(n5474), .B1(
        i_data_bus[943]), .B2(n6191), .ZN(n5817) );
  AOI22D1BWP30P140LVT U6123 ( .A1(i_data_bus[1007]), .A2(n6177), .B1(
        i_data_bus[239]), .B2(n6160), .ZN(n5816) );
  AOI22D1BWP30P140LVT U6124 ( .A1(i_data_bus[591]), .A2(n6179), .B1(
        i_data_bus[527]), .B2(n6181), .ZN(n5815) );
  AOI22D1BWP30P140LVT U6125 ( .A1(i_data_bus[559]), .A2(n6180), .B1(
        i_data_bus[623]), .B2(n6182), .ZN(n5814) );
  ND4D1BWP30P140LVT U6126 ( .A1(n5817), .A2(n5816), .A3(n5815), .A4(n5814), 
        .ZN(n5823) );
  AOI22D1BWP30P140LVT U6127 ( .A1(i_data_bus[175]), .A2(n5488), .B1(
        i_data_bus[143]), .B2(n6190), .ZN(n5821) );
  AOI22D1BWP30P140LVT U6128 ( .A1(i_data_bus[207]), .A2(n6189), .B1(
        i_data_bus[399]), .B2(n6192), .ZN(n5820) );
  AOI22D1BWP30P140LVT U6129 ( .A1(i_data_bus[975]), .A2(n6161), .B1(
        i_data_bus[271]), .B2(n6143), .ZN(n5819) );
  AOI22D1BWP30P140LVT U6130 ( .A1(i_data_bus[495]), .A2(n6174), .B1(
        i_data_bus[303]), .B2(n6193), .ZN(n5818) );
  ND4D1BWP30P140LVT U6131 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), 
        .ZN(n5822) );
  NR4D0BWP30P140LVT U6132 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), 
        .ZN(n5826) );
  ND4D1BWP30P140LVT U6133 ( .A1(n5829), .A2(n5828), .A3(n5827), .A4(n5826), 
        .ZN(o_data_bus[239]) );
  AOI22D1BWP30P140LVT U6134 ( .A1(i_data_bus[880]), .A2(n6168), .B1(
        i_data_bus[656]), .B2(n6156), .ZN(n5850) );
  AOI22D1BWP30P140LVT U6135 ( .A1(i_data_bus[80]), .A2(n6163), .B1(
        i_data_bus[720]), .B2(n6167), .ZN(n5849) );
  AOI22D1BWP30P140LVT U6136 ( .A1(i_data_bus[304]), .A2(n6193), .B1(
        i_data_bus[272]), .B2(n6143), .ZN(n5848) );
  AOI22D1BWP30P140LVT U6137 ( .A1(i_data_bus[784]), .A2(n6165), .B1(
        i_data_bus[848]), .B2(n6164), .ZN(n5833) );
  AOI22D1BWP30P140LVT U6138 ( .A1(i_data_bus[112]), .A2(n6162), .B1(
        i_data_bus[688]), .B2(n6158), .ZN(n5832) );
  AOI22D1BWP30P140LVT U6139 ( .A1(i_data_bus[48]), .A2(n6157), .B1(
        i_data_bus[752]), .B2(n6159), .ZN(n5831) );
  AOI22D1BWP30P140LVT U6140 ( .A1(i_data_bus[16]), .A2(n6169), .B1(
        i_data_bus[816]), .B2(n6166), .ZN(n5830) );
  ND4D1BWP30P140LVT U6141 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), 
        .ZN(n5846) );
  MOAI22D1BWP30P140LVT U6142 ( .A1(n5834), .A2(n119), .B1(i_data_bus[208]), 
        .B2(n6189), .ZN(n5845) );
  AOI22D1BWP30P140LVT U6143 ( .A1(i_data_bus[1008]), .A2(n6177), .B1(
        i_data_bus[432]), .B2(n5491), .ZN(n5838) );
  AOI22D1BWP30P140LVT U6144 ( .A1(i_data_bus[944]), .A2(n6191), .B1(
        i_data_bus[144]), .B2(n6190), .ZN(n5837) );
  AOI22D1BWP30P140LVT U6145 ( .A1(i_data_bus[560]), .A2(n6180), .B1(
        i_data_bus[592]), .B2(n6179), .ZN(n5836) );
  AOI22D1BWP30P140LVT U6146 ( .A1(i_data_bus[528]), .A2(n6181), .B1(
        i_data_bus[624]), .B2(n6182), .ZN(n5835) );
  ND4D1BWP30P140LVT U6147 ( .A1(n5838), .A2(n5837), .A3(n5836), .A4(n5835), 
        .ZN(n5844) );
  AOI22D1BWP30P140LVT U6148 ( .A1(i_data_bus[336]), .A2(n6178), .B1(
        i_data_bus[496]), .B2(n6174), .ZN(n5842) );
  AOI22D1BWP30P140LVT U6149 ( .A1(i_data_bus[976]), .A2(n6161), .B1(
        i_data_bus[464]), .B2(n6187), .ZN(n5841) );
  AOI22D1BWP30P140LVT U6150 ( .A1(i_data_bus[912]), .A2(n5474), .B1(
        i_data_bus[240]), .B2(n6160), .ZN(n5840) );
  AOI22D1BWP30P140LVT U6151 ( .A1(i_data_bus[176]), .A2(n5488), .B1(
        i_data_bus[368]), .B2(n6188), .ZN(n5839) );
  ND4D1BWP30P140LVT U6152 ( .A1(n5842), .A2(n5841), .A3(n5840), .A4(n5839), 
        .ZN(n5843) );
  NR4D0BWP30P140LVT U6153 ( .A1(n5846), .A2(n5845), .A3(n5844), .A4(n5843), 
        .ZN(n5847) );
  ND4D1BWP30P140LVT U6154 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), 
        .ZN(o_data_bus[240]) );
  AOI22D1BWP30P140LVT U6155 ( .A1(i_data_bus[657]), .A2(n6156), .B1(
        i_data_bus[753]), .B2(n6159), .ZN(n5871) );
  AOI22D1BWP30P140LVT U6156 ( .A1(i_data_bus[49]), .A2(n6157), .B1(
        i_data_bus[689]), .B2(n6158), .ZN(n5870) );
  AOI22D1BWP30P140LVT U6157 ( .A1(i_data_bus[1009]), .A2(n6177), .B1(
        i_data_bus[401]), .B2(n6192), .ZN(n5869) );
  AOI22D1BWP30P140LVT U6158 ( .A1(i_data_bus[17]), .A2(n6169), .B1(
        i_data_bus[849]), .B2(n6164), .ZN(n5854) );
  AOI22D1BWP30P140LVT U6159 ( .A1(i_data_bus[785]), .A2(n6165), .B1(
        i_data_bus[721]), .B2(n6167), .ZN(n5853) );
  AOI22D1BWP30P140LVT U6160 ( .A1(i_data_bus[881]), .A2(n6168), .B1(
        i_data_bus[817]), .B2(n6166), .ZN(n5852) );
  AOI22D1BWP30P140LVT U6161 ( .A1(i_data_bus[81]), .A2(n6163), .B1(
        i_data_bus[113]), .B2(n6162), .ZN(n5851) );
  ND4D1BWP30P140LVT U6162 ( .A1(n5854), .A2(n5853), .A3(n5852), .A4(n5851), 
        .ZN(n5867) );
  MOAI22D1BWP30P140LVT U6163 ( .A1(n5855), .A2(n6116), .B1(i_data_bus[497]), 
        .B2(n6174), .ZN(n5866) );
  AOI22D1BWP30P140LVT U6164 ( .A1(i_data_bus[241]), .A2(n6160), .B1(
        i_data_bus[273]), .B2(n6143), .ZN(n5859) );
  AOI22D1BWP30P140LVT U6165 ( .A1(i_data_bus[977]), .A2(n6161), .B1(
        i_data_bus[433]), .B2(n5491), .ZN(n5858) );
  AOI22D1BWP30P140LVT U6166 ( .A1(i_data_bus[593]), .A2(n6179), .B1(
        i_data_bus[561]), .B2(n6180), .ZN(n5857) );
  AOI22D1BWP30P140LVT U6167 ( .A1(i_data_bus[625]), .A2(n6182), .B1(
        i_data_bus[529]), .B2(n6181), .ZN(n5856) );
  ND4D1BWP30P140LVT U6168 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), 
        .ZN(n5865) );
  AOI22D1BWP30P140LVT U6169 ( .A1(i_data_bus[337]), .A2(n6178), .B1(
        i_data_bus[145]), .B2(n6190), .ZN(n5863) );
  AOI22D1BWP30P140LVT U6170 ( .A1(i_data_bus[209]), .A2(n6189), .B1(
        i_data_bus[305]), .B2(n6193), .ZN(n5862) );
  AOI22D1BWP30P140LVT U6171 ( .A1(i_data_bus[945]), .A2(n6191), .B1(
        i_data_bus[465]), .B2(n6187), .ZN(n5861) );
  AOI22D1BWP30P140LVT U6172 ( .A1(i_data_bus[913]), .A2(n5474), .B1(
        i_data_bus[177]), .B2(n5488), .ZN(n5860) );
  ND4D1BWP30P140LVT U6173 ( .A1(n5863), .A2(n5862), .A3(n5861), .A4(n5860), 
        .ZN(n5864) );
  NR4D0BWP30P140LVT U6174 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), 
        .ZN(n5868) );
  ND4D1BWP30P140LVT U6175 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), 
        .ZN(o_data_bus[241]) );
  AOI22D1BWP30P140LVT U6176 ( .A1(i_data_bus[658]), .A2(n6156), .B1(
        i_data_bus[754]), .B2(n6159), .ZN(n5893) );
  AOI22D1BWP30P140LVT U6177 ( .A1(i_data_bus[722]), .A2(n6167), .B1(
        i_data_bus[818]), .B2(n6166), .ZN(n5892) );
  AOI22D1BWP30P140LVT U6178 ( .A1(i_data_bus[178]), .A2(n5488), .B1(
        i_data_bus[306]), .B2(n6193), .ZN(n5891) );
  AOI22D1BWP30P140LVT U6179 ( .A1(i_data_bus[82]), .A2(n6163), .B1(
        i_data_bus[882]), .B2(n6168), .ZN(n5875) );
  AOI22D1BWP30P140LVT U6180 ( .A1(i_data_bus[690]), .A2(n6158), .B1(
        i_data_bus[850]), .B2(n6164), .ZN(n5874) );
  AOI22D1BWP30P140LVT U6181 ( .A1(i_data_bus[50]), .A2(n6157), .B1(
        i_data_bus[786]), .B2(n6165), .ZN(n5873) );
  AOI22D1BWP30P140LVT U6182 ( .A1(i_data_bus[114]), .A2(n6162), .B1(
        i_data_bus[18]), .B2(n6169), .ZN(n5872) );
  ND4D1BWP30P140LVT U6183 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), 
        .ZN(n5889) );
  MOAI22D1BWP30P140LVT U6184 ( .A1(n5877), .A2(n5876), .B1(i_data_bus[978]), 
        .B2(n6161), .ZN(n5888) );
  AOI22D1BWP30P140LVT U6185 ( .A1(i_data_bus[914]), .A2(n5474), .B1(
        i_data_bus[498]), .B2(n6174), .ZN(n5881) );
  AOI22D1BWP30P140LVT U6186 ( .A1(i_data_bus[1010]), .A2(n6177), .B1(
        i_data_bus[338]), .B2(n6178), .ZN(n5880) );
  AOI22D1BWP30P140LVT U6187 ( .A1(i_data_bus[530]), .A2(n6181), .B1(
        i_data_bus[562]), .B2(n6180), .ZN(n5879) );
  AOI22D1BWP30P140LVT U6188 ( .A1(i_data_bus[626]), .A2(n6182), .B1(
        i_data_bus[594]), .B2(n6179), .ZN(n5878) );
  ND4D1BWP30P140LVT U6189 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), 
        .ZN(n5887) );
  AOI22D1BWP30P140LVT U6190 ( .A1(i_data_bus[946]), .A2(n6191), .B1(
        i_data_bus[274]), .B2(n6143), .ZN(n5885) );
  AOI22D1BWP30P140LVT U6191 ( .A1(i_data_bus[402]), .A2(n6192), .B1(
        i_data_bus[210]), .B2(n6189), .ZN(n5884) );
  AOI22D1BWP30P140LVT U6192 ( .A1(i_data_bus[370]), .A2(n6188), .B1(
        i_data_bus[466]), .B2(n6187), .ZN(n5883) );
  AOI22D1BWP30P140LVT U6193 ( .A1(i_data_bus[242]), .A2(n6160), .B1(
        i_data_bus[434]), .B2(n5491), .ZN(n5882) );
  ND4D1BWP30P140LVT U6194 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), 
        .ZN(n5886) );
  NR4D0BWP30P140LVT U6195 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), 
        .ZN(n5890) );
  ND4D1BWP30P140LVT U6196 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), 
        .ZN(o_data_bus[242]) );
  AOI22D1BWP30P140LVT U6197 ( .A1(i_data_bus[115]), .A2(n6162), .B1(
        i_data_bus[819]), .B2(n6166), .ZN(n5915) );
  AOI22D1BWP30P140LVT U6198 ( .A1(i_data_bus[691]), .A2(n6158), .B1(
        i_data_bus[723]), .B2(n6167), .ZN(n5914) );
  AOI22D1BWP30P140LVT U6199 ( .A1(i_data_bus[307]), .A2(n6193), .B1(
        i_data_bus[275]), .B2(n6143), .ZN(n5913) );
  AOI22D1BWP30P140LVT U6200 ( .A1(i_data_bus[83]), .A2(n6163), .B1(
        i_data_bus[659]), .B2(n6156), .ZN(n5897) );
  AOI22D1BWP30P140LVT U6201 ( .A1(i_data_bus[19]), .A2(n6169), .B1(
        i_data_bus[851]), .B2(n6164), .ZN(n5896) );
  AOI22D1BWP30P140LVT U6202 ( .A1(i_data_bus[755]), .A2(n6159), .B1(
        i_data_bus[883]), .B2(n6168), .ZN(n5895) );
  AOI22D1BWP30P140LVT U6203 ( .A1(i_data_bus[51]), .A2(n6157), .B1(
        i_data_bus[787]), .B2(n6165), .ZN(n5894) );
  ND4D1BWP30P140LVT U6204 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), 
        .ZN(n5911) );
  MOAI22D1BWP30P140LVT U6205 ( .A1(n5899), .A2(n5898), .B1(i_data_bus[947]), 
        .B2(n6191), .ZN(n5910) );
  AOI22D1BWP30P140LVT U6206 ( .A1(i_data_bus[979]), .A2(n6161), .B1(
        i_data_bus[211]), .B2(n6189), .ZN(n5903) );
  AOI22D1BWP30P140LVT U6207 ( .A1(i_data_bus[1011]), .A2(n6177), .B1(
        i_data_bus[403]), .B2(n6192), .ZN(n5902) );
  AOI22D1BWP30P140LVT U6208 ( .A1(i_data_bus[531]), .A2(n6181), .B1(
        i_data_bus[595]), .B2(n6179), .ZN(n5901) );
  AOI22D1BWP30P140LVT U6209 ( .A1(i_data_bus[563]), .A2(n6180), .B1(
        i_data_bus[627]), .B2(n6182), .ZN(n5900) );
  ND4D1BWP30P140LVT U6210 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), 
        .ZN(n5909) );
  AOI22D1BWP30P140LVT U6211 ( .A1(i_data_bus[339]), .A2(n6178), .B1(
        i_data_bus[435]), .B2(n5491), .ZN(n5907) );
  AOI22D1BWP30P140LVT U6212 ( .A1(i_data_bus[915]), .A2(n5474), .B1(
        i_data_bus[467]), .B2(n6187), .ZN(n5906) );
  AOI22D1BWP30P140LVT U6213 ( .A1(i_data_bus[371]), .A2(n6188), .B1(
        i_data_bus[243]), .B2(n6160), .ZN(n5905) );
  AOI22D1BWP30P140LVT U6214 ( .A1(i_data_bus[179]), .A2(n5488), .B1(
        i_data_bus[147]), .B2(n6190), .ZN(n5904) );
  ND4D1BWP30P140LVT U6215 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), 
        .ZN(n5908) );
  NR4D0BWP30P140LVT U6216 ( .A1(n5911), .A2(n5910), .A3(n5909), .A4(n5908), 
        .ZN(n5912) );
  ND4D1BWP30P140LVT U6217 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), 
        .ZN(o_data_bus[243]) );
  AOI22D1BWP30P140LVT U6218 ( .A1(i_data_bus[788]), .A2(n6165), .B1(
        i_data_bus[692]), .B2(n6158), .ZN(n5937) );
  AOI22D1BWP30P140LVT U6219 ( .A1(i_data_bus[52]), .A2(n6157), .B1(
        i_data_bus[84]), .B2(n6163), .ZN(n5936) );
  AOI22D1BWP30P140LVT U6220 ( .A1(i_data_bus[244]), .A2(n6160), .B1(
        i_data_bus[436]), .B2(n5491), .ZN(n5935) );
  AOI22D1BWP30P140LVT U6221 ( .A1(i_data_bus[20]), .A2(n6169), .B1(
        i_data_bus[724]), .B2(n6167), .ZN(n5919) );
  AOI22D1BWP30P140LVT U6222 ( .A1(i_data_bus[820]), .A2(n6166), .B1(
        i_data_bus[660]), .B2(n6156), .ZN(n5918) );
  AOI22D1BWP30P140LVT U6223 ( .A1(i_data_bus[116]), .A2(n6162), .B1(
        i_data_bus[756]), .B2(n6159), .ZN(n5917) );
  AOI22D1BWP30P140LVT U6224 ( .A1(i_data_bus[852]), .A2(n6164), .B1(
        i_data_bus[884]), .B2(n6168), .ZN(n5916) );
  ND4D1BWP30P140LVT U6225 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), 
        .ZN(n5933) );
  MOAI22D1BWP30P140LVT U6226 ( .A1(n5921), .A2(n5920), .B1(i_data_bus[276]), 
        .B2(n6143), .ZN(n5932) );
  AOI22D1BWP30P140LVT U6227 ( .A1(i_data_bus[948]), .A2(n6191), .B1(
        i_data_bus[148]), .B2(n6190), .ZN(n5925) );
  AOI22D1BWP30P140LVT U6228 ( .A1(i_data_bus[980]), .A2(n6161), .B1(
        i_data_bus[404]), .B2(n6192), .ZN(n5924) );
  AOI22D1BWP30P140LVT U6229 ( .A1(i_data_bus[596]), .A2(n6179), .B1(
        i_data_bus[564]), .B2(n6180), .ZN(n5923) );
  AOI22D1BWP30P140LVT U6230 ( .A1(i_data_bus[532]), .A2(n6181), .B1(
        i_data_bus[628]), .B2(n6182), .ZN(n5922) );
  ND4D1BWP30P140LVT U6231 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), 
        .ZN(n5931) );
  AOI22D1BWP30P140LVT U6232 ( .A1(i_data_bus[340]), .A2(n6178), .B1(
        i_data_bus[500]), .B2(n6174), .ZN(n5929) );
  AOI22D1BWP30P140LVT U6233 ( .A1(i_data_bus[1012]), .A2(n6177), .B1(
        i_data_bus[180]), .B2(n5488), .ZN(n5928) );
  AOI22D1BWP30P140LVT U6234 ( .A1(i_data_bus[916]), .A2(n5474), .B1(
        i_data_bus[468]), .B2(n6187), .ZN(n5927) );
  AOI22D1BWP30P140LVT U6235 ( .A1(i_data_bus[212]), .A2(n6189), .B1(
        i_data_bus[372]), .B2(n6188), .ZN(n5926) );
  ND4D1BWP30P140LVT U6236 ( .A1(n5929), .A2(n5928), .A3(n5927), .A4(n5926), 
        .ZN(n5930) );
  NR4D0BWP30P140LVT U6237 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), 
        .ZN(n5934) );
  ND4D1BWP30P140LVT U6238 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), 
        .ZN(o_data_bus[244]) );
  AOI22D1BWP30P140LVT U6239 ( .A1(i_data_bus[789]), .A2(n6165), .B1(
        i_data_bus[725]), .B2(n6167), .ZN(n5958) );
  AOI22D1BWP30P140LVT U6240 ( .A1(i_data_bus[53]), .A2(n6157), .B1(
        i_data_bus[821]), .B2(n6166), .ZN(n5957) );
  AOI22D1BWP30P140LVT U6241 ( .A1(i_data_bus[213]), .A2(n6189), .B1(
        i_data_bus[277]), .B2(n6143), .ZN(n5956) );
  AOI22D1BWP30P140LVT U6242 ( .A1(i_data_bus[21]), .A2(n6169), .B1(
        i_data_bus[853]), .B2(n6164), .ZN(n5941) );
  AOI22D1BWP30P140LVT U6243 ( .A1(i_data_bus[661]), .A2(n6156), .B1(
        i_data_bus[693]), .B2(n6158), .ZN(n5940) );
  AOI22D1BWP30P140LVT U6244 ( .A1(i_data_bus[117]), .A2(n6162), .B1(
        i_data_bus[757]), .B2(n6159), .ZN(n5939) );
  AOI22D1BWP30P140LVT U6245 ( .A1(i_data_bus[85]), .A2(n6163), .B1(
        i_data_bus[885]), .B2(n6168), .ZN(n5938) );
  ND4D1BWP30P140LVT U6246 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), 
        .ZN(n5954) );
  MOAI22D1BWP30P140LVT U6247 ( .A1(n5942), .A2(n6116), .B1(i_data_bus[181]), 
        .B2(n5488), .ZN(n5953) );
  AOI22D1BWP30P140LVT U6248 ( .A1(i_data_bus[981]), .A2(n6161), .B1(
        i_data_bus[341]), .B2(n6178), .ZN(n5946) );
  AOI22D1BWP30P140LVT U6249 ( .A1(i_data_bus[917]), .A2(n5474), .B1(
        i_data_bus[1013]), .B2(n6177), .ZN(n5945) );
  AOI22D1BWP30P140LVT U6250 ( .A1(i_data_bus[597]), .A2(n6179), .B1(
        i_data_bus[565]), .B2(n6180), .ZN(n5944) );
  AOI22D1BWP30P140LVT U6251 ( .A1(i_data_bus[629]), .A2(n6182), .B1(
        i_data_bus[533]), .B2(n6181), .ZN(n5943) );
  ND4D1BWP30P140LVT U6252 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), 
        .ZN(n5952) );
  AOI22D1BWP30P140LVT U6253 ( .A1(i_data_bus[501]), .A2(n6174), .B1(
        i_data_bus[469]), .B2(n6187), .ZN(n5950) );
  AOI22D1BWP30P140LVT U6254 ( .A1(i_data_bus[949]), .A2(n6191), .B1(
        i_data_bus[149]), .B2(n6190), .ZN(n5949) );
  AOI22D1BWP30P140LVT U6255 ( .A1(i_data_bus[437]), .A2(n5491), .B1(
        i_data_bus[245]), .B2(n6160), .ZN(n5948) );
  AOI22D1BWP30P140LVT U6256 ( .A1(i_data_bus[309]), .A2(n6193), .B1(
        i_data_bus[405]), .B2(n6192), .ZN(n5947) );
  ND4D1BWP30P140LVT U6257 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), 
        .ZN(n5951) );
  NR4D0BWP30P140LVT U6258 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), 
        .ZN(n5955) );
  ND4D1BWP30P140LVT U6259 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), 
        .ZN(o_data_bus[245]) );
  AOI22D1BWP30P140LVT U6260 ( .A1(i_data_bus[822]), .A2(n6166), .B1(
        i_data_bus[662]), .B2(n6156), .ZN(n5980) );
  AOI22D1BWP30P140LVT U6261 ( .A1(i_data_bus[54]), .A2(n6157), .B1(
        i_data_bus[118]), .B2(n6162), .ZN(n5979) );
  AOI22D1BWP30P140LVT U6262 ( .A1(i_data_bus[182]), .A2(n5488), .B1(
        i_data_bus[470]), .B2(n6187), .ZN(n5978) );
  AOI22D1BWP30P140LVT U6263 ( .A1(i_data_bus[86]), .A2(n6163), .B1(
        i_data_bus[726]), .B2(n6167), .ZN(n5962) );
  AOI22D1BWP30P140LVT U6264 ( .A1(i_data_bus[22]), .A2(n6169), .B1(
        i_data_bus[790]), .B2(n6165), .ZN(n5961) );
  AOI22D1BWP30P140LVT U6265 ( .A1(i_data_bus[886]), .A2(n6168), .B1(
        i_data_bus[854]), .B2(n6164), .ZN(n5960) );
  AOI22D1BWP30P140LVT U6266 ( .A1(i_data_bus[694]), .A2(n6158), .B1(
        i_data_bus[758]), .B2(n6159), .ZN(n5959) );
  ND4D1BWP30P140LVT U6267 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), 
        .ZN(n5976) );
  MOAI22D1BWP30P140LVT U6268 ( .A1(n5964), .A2(n5963), .B1(i_data_bus[246]), 
        .B2(n6160), .ZN(n5975) );
  AOI22D1BWP30P140LVT U6269 ( .A1(i_data_bus[502]), .A2(n6174), .B1(
        i_data_bus[310]), .B2(n6193), .ZN(n5968) );
  AOI22D1BWP30P140LVT U6270 ( .A1(i_data_bus[1014]), .A2(n6177), .B1(
        i_data_bus[342]), .B2(n6178), .ZN(n5967) );
  AOI22D1BWP30P140LVT U6271 ( .A1(i_data_bus[534]), .A2(n6181), .B1(
        i_data_bus[630]), .B2(n6182), .ZN(n5966) );
  AOI22D1BWP30P140LVT U6272 ( .A1(i_data_bus[566]), .A2(n6180), .B1(
        i_data_bus[598]), .B2(n6179), .ZN(n5965) );
  ND4D1BWP30P140LVT U6273 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), 
        .ZN(n5974) );
  AOI22D1BWP30P140LVT U6274 ( .A1(i_data_bus[950]), .A2(n6191), .B1(
        i_data_bus[374]), .B2(n6188), .ZN(n5972) );
  AOI22D1BWP30P140LVT U6275 ( .A1(i_data_bus[150]), .A2(n6190), .B1(
        i_data_bus[278]), .B2(n6143), .ZN(n5971) );
  AOI22D1BWP30P140LVT U6276 ( .A1(i_data_bus[918]), .A2(n5474), .B1(
        i_data_bus[438]), .B2(n5491), .ZN(n5970) );
  AOI22D1BWP30P140LVT U6277 ( .A1(i_data_bus[982]), .A2(n6161), .B1(
        i_data_bus[406]), .B2(n6192), .ZN(n5969) );
  ND4D1BWP30P140LVT U6278 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), 
        .ZN(n5973) );
  NR4D0BWP30P140LVT U6279 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), 
        .ZN(n5977) );
  ND4D1BWP30P140LVT U6280 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), 
        .ZN(o_data_bus[246]) );
  AOI22D1BWP30P140LVT U6281 ( .A1(i_data_bus[695]), .A2(n6158), .B1(
        i_data_bus[791]), .B2(n6165), .ZN(n6003) );
  AOI22D1BWP30P140LVT U6282 ( .A1(i_data_bus[119]), .A2(n6162), .B1(
        i_data_bus[855]), .B2(n6164), .ZN(n6002) );
  AOI22D1BWP30P140LVT U6283 ( .A1(i_data_bus[1015]), .A2(n6177), .B1(
        i_data_bus[951]), .B2(n6191), .ZN(n6001) );
  AOI22D1BWP30P140LVT U6284 ( .A1(i_data_bus[23]), .A2(n6169), .B1(
        i_data_bus[727]), .B2(n6167), .ZN(n5984) );
  AOI22D1BWP30P140LVT U6285 ( .A1(i_data_bus[759]), .A2(n6159), .B1(
        i_data_bus[663]), .B2(n6156), .ZN(n5983) );
  AOI22D1BWP30P140LVT U6286 ( .A1(i_data_bus[87]), .A2(n6163), .B1(
        i_data_bus[887]), .B2(n6168), .ZN(n5982) );
  AOI22D1BWP30P140LVT U6287 ( .A1(i_data_bus[55]), .A2(n6157), .B1(
        i_data_bus[823]), .B2(n6166), .ZN(n5981) );
  ND4D1BWP30P140LVT U6288 ( .A1(n5984), .A2(n5983), .A3(n5982), .A4(n5981), 
        .ZN(n5999) );
  OAI22D1BWP30P140LVT U6289 ( .A1(n5987), .A2(n5986), .B1(n5985), .B2(n6116), 
        .ZN(n5998) );
  AOI22D1BWP30P140LVT U6290 ( .A1(i_data_bus[183]), .A2(n5488), .B1(
        i_data_bus[503]), .B2(n6174), .ZN(n5991) );
  AOI22D1BWP30P140LVT U6291 ( .A1(i_data_bus[215]), .A2(n6189), .B1(
        i_data_bus[343]), .B2(n6178), .ZN(n5990) );
  AOI22D1BWP30P140LVT U6292 ( .A1(i_data_bus[631]), .A2(n6182), .B1(
        i_data_bus[599]), .B2(n6179), .ZN(n5989) );
  AOI22D1BWP30P140LVT U6293 ( .A1(i_data_bus[535]), .A2(n6181), .B1(
        i_data_bus[567]), .B2(n6180), .ZN(n5988) );
  ND4D1BWP30P140LVT U6294 ( .A1(n5991), .A2(n5990), .A3(n5989), .A4(n5988), 
        .ZN(n5997) );
  AOI22D1BWP30P140LVT U6295 ( .A1(i_data_bus[279]), .A2(n6143), .B1(
        i_data_bus[407]), .B2(n6192), .ZN(n5995) );
  AOI22D1BWP30P140LVT U6296 ( .A1(i_data_bus[247]), .A2(n6160), .B1(
        i_data_bus[311]), .B2(n6193), .ZN(n5994) );
  AOI22D1BWP30P140LVT U6297 ( .A1(i_data_bus[471]), .A2(n6187), .B1(
        i_data_bus[151]), .B2(n6190), .ZN(n5993) );
  AOI22D1BWP30P140LVT U6298 ( .A1(i_data_bus[983]), .A2(n6161), .B1(
        i_data_bus[919]), .B2(n5474), .ZN(n5992) );
  ND4D1BWP30P140LVT U6299 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), 
        .ZN(n5996) );
  NR4D0BWP30P140LVT U6300 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), 
        .ZN(n6000) );
  ND4D1BWP30P140LVT U6301 ( .A1(n6003), .A2(n6002), .A3(n6001), .A4(n6000), 
        .ZN(o_data_bus[247]) );
  AOI22D1BWP30P140LVT U6302 ( .A1(i_data_bus[120]), .A2(n6162), .B1(
        i_data_bus[696]), .B2(n6158), .ZN(n6024) );
  AOI22D1BWP30P140LVT U6303 ( .A1(i_data_bus[824]), .A2(n6166), .B1(
        i_data_bus[760]), .B2(n6159), .ZN(n6023) );
  AOI22D1BWP30P140LVT U6304 ( .A1(i_data_bus[344]), .A2(n6178), .B1(
        i_data_bus[376]), .B2(n6188), .ZN(n6022) );
  AOI22D1BWP30P140LVT U6305 ( .A1(i_data_bus[56]), .A2(n6157), .B1(
        i_data_bus[664]), .B2(n6156), .ZN(n6007) );
  AOI22D1BWP30P140LVT U6306 ( .A1(i_data_bus[856]), .A2(n6164), .B1(
        i_data_bus[728]), .B2(n6167), .ZN(n6006) );
  AOI22D1BWP30P140LVT U6307 ( .A1(i_data_bus[24]), .A2(n6169), .B1(
        i_data_bus[792]), .B2(n6165), .ZN(n6005) );
  AOI22D1BWP30P140LVT U6308 ( .A1(i_data_bus[88]), .A2(n6163), .B1(
        i_data_bus[888]), .B2(n6168), .ZN(n6004) );
  ND4D1BWP30P140LVT U6309 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), 
        .ZN(n6020) );
  MOAI22D1BWP30P140LVT U6310 ( .A1(n6008), .A2(n120), .B1(i_data_bus[152]), 
        .B2(n6190), .ZN(n6019) );
  AOI22D1BWP30P140LVT U6311 ( .A1(i_data_bus[1016]), .A2(n6177), .B1(
        i_data_bus[472]), .B2(n6187), .ZN(n6012) );
  AOI22D1BWP30P140LVT U6312 ( .A1(i_data_bus[248]), .A2(n6160), .B1(
        i_data_bus[312]), .B2(n6193), .ZN(n6011) );
  AOI22D1BWP30P140LVT U6313 ( .A1(i_data_bus[632]), .A2(n6182), .B1(
        i_data_bus[568]), .B2(n6180), .ZN(n6010) );
  AOI22D1BWP30P140LVT U6314 ( .A1(i_data_bus[600]), .A2(n6179), .B1(
        i_data_bus[536]), .B2(n6181), .ZN(n6009) );
  ND4D1BWP30P140LVT U6315 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), 
        .ZN(n6018) );
  AOI22D1BWP30P140LVT U6316 ( .A1(i_data_bus[216]), .A2(n6189), .B1(
        i_data_bus[504]), .B2(n6174), .ZN(n6016) );
  AOI22D1BWP30P140LVT U6317 ( .A1(i_data_bus[984]), .A2(n6161), .B1(
        i_data_bus[952]), .B2(n6191), .ZN(n6015) );
  AOI22D1BWP30P140LVT U6318 ( .A1(i_data_bus[920]), .A2(n5474), .B1(
        i_data_bus[184]), .B2(n5488), .ZN(n6014) );
  AOI22D1BWP30P140LVT U6319 ( .A1(i_data_bus[408]), .A2(n6192), .B1(
        i_data_bus[440]), .B2(n5491), .ZN(n6013) );
  ND4D1BWP30P140LVT U6320 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), 
        .ZN(n6017) );
  NR4D0BWP30P140LVT U6321 ( .A1(n6020), .A2(n6019), .A3(n6018), .A4(n6017), 
        .ZN(n6021) );
  ND4D1BWP30P140LVT U6322 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), 
        .ZN(o_data_bus[248]) );
  AOI22D1BWP30P140LVT U6323 ( .A1(i_data_bus[761]), .A2(n6159), .B1(
        i_data_bus[889]), .B2(n6168), .ZN(n6045) );
  AOI22D1BWP30P140LVT U6324 ( .A1(i_data_bus[57]), .A2(n6157), .B1(
        i_data_bus[121]), .B2(n6162), .ZN(n6044) );
  AOI22D1BWP30P140LVT U6325 ( .A1(i_data_bus[377]), .A2(n6188), .B1(
        i_data_bus[313]), .B2(n6193), .ZN(n6043) );
  AOI22D1BWP30P140LVT U6326 ( .A1(i_data_bus[665]), .A2(n6156), .B1(
        i_data_bus[793]), .B2(n6165), .ZN(n6028) );
  AOI22D1BWP30P140LVT U6327 ( .A1(i_data_bus[825]), .A2(n6166), .B1(
        i_data_bus[857]), .B2(n6164), .ZN(n6027) );
  AOI22D1BWP30P140LVT U6328 ( .A1(i_data_bus[729]), .A2(n6167), .B1(
        i_data_bus[697]), .B2(n6158), .ZN(n6026) );
  AOI22D1BWP30P140LVT U6329 ( .A1(i_data_bus[25]), .A2(n6169), .B1(
        i_data_bus[89]), .B2(n6163), .ZN(n6025) );
  ND4D1BWP30P140LVT U6330 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), 
        .ZN(n6041) );
  MOAI22D1BWP30P140LVT U6331 ( .A1(n6029), .A2(n119), .B1(i_data_bus[1017]), 
        .B2(n6177), .ZN(n6040) );
  AOI22D1BWP30P140LVT U6332 ( .A1(i_data_bus[921]), .A2(n5474), .B1(
        i_data_bus[985]), .B2(n6161), .ZN(n6033) );
  AOI22D1BWP30P140LVT U6333 ( .A1(i_data_bus[153]), .A2(n6190), .B1(
        i_data_bus[217]), .B2(n6189), .ZN(n6032) );
  AOI22D1BWP30P140LVT U6334 ( .A1(i_data_bus[569]), .A2(n6180), .B1(
        i_data_bus[537]), .B2(n6181), .ZN(n6031) );
  AOI22D1BWP30P140LVT U6335 ( .A1(i_data_bus[633]), .A2(n6182), .B1(
        i_data_bus[601]), .B2(n6179), .ZN(n6030) );
  ND4D1BWP30P140LVT U6336 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), 
        .ZN(n6039) );
  AOI22D1BWP30P140LVT U6337 ( .A1(i_data_bus[345]), .A2(n6178), .B1(
        i_data_bus[281]), .B2(n6143), .ZN(n6037) );
  AOI22D1BWP30P140LVT U6338 ( .A1(i_data_bus[185]), .A2(n5488), .B1(
        i_data_bus[441]), .B2(n5491), .ZN(n6036) );
  AOI22D1BWP30P140LVT U6339 ( .A1(i_data_bus[473]), .A2(n6187), .B1(
        i_data_bus[505]), .B2(n6174), .ZN(n6035) );
  AOI22D1BWP30P140LVT U6340 ( .A1(i_data_bus[953]), .A2(n6191), .B1(
        i_data_bus[249]), .B2(n6160), .ZN(n6034) );
  ND4D1BWP30P140LVT U6341 ( .A1(n6037), .A2(n6036), .A3(n6035), .A4(n6034), 
        .ZN(n6038) );
  NR4D0BWP30P140LVT U6342 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), 
        .ZN(n6042) );
  ND4D1BWP30P140LVT U6343 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), 
        .ZN(o_data_bus[249]) );
  AOI22D1BWP30P140LVT U6344 ( .A1(i_data_bus[90]), .A2(n6163), .B1(
        i_data_bus[730]), .B2(n6167), .ZN(n6066) );
  AOI22D1BWP30P140LVT U6345 ( .A1(i_data_bus[698]), .A2(n6158), .B1(
        i_data_bus[794]), .B2(n6165), .ZN(n6065) );
  AOI22D1BWP30P140LVT U6346 ( .A1(i_data_bus[1018]), .A2(n6177), .B1(
        i_data_bus[314]), .B2(n6193), .ZN(n6064) );
  AOI22D1BWP30P140LVT U6347 ( .A1(i_data_bus[58]), .A2(n6157), .B1(
        i_data_bus[826]), .B2(n6166), .ZN(n6049) );
  AOI22D1BWP30P140LVT U6348 ( .A1(i_data_bus[890]), .A2(n6168), .B1(
        i_data_bus[858]), .B2(n6164), .ZN(n6048) );
  AOI22D1BWP30P140LVT U6349 ( .A1(i_data_bus[122]), .A2(n6162), .B1(
        i_data_bus[666]), .B2(n6156), .ZN(n6047) );
  AOI22D1BWP30P140LVT U6350 ( .A1(i_data_bus[26]), .A2(n6169), .B1(
        i_data_bus[762]), .B2(n6159), .ZN(n6046) );
  ND4D1BWP30P140LVT U6351 ( .A1(n6049), .A2(n6048), .A3(n6047), .A4(n6046), 
        .ZN(n6062) );
  MOAI22D1BWP30P140LVT U6352 ( .A1(n6050), .A2(n6116), .B1(i_data_bus[250]), 
        .B2(n6160), .ZN(n6061) );
  AOI22D1BWP30P140LVT U6353 ( .A1(i_data_bus[954]), .A2(n6191), .B1(
        i_data_bus[282]), .B2(n6143), .ZN(n6054) );
  AOI22D1BWP30P140LVT U6354 ( .A1(i_data_bus[346]), .A2(n6178), .B1(
        i_data_bus[186]), .B2(n5488), .ZN(n6053) );
  AOI22D1BWP30P140LVT U6355 ( .A1(i_data_bus[538]), .A2(n6181), .B1(
        i_data_bus[570]), .B2(n6180), .ZN(n6052) );
  AOI22D1BWP30P140LVT U6356 ( .A1(i_data_bus[602]), .A2(n6179), .B1(
        i_data_bus[634]), .B2(n6182), .ZN(n6051) );
  ND4D1BWP30P140LVT U6357 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), 
        .ZN(n6060) );
  AOI22D1BWP30P140LVT U6358 ( .A1(i_data_bus[922]), .A2(n5474), .B1(
        i_data_bus[506]), .B2(n6174), .ZN(n6058) );
  AOI22D1BWP30P140LVT U6359 ( .A1(i_data_bus[154]), .A2(n6190), .B1(
        i_data_bus[474]), .B2(n6187), .ZN(n6057) );
  AOI22D1BWP30P140LVT U6360 ( .A1(i_data_bus[986]), .A2(n6161), .B1(
        i_data_bus[410]), .B2(n6192), .ZN(n6056) );
  AOI22D1BWP30P140LVT U6361 ( .A1(i_data_bus[442]), .A2(n5491), .B1(
        i_data_bus[218]), .B2(n6189), .ZN(n6055) );
  ND4D1BWP30P140LVT U6362 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), 
        .ZN(n6059) );
  NR4D0BWP30P140LVT U6363 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), 
        .ZN(n6063) );
  ND4D1BWP30P140LVT U6364 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), 
        .ZN(o_data_bus[250]) );
  AOI22D1BWP30P140LVT U6365 ( .A1(i_data_bus[59]), .A2(n6157), .B1(
        i_data_bus[827]), .B2(n6166), .ZN(n6088) );
  AOI22D1BWP30P140LVT U6366 ( .A1(i_data_bus[123]), .A2(n6162), .B1(
        i_data_bus[859]), .B2(n6164), .ZN(n6087) );
  AOI22D1BWP30P140LVT U6367 ( .A1(i_data_bus[507]), .A2(n6174), .B1(
        i_data_bus[155]), .B2(n6190), .ZN(n6086) );
  AOI22D1BWP30P140LVT U6368 ( .A1(i_data_bus[91]), .A2(n6163), .B1(
        i_data_bus[731]), .B2(n6167), .ZN(n6070) );
  AOI22D1BWP30P140LVT U6369 ( .A1(i_data_bus[667]), .A2(n6156), .B1(
        i_data_bus[699]), .B2(n6158), .ZN(n6069) );
  AOI22D1BWP30P140LVT U6370 ( .A1(i_data_bus[27]), .A2(n6169), .B1(
        i_data_bus[795]), .B2(n6165), .ZN(n6068) );
  AOI22D1BWP30P140LVT U6371 ( .A1(i_data_bus[891]), .A2(n6168), .B1(
        i_data_bus[763]), .B2(n6159), .ZN(n6067) );
  ND4D1BWP30P140LVT U6372 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), 
        .ZN(n6084) );
  OAI22D1BWP30P140LVT U6373 ( .A1(n6072), .A2(n6094), .B1(n6071), .B2(n6175), 
        .ZN(n6083) );
  AOI22D1BWP30P140LVT U6374 ( .A1(i_data_bus[219]), .A2(n6189), .B1(
        i_data_bus[283]), .B2(n6143), .ZN(n6076) );
  AOI22D1BWP30P140LVT U6375 ( .A1(i_data_bus[1019]), .A2(n6177), .B1(
        i_data_bus[379]), .B2(n6188), .ZN(n6075) );
  AOI22D1BWP30P140LVT U6376 ( .A1(i_data_bus[571]), .A2(n6180), .B1(
        i_data_bus[539]), .B2(n6181), .ZN(n6074) );
  AOI22D1BWP30P140LVT U6377 ( .A1(i_data_bus[603]), .A2(n6179), .B1(
        i_data_bus[635]), .B2(n6182), .ZN(n6073) );
  ND4D1BWP30P140LVT U6378 ( .A1(n6076), .A2(n6075), .A3(n6074), .A4(n6073), 
        .ZN(n6082) );
  AOI22D1BWP30P140LVT U6379 ( .A1(i_data_bus[315]), .A2(n6193), .B1(
        i_data_bus[475]), .B2(n6187), .ZN(n6080) );
  AOI22D1BWP30P140LVT U6380 ( .A1(i_data_bus[987]), .A2(n6161), .B1(
        i_data_bus[443]), .B2(n5491), .ZN(n6079) );
  AOI22D1BWP30P140LVT U6381 ( .A1(i_data_bus[411]), .A2(n6192), .B1(
        i_data_bus[251]), .B2(n6160), .ZN(n6078) );
  AOI22D1BWP30P140LVT U6382 ( .A1(i_data_bus[923]), .A2(n5474), .B1(
        i_data_bus[955]), .B2(n6191), .ZN(n6077) );
  ND4D1BWP30P140LVT U6383 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), 
        .ZN(n6081) );
  NR4D0BWP30P140LVT U6384 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), 
        .ZN(n6085) );
  ND4D1BWP30P140LVT U6385 ( .A1(n6088), .A2(n6087), .A3(n6086), .A4(n6085), 
        .ZN(o_data_bus[251]) );
  AOI22D1BWP30P140LVT U6386 ( .A1(i_data_bus[124]), .A2(n6162), .B1(
        i_data_bus[860]), .B2(n6164), .ZN(n6111) );
  AOI22D1BWP30P140LVT U6387 ( .A1(i_data_bus[92]), .A2(n6163), .B1(
        i_data_bus[668]), .B2(n6156), .ZN(n6110) );
  AOI22D1BWP30P140LVT U6388 ( .A1(i_data_bus[988]), .A2(n6161), .B1(
        i_data_bus[284]), .B2(n6143), .ZN(n6109) );
  AOI22D1BWP30P140LVT U6389 ( .A1(i_data_bus[28]), .A2(n6169), .B1(
        i_data_bus[732]), .B2(n6167), .ZN(n6092) );
  AOI22D1BWP30P140LVT U6390 ( .A1(i_data_bus[828]), .A2(n6166), .B1(
        i_data_bus[700]), .B2(n6158), .ZN(n6091) );
  AOI22D1BWP30P140LVT U6391 ( .A1(i_data_bus[796]), .A2(n6165), .B1(
        i_data_bus[764]), .B2(n6159), .ZN(n6090) );
  AOI22D1BWP30P140LVT U6392 ( .A1(i_data_bus[60]), .A2(n6157), .B1(
        i_data_bus[892]), .B2(n6168), .ZN(n6089) );
  ND4D1BWP30P140LVT U6393 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), 
        .ZN(n6107) );
  OAI22D1BWP30P140LVT U6394 ( .A1(n6095), .A2(n6094), .B1(n6093), .B2(n119), 
        .ZN(n6106) );
  AOI22D1BWP30P140LVT U6395 ( .A1(i_data_bus[924]), .A2(n5474), .B1(
        i_data_bus[444]), .B2(n5491), .ZN(n6099) );
  AOI22D1BWP30P140LVT U6396 ( .A1(i_data_bus[380]), .A2(n6188), .B1(
        i_data_bus[220]), .B2(n6189), .ZN(n6098) );
  AOI22D1BWP30P140LVT U6397 ( .A1(i_data_bus[636]), .A2(n6182), .B1(
        i_data_bus[604]), .B2(n6179), .ZN(n6097) );
  AOI22D1BWP30P140LVT U6398 ( .A1(i_data_bus[540]), .A2(n6181), .B1(
        i_data_bus[572]), .B2(n6180), .ZN(n6096) );
  ND4D1BWP30P140LVT U6399 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), 
        .ZN(n6105) );
  AOI22D1BWP30P140LVT U6400 ( .A1(i_data_bus[956]), .A2(n6191), .B1(
        i_data_bus[316]), .B2(n6193), .ZN(n6103) );
  AOI22D1BWP30P140LVT U6401 ( .A1(i_data_bus[1020]), .A2(n6177), .B1(
        i_data_bus[156]), .B2(n6190), .ZN(n6102) );
  AOI22D1BWP30P140LVT U6402 ( .A1(i_data_bus[188]), .A2(n5488), .B1(
        i_data_bus[476]), .B2(n6187), .ZN(n6101) );
  AOI22D1BWP30P140LVT U6403 ( .A1(i_data_bus[252]), .A2(n6160), .B1(
        i_data_bus[508]), .B2(n6174), .ZN(n6100) );
  ND4D1BWP30P140LVT U6404 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), 
        .ZN(n6104) );
  NR4D0BWP30P140LVT U6405 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), 
        .ZN(n6108) );
  ND4D1BWP30P140LVT U6406 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), 
        .ZN(o_data_bus[252]) );
  AOI22D1BWP30P140LVT U6407 ( .A1(i_data_bus[765]), .A2(n6159), .B1(
        i_data_bus[797]), .B2(n6165), .ZN(n6133) );
  AOI22D1BWP30P140LVT U6408 ( .A1(i_data_bus[669]), .A2(n6156), .B1(
        i_data_bus[829]), .B2(n6166), .ZN(n6132) );
  AOI22D1BWP30P140LVT U6409 ( .A1(i_data_bus[349]), .A2(n6178), .B1(
        i_data_bus[285]), .B2(n6143), .ZN(n6131) );
  AOI22D1BWP30P140LVT U6410 ( .A1(i_data_bus[29]), .A2(n6169), .B1(
        i_data_bus[125]), .B2(n6162), .ZN(n6115) );
  AOI22D1BWP30P140LVT U6411 ( .A1(i_data_bus[61]), .A2(n6157), .B1(
        i_data_bus[893]), .B2(n6168), .ZN(n6114) );
  AOI22D1BWP30P140LVT U6412 ( .A1(i_data_bus[93]), .A2(n6163), .B1(
        i_data_bus[861]), .B2(n6164), .ZN(n6113) );
  AOI22D1BWP30P140LVT U6413 ( .A1(i_data_bus[701]), .A2(n6158), .B1(
        i_data_bus[733]), .B2(n6167), .ZN(n6112) );
  ND4D1BWP30P140LVT U6414 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), 
        .ZN(n6129) );
  MOAI22D1BWP30P140LVT U6415 ( .A1(n6117), .A2(n6116), .B1(i_data_bus[157]), 
        .B2(n6190), .ZN(n6128) );
  AOI22D1BWP30P140LVT U6416 ( .A1(i_data_bus[925]), .A2(n5474), .B1(
        i_data_bus[957]), .B2(n6191), .ZN(n6121) );
  AOI22D1BWP30P140LVT U6417 ( .A1(i_data_bus[989]), .A2(n6161), .B1(
        i_data_bus[413]), .B2(n6192), .ZN(n6120) );
  AOI22D1BWP30P140LVT U6418 ( .A1(i_data_bus[573]), .A2(n6180), .B1(
        i_data_bus[541]), .B2(n6181), .ZN(n6119) );
  AOI22D1BWP30P140LVT U6419 ( .A1(i_data_bus[637]), .A2(n6182), .B1(
        i_data_bus[605]), .B2(n6179), .ZN(n6118) );
  ND4D1BWP30P140LVT U6420 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), 
        .ZN(n6127) );
  AOI22D1BWP30P140LVT U6421 ( .A1(i_data_bus[1021]), .A2(n6177), .B1(
        i_data_bus[221]), .B2(n6189), .ZN(n6125) );
  AOI22D1BWP30P140LVT U6422 ( .A1(i_data_bus[445]), .A2(n5491), .B1(
        i_data_bus[253]), .B2(n6160), .ZN(n6124) );
  AOI22D1BWP30P140LVT U6423 ( .A1(i_data_bus[317]), .A2(n6193), .B1(
        i_data_bus[509]), .B2(n6174), .ZN(n6123) );
  AOI22D1BWP30P140LVT U6424 ( .A1(i_data_bus[189]), .A2(n5488), .B1(
        i_data_bus[477]), .B2(n6187), .ZN(n6122) );
  ND4D1BWP30P140LVT U6425 ( .A1(n6125), .A2(n6124), .A3(n6123), .A4(n6122), 
        .ZN(n6126) );
  NR4D0BWP30P140LVT U6426 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), 
        .ZN(n6130) );
  ND4D1BWP30P140LVT U6427 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), 
        .ZN(o_data_bus[253]) );
  AOI22D1BWP30P140LVT U6428 ( .A1(i_data_bus[94]), .A2(n6163), .B1(
        i_data_bus[702]), .B2(n6158), .ZN(n6155) );
  AOI22D1BWP30P140LVT U6429 ( .A1(i_data_bus[62]), .A2(n6157), .B1(
        i_data_bus[126]), .B2(n6162), .ZN(n6154) );
  AOI22D1BWP30P140LVT U6430 ( .A1(i_data_bus[958]), .A2(n6191), .B1(
        i_data_bus[478]), .B2(n6187), .ZN(n6153) );
  AOI22D1BWP30P140LVT U6431 ( .A1(i_data_bus[862]), .A2(n6164), .B1(
        i_data_bus[734]), .B2(n6167), .ZN(n6137) );
  AOI22D1BWP30P140LVT U6432 ( .A1(i_data_bus[30]), .A2(n6169), .B1(
        i_data_bus[798]), .B2(n6165), .ZN(n6136) );
  AOI22D1BWP30P140LVT U6433 ( .A1(i_data_bus[670]), .A2(n6156), .B1(
        i_data_bus[830]), .B2(n6166), .ZN(n6135) );
  AOI22D1BWP30P140LVT U6434 ( .A1(i_data_bus[766]), .A2(n6159), .B1(
        i_data_bus[894]), .B2(n6168), .ZN(n6134) );
  ND4D1BWP30P140LVT U6435 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), 
        .ZN(n6151) );
  MOAI22D1BWP30P140LVT U6436 ( .A1(n6138), .A2(n119), .B1(i_data_bus[990]), 
        .B2(n6161), .ZN(n6150) );
  AOI22D1BWP30P140LVT U6437 ( .A1(i_data_bus[222]), .A2(n6189), .B1(
        i_data_bus[382]), .B2(n6188), .ZN(n6142) );
  AOI22D1BWP30P140LVT U6438 ( .A1(i_data_bus[1022]), .A2(n6177), .B1(
        i_data_bus[446]), .B2(n5491), .ZN(n6141) );
  AOI22D1BWP30P140LVT U6439 ( .A1(i_data_bus[542]), .A2(n6181), .B1(
        i_data_bus[606]), .B2(n6179), .ZN(n6140) );
  AOI22D1BWP30P140LVT U6440 ( .A1(i_data_bus[574]), .A2(n6180), .B1(
        i_data_bus[638]), .B2(n6182), .ZN(n6139) );
  ND4D1BWP30P140LVT U6441 ( .A1(n6142), .A2(n6141), .A3(n6140), .A4(n6139), 
        .ZN(n6149) );
  AOI22D1BWP30P140LVT U6442 ( .A1(i_data_bus[926]), .A2(n5474), .B1(
        i_data_bus[286]), .B2(n6143), .ZN(n6147) );
  AOI22D1BWP30P140LVT U6443 ( .A1(i_data_bus[318]), .A2(n6193), .B1(
        i_data_bus[190]), .B2(n5488), .ZN(n6146) );
  AOI22D1BWP30P140LVT U6444 ( .A1(i_data_bus[254]), .A2(n6160), .B1(
        i_data_bus[158]), .B2(n6190), .ZN(n6145) );
  AOI22D1BWP30P140LVT U6445 ( .A1(i_data_bus[350]), .A2(n6178), .B1(
        i_data_bus[510]), .B2(n6174), .ZN(n6144) );
  ND4D1BWP30P140LVT U6446 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), 
        .ZN(n6148) );
  NR4D0BWP30P140LVT U6447 ( .A1(n6151), .A2(n6150), .A3(n6149), .A4(n6148), 
        .ZN(n6152) );
  ND4D1BWP30P140LVT U6448 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), 
        .ZN(o_data_bus[254]) );
  AOI22D1BWP30P140LVT U6449 ( .A1(i_data_bus[63]), .A2(n6157), .B1(
        i_data_bus[671]), .B2(n6156), .ZN(n6205) );
  AOI22D1BWP30P140LVT U6450 ( .A1(i_data_bus[767]), .A2(n6159), .B1(
        i_data_bus[703]), .B2(n6158), .ZN(n6204) );
  AOI22D1BWP30P140LVT U6451 ( .A1(i_data_bus[991]), .A2(n6161), .B1(
        i_data_bus[255]), .B2(n6160), .ZN(n6203) );
  AOI22D1BWP30P140LVT U6452 ( .A1(i_data_bus[95]), .A2(n6163), .B1(
        i_data_bus[127]), .B2(n6162), .ZN(n6173) );
  AOI22D1BWP30P140LVT U6453 ( .A1(i_data_bus[799]), .A2(n6165), .B1(
        i_data_bus[863]), .B2(n6164), .ZN(n6172) );
  AOI22D1BWP30P140LVT U6454 ( .A1(i_data_bus[735]), .A2(n6167), .B1(
        i_data_bus[831]), .B2(n6166), .ZN(n6171) );
  AOI22D1BWP30P140LVT U6455 ( .A1(i_data_bus[31]), .A2(n6169), .B1(
        i_data_bus[895]), .B2(n6168), .ZN(n6170) );
  ND4D1BWP30P140LVT U6456 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), 
        .ZN(n6201) );
  MOAI22D1BWP30P140LVT U6457 ( .A1(n6176), .A2(n6175), .B1(i_data_bus[511]), 
        .B2(n6174), .ZN(n6200) );
  AOI22D1BWP30P140LVT U6458 ( .A1(i_data_bus[1023]), .A2(n6177), .B1(
        i_data_bus[287]), .B2(n6143), .ZN(n6186) );
  AOI22D1BWP30P140LVT U6459 ( .A1(i_data_bus[927]), .A2(n5474), .B1(
        i_data_bus[351]), .B2(n6178), .ZN(n6185) );
  AOI22D1BWP30P140LVT U6460 ( .A1(i_data_bus[575]), .A2(n6180), .B1(
        i_data_bus[607]), .B2(n6179), .ZN(n6184) );
  AOI22D1BWP30P140LVT U6461 ( .A1(i_data_bus[639]), .A2(n6182), .B1(
        i_data_bus[543]), .B2(n6181), .ZN(n6183) );
  ND4D1BWP30P140LVT U6462 ( .A1(n6186), .A2(n6185), .A3(n6184), .A4(n6183), 
        .ZN(n6199) );
  AOI22D1BWP30P140LVT U6463 ( .A1(i_data_bus[447]), .A2(n5491), .B1(
        i_data_bus[479]), .B2(n6187), .ZN(n6197) );
  AOI22D1BWP30P140LVT U6464 ( .A1(i_data_bus[223]), .A2(n6189), .B1(
        i_data_bus[383]), .B2(n6188), .ZN(n6196) );
  AOI22D1BWP30P140LVT U6465 ( .A1(i_data_bus[959]), .A2(n6191), .B1(
        i_data_bus[159]), .B2(n6190), .ZN(n6195) );
  AOI22D1BWP30P140LVT U6466 ( .A1(i_data_bus[319]), .A2(n6193), .B1(
        i_data_bus[415]), .B2(n6192), .ZN(n6194) );
  ND4D1BWP30P140LVT U6467 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), 
        .ZN(n6198) );
  NR4D0BWP30P140LVT U6468 ( .A1(n6201), .A2(n6200), .A3(n6199), .A4(n6198), 
        .ZN(n6202) );
  ND4D1BWP30P140LVT U6469 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), 
        .ZN(o_data_bus[255]) );
endmodule


module crossbar_one_hot_comb_wrapper_seq ( clk, rst, i_valid, i_data_bus, 
        o_valid, o_data_bus, i_en, i_cmd );
  input [31:0] i_valid;
  input [1023:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [255:0] i_cmd;
  input clk, rst, i_en;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N61, N62, N63, N64, N65, N66, N67, N103, N104, N105, N106, N107, N108,
         N109, N110, N115, N116, N117, N118, N119, N127, N128, N129, N130,
         N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141,
         N142, N143, N144, N145, N151, N152, N153, N154, N155, N156, N157,
         N158, N159, N160, N161, N162, N175, N176, N177, N178, N179, N180,
         N181, N182, N187, N188, N189, N190, N191, N247, N248, N249, N250,
         N251, N252, N253, N254, N259, N260, N261, N262, N263, N319, N320,
         N321, N322, N323, N324, N325, N326, N331, N332, N333, N334, N335,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617,
         N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628,
         N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639,
         N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650,
         N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661,
         N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672,
         N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683,
         N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694,
         N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705,
         N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716,
         N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727,
         N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738,
         N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749,
         N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760,
         N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771,
         N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782,
         N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793,
         N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804,
         N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815,
         N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826,
         N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837,
         N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848,
         N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859,
         N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870,
         N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881,
         N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892,
         N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903,
         N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914,
         N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925,
         N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936,
         N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947,
         N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958,
         N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969,
         N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980,
         N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991,
         N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002,
         N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012,
         N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022,
         N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032,
         N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042,
         N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052,
         N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062,
         N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072,
         N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082,
         N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092,
         N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102,
         N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112,
         N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122,
         N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132,
         N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142,
         N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152,
         N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162,
         N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172,
         N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182,
         N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192,
         N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202,
         N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212,
         N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222,
         N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232,
         N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242,
         N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252,
         N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262,
         N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272,
         N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282,
         N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292,
         N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302,
         N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312,
         N1313, N1314, n7, n8, n9, n10, n11, n12, n13, n14, n15;
  wire   [31:0] i_valid_reg;
  wire   [1023:0] i_data_bus_reg;
  wire   [255:0] i_cmd_reg;
  wire   [7:0] o_valid_wire;
  wire   [255:0] o_data_bus_wire;

  crossbar_one_hot_comb_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA32 dut ( 
        .i_valid(i_valid_reg), .i_data_bus(i_data_bus_reg), .o_valid(
        o_valid_wire), .o_data_bus(o_data_bus_wire), .i_en(i_en), .i_cmd(
        i_cmd_reg) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_255_ ( .D(N1314), .CP(clk), .Q(
        i_cmd_reg[255]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_254_ ( .D(N1313), .CP(clk), .Q(
        i_cmd_reg[254]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_253_ ( .D(N1312), .CP(clk), .Q(
        i_cmd_reg[253]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_252_ ( .D(N1311), .CP(clk), .Q(
        i_cmd_reg[252]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_251_ ( .D(N1310), .CP(clk), .Q(
        i_cmd_reg[251]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_250_ ( .D(N1309), .CP(clk), .Q(
        i_cmd_reg[250]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_249_ ( .D(N1308), .CP(clk), .Q(
        i_cmd_reg[249]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_248_ ( .D(N1307), .CP(clk), .Q(
        i_cmd_reg[248]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_247_ ( .D(N1306), .CP(clk), .Q(
        i_cmd_reg[247]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_246_ ( .D(N1305), .CP(clk), .Q(
        i_cmd_reg[246]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_245_ ( .D(N1304), .CP(clk), .Q(
        i_cmd_reg[245]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_244_ ( .D(N1303), .CP(clk), .Q(
        i_cmd_reg[244]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_243_ ( .D(N1302), .CP(clk), .Q(
        i_cmd_reg[243]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_242_ ( .D(N1301), .CP(clk), .Q(
        i_cmd_reg[242]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_241_ ( .D(N1300), .CP(clk), .Q(
        i_cmd_reg[241]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_240_ ( .D(N1299), .CP(clk), .Q(
        i_cmd_reg[240]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_239_ ( .D(N1298), .CP(clk), .Q(
        i_cmd_reg[239]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_238_ ( .D(N1297), .CP(clk), .Q(
        i_cmd_reg[238]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_237_ ( .D(N1296), .CP(clk), .Q(
        i_cmd_reg[237]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_236_ ( .D(N1295), .CP(clk), .Q(
        i_cmd_reg[236]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_235_ ( .D(N1294), .CP(clk), .Q(
        i_cmd_reg[235]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_234_ ( .D(N1293), .CP(clk), .Q(
        i_cmd_reg[234]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_233_ ( .D(N1292), .CP(clk), .Q(
        i_cmd_reg[233]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_232_ ( .D(N1291), .CP(clk), .Q(
        i_cmd_reg[232]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_231_ ( .D(N1290), .CP(clk), .Q(
        i_cmd_reg[231]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_230_ ( .D(N1289), .CP(clk), .Q(
        i_cmd_reg[230]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_229_ ( .D(N1288), .CP(clk), .Q(
        i_cmd_reg[229]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_228_ ( .D(N1287), .CP(clk), .Q(
        i_cmd_reg[228]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_227_ ( .D(N1286), .CP(clk), .Q(
        i_cmd_reg[227]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_226_ ( .D(N1285), .CP(clk), .Q(
        i_cmd_reg[226]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_225_ ( .D(N1284), .CP(clk), .Q(
        i_cmd_reg[225]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_224_ ( .D(N1283), .CP(clk), .Q(
        i_cmd_reg[224]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_223_ ( .D(N1282), .CP(clk), .Q(
        i_cmd_reg[223]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_222_ ( .D(N1281), .CP(clk), .Q(
        i_cmd_reg[222]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_220_ ( .D(N1279), .CP(clk), .Q(
        i_cmd_reg[220]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_219_ ( .D(N1278), .CP(clk), .Q(
        i_cmd_reg[219]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_218_ ( .D(N1277), .CP(clk), .Q(
        i_cmd_reg[218]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_217_ ( .D(N1276), .CP(clk), .Q(
        i_cmd_reg[217]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_216_ ( .D(N1275), .CP(clk), .Q(
        i_cmd_reg[216]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_215_ ( .D(N1274), .CP(clk), .Q(
        i_cmd_reg[215]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_214_ ( .D(N1273), .CP(clk), .Q(
        i_cmd_reg[214]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_213_ ( .D(N1272), .CP(clk), .Q(
        i_cmd_reg[213]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_212_ ( .D(N1271), .CP(clk), .Q(
        i_cmd_reg[212]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_211_ ( .D(N1270), .CP(clk), .Q(
        i_cmd_reg[211]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_210_ ( .D(N1269), .CP(clk), .Q(
        i_cmd_reg[210]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_209_ ( .D(N1268), .CP(clk), .Q(
        i_cmd_reg[209]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_208_ ( .D(N1267), .CP(clk), .Q(
        i_cmd_reg[208]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_207_ ( .D(N1266), .CP(clk), .Q(
        i_cmd_reg[207]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_206_ ( .D(N1265), .CP(clk), .Q(
        i_cmd_reg[206]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_205_ ( .D(N1264), .CP(clk), .Q(
        i_cmd_reg[205]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_204_ ( .D(N1263), .CP(clk), .Q(
        i_cmd_reg[204]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_203_ ( .D(N1262), .CP(clk), .Q(
        i_cmd_reg[203]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_202_ ( .D(N1261), .CP(clk), .Q(
        i_cmd_reg[202]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_201_ ( .D(N1260), .CP(clk), .Q(
        i_cmd_reg[201]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_200_ ( .D(N1259), .CP(clk), .Q(
        i_cmd_reg[200]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_199_ ( .D(N1258), .CP(clk), .Q(
        i_cmd_reg[199]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_198_ ( .D(N1257), .CP(clk), .Q(
        i_cmd_reg[198]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_197_ ( .D(N1256), .CP(clk), .Q(
        i_cmd_reg[197]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_196_ ( .D(N1255), .CP(clk), .Q(
        i_cmd_reg[196]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_195_ ( .D(N1254), .CP(clk), .Q(
        i_cmd_reg[195]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_194_ ( .D(N1253), .CP(clk), .Q(
        i_cmd_reg[194]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_193_ ( .D(N1252), .CP(clk), .Q(
        i_cmd_reg[193]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_192_ ( .D(N1251), .CP(clk), .Q(
        i_cmd_reg[192]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_191_ ( .D(N1250), .CP(clk), .Q(
        i_cmd_reg[191]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_190_ ( .D(N1249), .CP(clk), .Q(
        i_cmd_reg[190]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_189_ ( .D(N1248), .CP(clk), .Q(
        i_cmd_reg[189]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_188_ ( .D(N1247), .CP(clk), .Q(
        i_cmd_reg[188]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_187_ ( .D(N1246), .CP(clk), .Q(
        i_cmd_reg[187]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_186_ ( .D(N1245), .CP(clk), .Q(
        i_cmd_reg[186]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_185_ ( .D(N1244), .CP(clk), .Q(
        i_cmd_reg[185]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_184_ ( .D(N1243), .CP(clk), .Q(
        i_cmd_reg[184]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_183_ ( .D(N1242), .CP(clk), .Q(
        i_cmd_reg[183]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_182_ ( .D(N1241), .CP(clk), .Q(
        i_cmd_reg[182]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_181_ ( .D(N1240), .CP(clk), .Q(
        i_cmd_reg[181]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_180_ ( .D(N1239), .CP(clk), .Q(
        i_cmd_reg[180]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_179_ ( .D(N1238), .CP(clk), .Q(
        i_cmd_reg[179]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_178_ ( .D(N1237), .CP(clk), .Q(
        i_cmd_reg[178]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_177_ ( .D(N1236), .CP(clk), .Q(
        i_cmd_reg[177]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_176_ ( .D(N1235), .CP(clk), .Q(
        i_cmd_reg[176]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_175_ ( .D(N1234), .CP(clk), .Q(
        i_cmd_reg[175]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_174_ ( .D(N1233), .CP(clk), .Q(
        i_cmd_reg[174]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_173_ ( .D(N1232), .CP(clk), .Q(
        i_cmd_reg[173]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_172_ ( .D(N1231), .CP(clk), .Q(
        i_cmd_reg[172]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_171_ ( .D(N1230), .CP(clk), .Q(
        i_cmd_reg[171]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_170_ ( .D(N1229), .CP(clk), .Q(
        i_cmd_reg[170]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_169_ ( .D(N1228), .CP(clk), .Q(
        i_cmd_reg[169]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_168_ ( .D(N1227), .CP(clk), .Q(
        i_cmd_reg[168]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_167_ ( .D(N1226), .CP(clk), .Q(
        i_cmd_reg[167]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_166_ ( .D(N1225), .CP(clk), .Q(
        i_cmd_reg[166]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_165_ ( .D(N1224), .CP(clk), .Q(
        i_cmd_reg[165]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_164_ ( .D(N1223), .CP(clk), .Q(
        i_cmd_reg[164]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_163_ ( .D(N1222), .CP(clk), .Q(
        i_cmd_reg[163]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_162_ ( .D(N1221), .CP(clk), .Q(
        i_cmd_reg[162]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_161_ ( .D(N1220), .CP(clk), .Q(
        i_cmd_reg[161]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_160_ ( .D(N1219), .CP(clk), .Q(
        i_cmd_reg[160]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_159_ ( .D(N1218), .CP(clk), .Q(
        i_cmd_reg[159]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_158_ ( .D(N1217), .CP(clk), .Q(
        i_cmd_reg[158]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_157_ ( .D(N1216), .CP(clk), .Q(
        i_cmd_reg[157]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_156_ ( .D(N1215), .CP(clk), .Q(
        i_cmd_reg[156]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_155_ ( .D(N1214), .CP(clk), .Q(
        i_cmd_reg[155]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_154_ ( .D(N1213), .CP(clk), .Q(
        i_cmd_reg[154]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_153_ ( .D(N1212), .CP(clk), .Q(
        i_cmd_reg[153]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_152_ ( .D(N1211), .CP(clk), .Q(
        i_cmd_reg[152]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_151_ ( .D(N1210), .CP(clk), .Q(
        i_cmd_reg[151]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_150_ ( .D(N1209), .CP(clk), .Q(
        i_cmd_reg[150]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_149_ ( .D(N1208), .CP(clk), .Q(
        i_cmd_reg[149]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_148_ ( .D(N1207), .CP(clk), .Q(
        i_cmd_reg[148]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_146_ ( .D(N1205), .CP(clk), .Q(
        i_cmd_reg[146]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_145_ ( .D(N1204), .CP(clk), .Q(
        i_cmd_reg[145]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_144_ ( .D(N1203), .CP(clk), .Q(
        i_cmd_reg[144]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_143_ ( .D(N1202), .CP(clk), .Q(
        i_cmd_reg[143]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_142_ ( .D(N1201), .CP(clk), .Q(
        i_cmd_reg[142]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_141_ ( .D(N1200), .CP(clk), .Q(
        i_cmd_reg[141]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_140_ ( .D(N1199), .CP(clk), .Q(
        i_cmd_reg[140]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_138_ ( .D(N1197), .CP(clk), .Q(
        i_cmd_reg[138]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_137_ ( .D(N1196), .CP(clk), .Q(
        i_cmd_reg[137]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_136_ ( .D(N1195), .CP(clk), .Q(
        i_cmd_reg[136]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_135_ ( .D(N1194), .CP(clk), .Q(
        i_cmd_reg[135]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_134_ ( .D(N1193), .CP(clk), .Q(
        i_cmd_reg[134]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_133_ ( .D(N1192), .CP(clk), .Q(
        i_cmd_reg[133]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_132_ ( .D(N1191), .CP(clk), .Q(
        i_cmd_reg[132]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_131_ ( .D(N1190), .CP(clk), .Q(
        i_cmd_reg[131]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_130_ ( .D(N1189), .CP(clk), .Q(
        i_cmd_reg[130]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_129_ ( .D(N1188), .CP(clk), .Q(
        i_cmd_reg[129]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_128_ ( .D(N1187), .CP(clk), .Q(
        i_cmd_reg[128]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_127_ ( .D(N1186), .CP(clk), .Q(
        i_cmd_reg[127]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_126_ ( .D(N1185), .CP(clk), .Q(
        i_cmd_reg[126]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_125_ ( .D(N1184), .CP(clk), .Q(
        i_cmd_reg[125]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_124_ ( .D(N1183), .CP(clk), .Q(
        i_cmd_reg[124]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_123_ ( .D(N1182), .CP(clk), .Q(
        i_cmd_reg[123]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_122_ ( .D(N1181), .CP(clk), .Q(
        i_cmd_reg[122]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_121_ ( .D(N1180), .CP(clk), .Q(
        i_cmd_reg[121]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_120_ ( .D(N1179), .CP(clk), .Q(
        i_cmd_reg[120]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_119_ ( .D(N1178), .CP(clk), .Q(
        i_cmd_reg[119]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_118_ ( .D(N1177), .CP(clk), .Q(
        i_cmd_reg[118]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_117_ ( .D(N1176), .CP(clk), .Q(
        i_cmd_reg[117]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_116_ ( .D(N1175), .CP(clk), .Q(
        i_cmd_reg[116]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_115_ ( .D(N1174), .CP(clk), .Q(
        i_cmd_reg[115]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_114_ ( .D(N1173), .CP(clk), .Q(
        i_cmd_reg[114]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_113_ ( .D(N1172), .CP(clk), .Q(
        i_cmd_reg[113]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_112_ ( .D(N1171), .CP(clk), .Q(
        i_cmd_reg[112]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_111_ ( .D(N1170), .CP(clk), .Q(
        i_cmd_reg[111]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_110_ ( .D(N1169), .CP(clk), .Q(
        i_cmd_reg[110]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_109_ ( .D(N1168), .CP(clk), .Q(
        i_cmd_reg[109]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_108_ ( .D(N1167), .CP(clk), .Q(
        i_cmd_reg[108]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_107_ ( .D(N1166), .CP(clk), .Q(
        i_cmd_reg[107]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_106_ ( .D(N1165), .CP(clk), .Q(
        i_cmd_reg[106]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_105_ ( .D(N1164), .CP(clk), .Q(
        i_cmd_reg[105]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_104_ ( .D(N1163), .CP(clk), .Q(
        i_cmd_reg[104]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_103_ ( .D(N1162), .CP(clk), .Q(
        i_cmd_reg[103]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_102_ ( .D(N1161), .CP(clk), .Q(
        i_cmd_reg[102]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_101_ ( .D(N1160), .CP(clk), .Q(
        i_cmd_reg[101]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_100_ ( .D(N1159), .CP(clk), .Q(
        i_cmd_reg[100]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_99_ ( .D(N1158), .CP(clk), .Q(i_cmd_reg[99])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_98_ ( .D(N1157), .CP(clk), .Q(i_cmd_reg[98])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_97_ ( .D(N1156), .CP(clk), .Q(i_cmd_reg[97])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_96_ ( .D(N1155), .CP(clk), .Q(i_cmd_reg[96])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_95_ ( .D(N1154), .CP(clk), .Q(i_cmd_reg[95])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_94_ ( .D(N1153), .CP(clk), .Q(i_cmd_reg[94])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_93_ ( .D(N1152), .CP(clk), .Q(i_cmd_reg[93])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_92_ ( .D(N1151), .CP(clk), .Q(i_cmd_reg[92])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_91_ ( .D(N1150), .CP(clk), .Q(i_cmd_reg[91])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_90_ ( .D(N1149), .CP(clk), .Q(i_cmd_reg[90])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_89_ ( .D(N1148), .CP(clk), .Q(i_cmd_reg[89])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_88_ ( .D(N1147), .CP(clk), .Q(i_cmd_reg[88])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_87_ ( .D(N1146), .CP(clk), .Q(i_cmd_reg[87])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_86_ ( .D(N1145), .CP(clk), .Q(i_cmd_reg[86])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_85_ ( .D(N1144), .CP(clk), .Q(i_cmd_reg[85])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_84_ ( .D(N1143), .CP(clk), .Q(i_cmd_reg[84])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_83_ ( .D(N1142), .CP(clk), .Q(i_cmd_reg[83])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_82_ ( .D(N1141), .CP(clk), .Q(i_cmd_reg[82])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_81_ ( .D(N1140), .CP(clk), .Q(i_cmd_reg[81])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_80_ ( .D(N1139), .CP(clk), .Q(i_cmd_reg[80])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_79_ ( .D(N1138), .CP(clk), .Q(i_cmd_reg[79])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_78_ ( .D(N1137), .CP(clk), .Q(i_cmd_reg[78])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_77_ ( .D(N1136), .CP(clk), .Q(i_cmd_reg[77])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_76_ ( .D(N1135), .CP(clk), .Q(i_cmd_reg[76])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_75_ ( .D(N1134), .CP(clk), .Q(i_cmd_reg[75])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_74_ ( .D(N1133), .CP(clk), .Q(i_cmd_reg[74])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_73_ ( .D(N1132), .CP(clk), .Q(i_cmd_reg[73])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_72_ ( .D(N1131), .CP(clk), .Q(i_cmd_reg[72])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_71_ ( .D(N1130), .CP(clk), .Q(i_cmd_reg[71])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_70_ ( .D(N1129), .CP(clk), .Q(i_cmd_reg[70])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_69_ ( .D(N1128), .CP(clk), .Q(i_cmd_reg[69])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_68_ ( .D(N1127), .CP(clk), .Q(i_cmd_reg[68])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_67_ ( .D(N1126), .CP(clk), .Q(i_cmd_reg[67])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_66_ ( .D(N1125), .CP(clk), .Q(i_cmd_reg[66])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_65_ ( .D(N1124), .CP(clk), .Q(i_cmd_reg[65])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_64_ ( .D(N1123), .CP(clk), .Q(i_cmd_reg[64])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_63_ ( .D(N1122), .CP(clk), .Q(i_cmd_reg[63])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_62_ ( .D(N1121), .CP(clk), .Q(i_cmd_reg[62])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_61_ ( .D(N1120), .CP(clk), .Q(i_cmd_reg[61])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_60_ ( .D(N1119), .CP(clk), .Q(i_cmd_reg[60])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_59_ ( .D(N1118), .CP(clk), .Q(i_cmd_reg[59])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_58_ ( .D(N1117), .CP(clk), .Q(i_cmd_reg[58])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_57_ ( .D(N1116), .CP(clk), .Q(i_cmd_reg[57])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_56_ ( .D(N1115), .CP(clk), .Q(i_cmd_reg[56])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_55_ ( .D(N1114), .CP(clk), .Q(i_cmd_reg[55])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_54_ ( .D(N1113), .CP(clk), .Q(i_cmd_reg[54])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_53_ ( .D(N1112), .CP(clk), .Q(i_cmd_reg[53])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_52_ ( .D(N1111), .CP(clk), .Q(i_cmd_reg[52])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_51_ ( .D(N1110), .CP(clk), .Q(i_cmd_reg[51])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_50_ ( .D(N1109), .CP(clk), .Q(i_cmd_reg[50])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_49_ ( .D(N1108), .CP(clk), .Q(i_cmd_reg[49])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_48_ ( .D(N1107), .CP(clk), .Q(i_cmd_reg[48])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_47_ ( .D(N1106), .CP(clk), .Q(i_cmd_reg[47])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_46_ ( .D(N1105), .CP(clk), .Q(i_cmd_reg[46])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_45_ ( .D(N1104), .CP(clk), .Q(i_cmd_reg[45])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_44_ ( .D(N1103), .CP(clk), .Q(i_cmd_reg[44])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_43_ ( .D(N1102), .CP(clk), .Q(i_cmd_reg[43])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_42_ ( .D(N1101), .CP(clk), .Q(i_cmd_reg[42])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_41_ ( .D(N1100), .CP(clk), .Q(i_cmd_reg[41])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_40_ ( .D(N1099), .CP(clk), .Q(i_cmd_reg[40])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_39_ ( .D(N1098), .CP(clk), .Q(i_cmd_reg[39])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_38_ ( .D(N1097), .CP(clk), .Q(i_cmd_reg[38])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_37_ ( .D(N1096), .CP(clk), .Q(i_cmd_reg[37])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_36_ ( .D(N1095), .CP(clk), .Q(i_cmd_reg[36])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_35_ ( .D(N1094), .CP(clk), .Q(i_cmd_reg[35])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_34_ ( .D(N1093), .CP(clk), .Q(i_cmd_reg[34])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_33_ ( .D(N1092), .CP(clk), .Q(i_cmd_reg[33])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_32_ ( .D(N1091), .CP(clk), .Q(i_cmd_reg[32])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_31_ ( .D(N1090), .CP(clk), .Q(i_cmd_reg[31])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_30_ ( .D(N1089), .CP(clk), .Q(i_cmd_reg[30])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_29_ ( .D(N1088), .CP(clk), .Q(i_cmd_reg[29])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_28_ ( .D(N1087), .CP(clk), .Q(i_cmd_reg[28])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_27_ ( .D(N1086), .CP(clk), .Q(i_cmd_reg[27])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_26_ ( .D(N1085), .CP(clk), .Q(i_cmd_reg[26])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_25_ ( .D(N1084), .CP(clk), .Q(i_cmd_reg[25])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_24_ ( .D(N1083), .CP(clk), .Q(i_cmd_reg[24])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_23_ ( .D(N1082), .CP(clk), .Q(i_cmd_reg[23])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_22_ ( .D(N1081), .CP(clk), .Q(i_cmd_reg[22])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_21_ ( .D(N1080), .CP(clk), .Q(i_cmd_reg[21])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_20_ ( .D(N1079), .CP(clk), .Q(i_cmd_reg[20])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_19_ ( .D(N1078), .CP(clk), .Q(i_cmd_reg[19])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_18_ ( .D(N1077), .CP(clk), .Q(i_cmd_reg[18])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_17_ ( .D(N1076), .CP(clk), .Q(i_cmd_reg[17])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_16_ ( .D(N1075), .CP(clk), .Q(i_cmd_reg[16])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_15_ ( .D(N1074), .CP(clk), .Q(i_cmd_reg[15])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_14_ ( .D(N1073), .CP(clk), .Q(i_cmd_reg[14])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_13_ ( .D(N1072), .CP(clk), .Q(i_cmd_reg[13])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_12_ ( .D(N1071), .CP(clk), .Q(i_cmd_reg[12])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_11_ ( .D(N1070), .CP(clk), .Q(i_cmd_reg[11])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_10_ ( .D(N1069), .CP(clk), .Q(i_cmd_reg[10])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_9_ ( .D(N1068), .CP(clk), .Q(i_cmd_reg[9])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_8_ ( .D(N1067), .CP(clk), .Q(i_cmd_reg[8])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_7_ ( .D(N1066), .CP(clk), .Q(i_cmd_reg[7])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_6_ ( .D(N1065), .CP(clk), .Q(i_cmd_reg[6])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_5_ ( .D(N1064), .CP(clk), .Q(i_cmd_reg[5])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_4_ ( .D(N1063), .CP(clk), .Q(i_cmd_reg[4])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_3_ ( .D(N1062), .CP(clk), .Q(i_cmd_reg[3])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_2_ ( .D(N1061), .CP(clk), .Q(i_cmd_reg[2])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_1_ ( .D(N1060), .CP(clk), .Q(i_cmd_reg[1])
         );
  DFQD1BWP30P140LVT i_cmd_reg_reg_0_ ( .D(N1059), .CP(clk), .Q(i_cmd_reg[0])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_31_ ( .D(N34), .CP(clk), .Q(
        i_valid_reg[31]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_30_ ( .D(N33), .CP(clk), .Q(
        i_valid_reg[30]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_29_ ( .D(N32), .CP(clk), .Q(
        i_valid_reg[29]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_28_ ( .D(N31), .CP(clk), .Q(
        i_valid_reg[28]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_27_ ( .D(N30), .CP(clk), .Q(
        i_valid_reg[27]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_26_ ( .D(N29), .CP(clk), .Q(
        i_valid_reg[26]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_25_ ( .D(N28), .CP(clk), .Q(
        i_valid_reg[25]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_24_ ( .D(N27), .CP(clk), .Q(
        i_valid_reg[24]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_23_ ( .D(N26), .CP(clk), .Q(
        i_valid_reg[23]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_22_ ( .D(N25), .CP(clk), .Q(
        i_valid_reg[22]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_21_ ( .D(N24), .CP(clk), .Q(
        i_valid_reg[21]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_20_ ( .D(N23), .CP(clk), .Q(
        i_valid_reg[20]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_19_ ( .D(N22), .CP(clk), .Q(
        i_valid_reg[19]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_18_ ( .D(N21), .CP(clk), .Q(
        i_valid_reg[18]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_17_ ( .D(N20), .CP(clk), .Q(
        i_valid_reg[17]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_16_ ( .D(N19), .CP(clk), .Q(
        i_valid_reg[16]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_15_ ( .D(N18), .CP(clk), .Q(
        i_valid_reg[15]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_14_ ( .D(N17), .CP(clk), .Q(
        i_valid_reg[14]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_13_ ( .D(N16), .CP(clk), .Q(
        i_valid_reg[13]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_12_ ( .D(N15), .CP(clk), .Q(
        i_valid_reg[12]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_11_ ( .D(N14), .CP(clk), .Q(
        i_valid_reg[11]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_10_ ( .D(N13), .CP(clk), .Q(
        i_valid_reg[10]) );
  DFQD1BWP30P140LVT i_valid_reg_reg_9_ ( .D(N12), .CP(clk), .Q(i_valid_reg[9])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_8_ ( .D(N11), .CP(clk), .Q(i_valid_reg[8])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_7_ ( .D(N10), .CP(clk), .Q(i_valid_reg[7])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_6_ ( .D(N9), .CP(clk), .Q(i_valid_reg[6])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_5_ ( .D(N8), .CP(clk), .Q(i_valid_reg[5])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_4_ ( .D(N7), .CP(clk), .Q(i_valid_reg[4])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_3_ ( .D(N6), .CP(clk), .Q(i_valid_reg[3])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_2_ ( .D(N5), .CP(clk), .Q(i_valid_reg[2])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_1_ ( .D(N4), .CP(clk), .Q(i_valid_reg[1])
         );
  DFQD1BWP30P140LVT i_valid_reg_reg_0_ ( .D(N3), .CP(clk), .Q(i_valid_reg[0])
         );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1023_ ( .D(N1058), .CP(clk), .Q(
        i_data_bus_reg[1023]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1022_ ( .D(N1057), .CP(clk), .Q(
        i_data_bus_reg[1022]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1021_ ( .D(N1056), .CP(clk), .Q(
        i_data_bus_reg[1021]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1020_ ( .D(N1055), .CP(clk), .Q(
        i_data_bus_reg[1020]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1019_ ( .D(N1054), .CP(clk), .Q(
        i_data_bus_reg[1019]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1018_ ( .D(N1053), .CP(clk), .Q(
        i_data_bus_reg[1018]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1017_ ( .D(N1052), .CP(clk), .Q(
        i_data_bus_reg[1017]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1016_ ( .D(N1051), .CP(clk), .Q(
        i_data_bus_reg[1016]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1015_ ( .D(N1050), .CP(clk), .Q(
        i_data_bus_reg[1015]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1014_ ( .D(N1049), .CP(clk), .Q(
        i_data_bus_reg[1014]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1013_ ( .D(N1048), .CP(clk), .Q(
        i_data_bus_reg[1013]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1012_ ( .D(N1047), .CP(clk), .Q(
        i_data_bus_reg[1012]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1011_ ( .D(N1046), .CP(clk), .Q(
        i_data_bus_reg[1011]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1010_ ( .D(N1045), .CP(clk), .Q(
        i_data_bus_reg[1010]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1009_ ( .D(N1044), .CP(clk), .Q(
        i_data_bus_reg[1009]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1008_ ( .D(N1043), .CP(clk), .Q(
        i_data_bus_reg[1008]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1007_ ( .D(N1042), .CP(clk), .Q(
        i_data_bus_reg[1007]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1006_ ( .D(N1041), .CP(clk), .Q(
        i_data_bus_reg[1006]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1005_ ( .D(N1040), .CP(clk), .Q(
        i_data_bus_reg[1005]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1004_ ( .D(N1039), .CP(clk), .Q(
        i_data_bus_reg[1004]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1003_ ( .D(N1038), .CP(clk), .Q(
        i_data_bus_reg[1003]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1002_ ( .D(N1037), .CP(clk), .Q(
        i_data_bus_reg[1002]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1001_ ( .D(N1036), .CP(clk), .Q(
        i_data_bus_reg[1001]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1000_ ( .D(N1035), .CP(clk), .Q(
        i_data_bus_reg[1000]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_999_ ( .D(N1034), .CP(clk), .Q(
        i_data_bus_reg[999]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_998_ ( .D(N1033), .CP(clk), .Q(
        i_data_bus_reg[998]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_997_ ( .D(N1032), .CP(clk), .Q(
        i_data_bus_reg[997]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_996_ ( .D(N1031), .CP(clk), .Q(
        i_data_bus_reg[996]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_995_ ( .D(N1030), .CP(clk), .Q(
        i_data_bus_reg[995]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_994_ ( .D(N1029), .CP(clk), .Q(
        i_data_bus_reg[994]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_993_ ( .D(N1028), .CP(clk), .Q(
        i_data_bus_reg[993]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_992_ ( .D(N1027), .CP(clk), .Q(
        i_data_bus_reg[992]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_991_ ( .D(N1026), .CP(clk), .Q(
        i_data_bus_reg[991]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_990_ ( .D(N1025), .CP(clk), .Q(
        i_data_bus_reg[990]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_989_ ( .D(N1024), .CP(clk), .Q(
        i_data_bus_reg[989]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_988_ ( .D(N1023), .CP(clk), .Q(
        i_data_bus_reg[988]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_987_ ( .D(N1022), .CP(clk), .Q(
        i_data_bus_reg[987]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_986_ ( .D(N1021), .CP(clk), .Q(
        i_data_bus_reg[986]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_985_ ( .D(N1020), .CP(clk), .Q(
        i_data_bus_reg[985]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_984_ ( .D(N1019), .CP(clk), .Q(
        i_data_bus_reg[984]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_983_ ( .D(N1018), .CP(clk), .Q(
        i_data_bus_reg[983]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_982_ ( .D(N1017), .CP(clk), .Q(
        i_data_bus_reg[982]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_981_ ( .D(N1016), .CP(clk), .Q(
        i_data_bus_reg[981]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_980_ ( .D(N1015), .CP(clk), .Q(
        i_data_bus_reg[980]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_979_ ( .D(N1014), .CP(clk), .Q(
        i_data_bus_reg[979]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_978_ ( .D(N1013), .CP(clk), .Q(
        i_data_bus_reg[978]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_977_ ( .D(N1012), .CP(clk), .Q(
        i_data_bus_reg[977]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_976_ ( .D(N1011), .CP(clk), .Q(
        i_data_bus_reg[976]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_975_ ( .D(N1010), .CP(clk), .Q(
        i_data_bus_reg[975]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_974_ ( .D(N1009), .CP(clk), .Q(
        i_data_bus_reg[974]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_973_ ( .D(N1008), .CP(clk), .Q(
        i_data_bus_reg[973]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_972_ ( .D(N1007), .CP(clk), .Q(
        i_data_bus_reg[972]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_971_ ( .D(N1006), .CP(clk), .Q(
        i_data_bus_reg[971]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_970_ ( .D(N1005), .CP(clk), .Q(
        i_data_bus_reg[970]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_969_ ( .D(N1004), .CP(clk), .Q(
        i_data_bus_reg[969]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_968_ ( .D(N1003), .CP(clk), .Q(
        i_data_bus_reg[968]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_967_ ( .D(N1002), .CP(clk), .Q(
        i_data_bus_reg[967]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_966_ ( .D(N1001), .CP(clk), .Q(
        i_data_bus_reg[966]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_965_ ( .D(N1000), .CP(clk), .Q(
        i_data_bus_reg[965]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_964_ ( .D(N999), .CP(clk), .Q(
        i_data_bus_reg[964]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_963_ ( .D(N998), .CP(clk), .Q(
        i_data_bus_reg[963]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_962_ ( .D(N997), .CP(clk), .Q(
        i_data_bus_reg[962]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_961_ ( .D(N996), .CP(clk), .Q(
        i_data_bus_reg[961]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_960_ ( .D(N995), .CP(clk), .Q(
        i_data_bus_reg[960]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_959_ ( .D(N994), .CP(clk), .Q(
        i_data_bus_reg[959]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_958_ ( .D(N993), .CP(clk), .Q(
        i_data_bus_reg[958]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_957_ ( .D(N992), .CP(clk), .Q(
        i_data_bus_reg[957]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_956_ ( .D(N991), .CP(clk), .Q(
        i_data_bus_reg[956]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_955_ ( .D(N990), .CP(clk), .Q(
        i_data_bus_reg[955]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_954_ ( .D(N989), .CP(clk), .Q(
        i_data_bus_reg[954]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_953_ ( .D(N988), .CP(clk), .Q(
        i_data_bus_reg[953]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_952_ ( .D(N987), .CP(clk), .Q(
        i_data_bus_reg[952]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_951_ ( .D(N986), .CP(clk), .Q(
        i_data_bus_reg[951]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_950_ ( .D(N985), .CP(clk), .Q(
        i_data_bus_reg[950]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_949_ ( .D(N984), .CP(clk), .Q(
        i_data_bus_reg[949]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_948_ ( .D(N983), .CP(clk), .Q(
        i_data_bus_reg[948]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_947_ ( .D(N982), .CP(clk), .Q(
        i_data_bus_reg[947]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_946_ ( .D(N981), .CP(clk), .Q(
        i_data_bus_reg[946]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_945_ ( .D(N980), .CP(clk), .Q(
        i_data_bus_reg[945]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_944_ ( .D(N979), .CP(clk), .Q(
        i_data_bus_reg[944]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_943_ ( .D(N978), .CP(clk), .Q(
        i_data_bus_reg[943]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_942_ ( .D(N977), .CP(clk), .Q(
        i_data_bus_reg[942]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_941_ ( .D(N976), .CP(clk), .Q(
        i_data_bus_reg[941]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_940_ ( .D(N975), .CP(clk), .Q(
        i_data_bus_reg[940]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_939_ ( .D(N974), .CP(clk), .Q(
        i_data_bus_reg[939]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_938_ ( .D(N973), .CP(clk), .Q(
        i_data_bus_reg[938]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_937_ ( .D(N972), .CP(clk), .Q(
        i_data_bus_reg[937]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_936_ ( .D(N971), .CP(clk), .Q(
        i_data_bus_reg[936]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_935_ ( .D(N970), .CP(clk), .Q(
        i_data_bus_reg[935]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_934_ ( .D(N969), .CP(clk), .Q(
        i_data_bus_reg[934]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_933_ ( .D(N968), .CP(clk), .Q(
        i_data_bus_reg[933]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_932_ ( .D(N967), .CP(clk), .Q(
        i_data_bus_reg[932]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_931_ ( .D(N966), .CP(clk), .Q(
        i_data_bus_reg[931]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_930_ ( .D(N965), .CP(clk), .Q(
        i_data_bus_reg[930]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_929_ ( .D(N964), .CP(clk), .Q(
        i_data_bus_reg[929]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_928_ ( .D(N963), .CP(clk), .Q(
        i_data_bus_reg[928]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_927_ ( .D(N962), .CP(clk), .Q(
        i_data_bus_reg[927]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_926_ ( .D(N961), .CP(clk), .Q(
        i_data_bus_reg[926]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_925_ ( .D(N960), .CP(clk), .Q(
        i_data_bus_reg[925]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_924_ ( .D(N959), .CP(clk), .Q(
        i_data_bus_reg[924]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_923_ ( .D(N958), .CP(clk), .Q(
        i_data_bus_reg[923]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_922_ ( .D(N957), .CP(clk), .Q(
        i_data_bus_reg[922]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_921_ ( .D(N956), .CP(clk), .Q(
        i_data_bus_reg[921]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_920_ ( .D(N955), .CP(clk), .Q(
        i_data_bus_reg[920]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_919_ ( .D(N954), .CP(clk), .Q(
        i_data_bus_reg[919]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_918_ ( .D(N953), .CP(clk), .Q(
        i_data_bus_reg[918]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_917_ ( .D(N952), .CP(clk), .Q(
        i_data_bus_reg[917]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_916_ ( .D(N951), .CP(clk), .Q(
        i_data_bus_reg[916]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_915_ ( .D(N950), .CP(clk), .Q(
        i_data_bus_reg[915]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_914_ ( .D(N949), .CP(clk), .Q(
        i_data_bus_reg[914]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_913_ ( .D(N948), .CP(clk), .Q(
        i_data_bus_reg[913]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_912_ ( .D(N947), .CP(clk), .Q(
        i_data_bus_reg[912]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_911_ ( .D(N946), .CP(clk), .Q(
        i_data_bus_reg[911]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_910_ ( .D(N945), .CP(clk), .Q(
        i_data_bus_reg[910]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_909_ ( .D(N944), .CP(clk), .Q(
        i_data_bus_reg[909]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_908_ ( .D(N943), .CP(clk), .Q(
        i_data_bus_reg[908]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_907_ ( .D(N942), .CP(clk), .Q(
        i_data_bus_reg[907]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_906_ ( .D(N941), .CP(clk), .Q(
        i_data_bus_reg[906]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_905_ ( .D(N940), .CP(clk), .Q(
        i_data_bus_reg[905]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_904_ ( .D(N939), .CP(clk), .Q(
        i_data_bus_reg[904]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_903_ ( .D(N938), .CP(clk), .Q(
        i_data_bus_reg[903]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_902_ ( .D(N937), .CP(clk), .Q(
        i_data_bus_reg[902]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_901_ ( .D(N936), .CP(clk), .Q(
        i_data_bus_reg[901]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_900_ ( .D(N935), .CP(clk), .Q(
        i_data_bus_reg[900]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_899_ ( .D(N934), .CP(clk), .Q(
        i_data_bus_reg[899]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_898_ ( .D(N933), .CP(clk), .Q(
        i_data_bus_reg[898]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_897_ ( .D(N932), .CP(clk), .Q(
        i_data_bus_reg[897]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_896_ ( .D(N931), .CP(clk), .Q(
        i_data_bus_reg[896]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_895_ ( .D(N930), .CP(clk), .Q(
        i_data_bus_reg[895]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_894_ ( .D(N929), .CP(clk), .Q(
        i_data_bus_reg[894]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_893_ ( .D(N928), .CP(clk), .Q(
        i_data_bus_reg[893]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_892_ ( .D(N927), .CP(clk), .Q(
        i_data_bus_reg[892]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_891_ ( .D(N926), .CP(clk), .Q(
        i_data_bus_reg[891]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_890_ ( .D(N925), .CP(clk), .Q(
        i_data_bus_reg[890]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_889_ ( .D(N924), .CP(clk), .Q(
        i_data_bus_reg[889]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_888_ ( .D(N923), .CP(clk), .Q(
        i_data_bus_reg[888]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_887_ ( .D(N922), .CP(clk), .Q(
        i_data_bus_reg[887]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_886_ ( .D(N921), .CP(clk), .Q(
        i_data_bus_reg[886]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_885_ ( .D(N920), .CP(clk), .Q(
        i_data_bus_reg[885]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_884_ ( .D(N919), .CP(clk), .Q(
        i_data_bus_reg[884]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_883_ ( .D(N918), .CP(clk), .Q(
        i_data_bus_reg[883]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_882_ ( .D(N917), .CP(clk), .Q(
        i_data_bus_reg[882]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_881_ ( .D(N916), .CP(clk), .Q(
        i_data_bus_reg[881]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_880_ ( .D(N915), .CP(clk), .Q(
        i_data_bus_reg[880]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_879_ ( .D(N914), .CP(clk), .Q(
        i_data_bus_reg[879]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_878_ ( .D(N913), .CP(clk), .Q(
        i_data_bus_reg[878]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_877_ ( .D(N912), .CP(clk), .Q(
        i_data_bus_reg[877]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_876_ ( .D(N911), .CP(clk), .Q(
        i_data_bus_reg[876]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_875_ ( .D(N910), .CP(clk), .Q(
        i_data_bus_reg[875]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_874_ ( .D(N909), .CP(clk), .Q(
        i_data_bus_reg[874]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_873_ ( .D(N908), .CP(clk), .Q(
        i_data_bus_reg[873]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_872_ ( .D(N907), .CP(clk), .Q(
        i_data_bus_reg[872]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_871_ ( .D(N906), .CP(clk), .Q(
        i_data_bus_reg[871]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_870_ ( .D(N905), .CP(clk), .Q(
        i_data_bus_reg[870]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_869_ ( .D(N904), .CP(clk), .Q(
        i_data_bus_reg[869]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_868_ ( .D(N903), .CP(clk), .Q(
        i_data_bus_reg[868]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_867_ ( .D(N902), .CP(clk), .Q(
        i_data_bus_reg[867]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_866_ ( .D(N901), .CP(clk), .Q(
        i_data_bus_reg[866]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_865_ ( .D(N900), .CP(clk), .Q(
        i_data_bus_reg[865]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_864_ ( .D(N899), .CP(clk), .Q(
        i_data_bus_reg[864]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_863_ ( .D(N898), .CP(clk), .Q(
        i_data_bus_reg[863]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_862_ ( .D(N897), .CP(clk), .Q(
        i_data_bus_reg[862]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_861_ ( .D(N896), .CP(clk), .Q(
        i_data_bus_reg[861]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_860_ ( .D(N895), .CP(clk), .Q(
        i_data_bus_reg[860]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_859_ ( .D(N894), .CP(clk), .Q(
        i_data_bus_reg[859]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_858_ ( .D(N893), .CP(clk), .Q(
        i_data_bus_reg[858]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_857_ ( .D(N892), .CP(clk), .Q(
        i_data_bus_reg[857]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_856_ ( .D(N891), .CP(clk), .Q(
        i_data_bus_reg[856]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_855_ ( .D(N890), .CP(clk), .Q(
        i_data_bus_reg[855]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_854_ ( .D(N889), .CP(clk), .Q(
        i_data_bus_reg[854]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_853_ ( .D(N888), .CP(clk), .Q(
        i_data_bus_reg[853]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_852_ ( .D(N887), .CP(clk), .Q(
        i_data_bus_reg[852]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_851_ ( .D(N886), .CP(clk), .Q(
        i_data_bus_reg[851]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_850_ ( .D(N885), .CP(clk), .Q(
        i_data_bus_reg[850]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_849_ ( .D(N884), .CP(clk), .Q(
        i_data_bus_reg[849]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_848_ ( .D(N883), .CP(clk), .Q(
        i_data_bus_reg[848]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_847_ ( .D(N882), .CP(clk), .Q(
        i_data_bus_reg[847]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_846_ ( .D(N881), .CP(clk), .Q(
        i_data_bus_reg[846]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_845_ ( .D(N880), .CP(clk), .Q(
        i_data_bus_reg[845]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_844_ ( .D(N879), .CP(clk), .Q(
        i_data_bus_reg[844]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_843_ ( .D(N878), .CP(clk), .Q(
        i_data_bus_reg[843]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_842_ ( .D(N877), .CP(clk), .Q(
        i_data_bus_reg[842]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_841_ ( .D(N876), .CP(clk), .Q(
        i_data_bus_reg[841]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_840_ ( .D(N875), .CP(clk), .Q(
        i_data_bus_reg[840]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_839_ ( .D(N874), .CP(clk), .Q(
        i_data_bus_reg[839]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_838_ ( .D(N873), .CP(clk), .Q(
        i_data_bus_reg[838]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_837_ ( .D(N872), .CP(clk), .Q(
        i_data_bus_reg[837]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_836_ ( .D(N871), .CP(clk), .Q(
        i_data_bus_reg[836]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_835_ ( .D(N870), .CP(clk), .Q(
        i_data_bus_reg[835]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_834_ ( .D(N869), .CP(clk), .Q(
        i_data_bus_reg[834]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_833_ ( .D(N868), .CP(clk), .Q(
        i_data_bus_reg[833]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_832_ ( .D(N867), .CP(clk), .Q(
        i_data_bus_reg[832]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_831_ ( .D(N866), .CP(clk), .Q(
        i_data_bus_reg[831]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_830_ ( .D(N865), .CP(clk), .Q(
        i_data_bus_reg[830]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_829_ ( .D(N864), .CP(clk), .Q(
        i_data_bus_reg[829]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_828_ ( .D(N863), .CP(clk), .Q(
        i_data_bus_reg[828]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_827_ ( .D(N862), .CP(clk), .Q(
        i_data_bus_reg[827]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_826_ ( .D(N861), .CP(clk), .Q(
        i_data_bus_reg[826]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_825_ ( .D(N860), .CP(clk), .Q(
        i_data_bus_reg[825]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_824_ ( .D(N859), .CP(clk), .Q(
        i_data_bus_reg[824]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_823_ ( .D(N858), .CP(clk), .Q(
        i_data_bus_reg[823]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_822_ ( .D(N857), .CP(clk), .Q(
        i_data_bus_reg[822]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_821_ ( .D(N856), .CP(clk), .Q(
        i_data_bus_reg[821]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_820_ ( .D(N855), .CP(clk), .Q(
        i_data_bus_reg[820]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_819_ ( .D(N854), .CP(clk), .Q(
        i_data_bus_reg[819]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_818_ ( .D(N853), .CP(clk), .Q(
        i_data_bus_reg[818]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_817_ ( .D(N852), .CP(clk), .Q(
        i_data_bus_reg[817]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_816_ ( .D(N851), .CP(clk), .Q(
        i_data_bus_reg[816]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_815_ ( .D(N850), .CP(clk), .Q(
        i_data_bus_reg[815]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_814_ ( .D(N849), .CP(clk), .Q(
        i_data_bus_reg[814]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_813_ ( .D(N848), .CP(clk), .Q(
        i_data_bus_reg[813]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_812_ ( .D(N847), .CP(clk), .Q(
        i_data_bus_reg[812]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_811_ ( .D(N846), .CP(clk), .Q(
        i_data_bus_reg[811]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_810_ ( .D(N845), .CP(clk), .Q(
        i_data_bus_reg[810]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_809_ ( .D(N844), .CP(clk), .Q(
        i_data_bus_reg[809]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_808_ ( .D(N843), .CP(clk), .Q(
        i_data_bus_reg[808]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_807_ ( .D(N842), .CP(clk), .Q(
        i_data_bus_reg[807]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_806_ ( .D(N841), .CP(clk), .Q(
        i_data_bus_reg[806]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_805_ ( .D(N840), .CP(clk), .Q(
        i_data_bus_reg[805]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_804_ ( .D(N839), .CP(clk), .Q(
        i_data_bus_reg[804]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_803_ ( .D(N838), .CP(clk), .Q(
        i_data_bus_reg[803]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_802_ ( .D(N837), .CP(clk), .Q(
        i_data_bus_reg[802]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_801_ ( .D(N836), .CP(clk), .Q(
        i_data_bus_reg[801]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_800_ ( .D(N835), .CP(clk), .Q(
        i_data_bus_reg[800]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_799_ ( .D(N834), .CP(clk), .Q(
        i_data_bus_reg[799]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_798_ ( .D(N833), .CP(clk), .Q(
        i_data_bus_reg[798]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_797_ ( .D(N832), .CP(clk), .Q(
        i_data_bus_reg[797]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_796_ ( .D(N831), .CP(clk), .Q(
        i_data_bus_reg[796]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_795_ ( .D(N830), .CP(clk), .Q(
        i_data_bus_reg[795]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_794_ ( .D(N829), .CP(clk), .Q(
        i_data_bus_reg[794]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_793_ ( .D(N828), .CP(clk), .Q(
        i_data_bus_reg[793]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_792_ ( .D(N827), .CP(clk), .Q(
        i_data_bus_reg[792]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_791_ ( .D(N826), .CP(clk), .Q(
        i_data_bus_reg[791]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_790_ ( .D(N825), .CP(clk), .Q(
        i_data_bus_reg[790]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_789_ ( .D(N824), .CP(clk), .Q(
        i_data_bus_reg[789]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_788_ ( .D(N823), .CP(clk), .Q(
        i_data_bus_reg[788]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_787_ ( .D(N822), .CP(clk), .Q(
        i_data_bus_reg[787]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_786_ ( .D(N821), .CP(clk), .Q(
        i_data_bus_reg[786]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_785_ ( .D(N820), .CP(clk), .Q(
        i_data_bus_reg[785]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_784_ ( .D(N819), .CP(clk), .Q(
        i_data_bus_reg[784]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_783_ ( .D(N818), .CP(clk), .Q(
        i_data_bus_reg[783]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_782_ ( .D(N817), .CP(clk), .Q(
        i_data_bus_reg[782]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_781_ ( .D(N816), .CP(clk), .Q(
        i_data_bus_reg[781]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_780_ ( .D(N815), .CP(clk), .Q(
        i_data_bus_reg[780]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_779_ ( .D(N814), .CP(clk), .Q(
        i_data_bus_reg[779]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_778_ ( .D(N813), .CP(clk), .Q(
        i_data_bus_reg[778]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_777_ ( .D(N812), .CP(clk), .Q(
        i_data_bus_reg[777]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_776_ ( .D(N811), .CP(clk), .Q(
        i_data_bus_reg[776]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_775_ ( .D(N810), .CP(clk), .Q(
        i_data_bus_reg[775]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_774_ ( .D(N809), .CP(clk), .Q(
        i_data_bus_reg[774]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_773_ ( .D(N808), .CP(clk), .Q(
        i_data_bus_reg[773]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_772_ ( .D(N807), .CP(clk), .Q(
        i_data_bus_reg[772]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_771_ ( .D(N806), .CP(clk), .Q(
        i_data_bus_reg[771]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_770_ ( .D(N805), .CP(clk), .Q(
        i_data_bus_reg[770]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_769_ ( .D(N804), .CP(clk), .Q(
        i_data_bus_reg[769]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_768_ ( .D(N803), .CP(clk), .Q(
        i_data_bus_reg[768]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_767_ ( .D(N802), .CP(clk), .Q(
        i_data_bus_reg[767]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_766_ ( .D(N801), .CP(clk), .Q(
        i_data_bus_reg[766]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_765_ ( .D(N800), .CP(clk), .Q(
        i_data_bus_reg[765]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_764_ ( .D(N799), .CP(clk), .Q(
        i_data_bus_reg[764]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_763_ ( .D(N798), .CP(clk), .Q(
        i_data_bus_reg[763]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_762_ ( .D(N797), .CP(clk), .Q(
        i_data_bus_reg[762]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_761_ ( .D(N796), .CP(clk), .Q(
        i_data_bus_reg[761]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_760_ ( .D(N795), .CP(clk), .Q(
        i_data_bus_reg[760]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_759_ ( .D(N794), .CP(clk), .Q(
        i_data_bus_reg[759]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_758_ ( .D(N793), .CP(clk), .Q(
        i_data_bus_reg[758]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_757_ ( .D(N792), .CP(clk), .Q(
        i_data_bus_reg[757]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_756_ ( .D(N791), .CP(clk), .Q(
        i_data_bus_reg[756]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_755_ ( .D(N790), .CP(clk), .Q(
        i_data_bus_reg[755]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_754_ ( .D(N789), .CP(clk), .Q(
        i_data_bus_reg[754]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_753_ ( .D(N788), .CP(clk), .Q(
        i_data_bus_reg[753]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_752_ ( .D(N787), .CP(clk), .Q(
        i_data_bus_reg[752]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_751_ ( .D(N786), .CP(clk), .Q(
        i_data_bus_reg[751]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_750_ ( .D(N785), .CP(clk), .Q(
        i_data_bus_reg[750]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_749_ ( .D(N784), .CP(clk), .Q(
        i_data_bus_reg[749]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_748_ ( .D(N783), .CP(clk), .Q(
        i_data_bus_reg[748]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_747_ ( .D(N782), .CP(clk), .Q(
        i_data_bus_reg[747]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_746_ ( .D(N781), .CP(clk), .Q(
        i_data_bus_reg[746]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_745_ ( .D(N780), .CP(clk), .Q(
        i_data_bus_reg[745]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_744_ ( .D(N779), .CP(clk), .Q(
        i_data_bus_reg[744]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_743_ ( .D(N778), .CP(clk), .Q(
        i_data_bus_reg[743]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_742_ ( .D(N777), .CP(clk), .Q(
        i_data_bus_reg[742]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_741_ ( .D(N776), .CP(clk), .Q(
        i_data_bus_reg[741]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_740_ ( .D(N775), .CP(clk), .Q(
        i_data_bus_reg[740]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_739_ ( .D(N774), .CP(clk), .Q(
        i_data_bus_reg[739]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_738_ ( .D(N773), .CP(clk), .Q(
        i_data_bus_reg[738]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_737_ ( .D(N772), .CP(clk), .Q(
        i_data_bus_reg[737]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_736_ ( .D(N771), .CP(clk), .Q(
        i_data_bus_reg[736]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_735_ ( .D(N770), .CP(clk), .Q(
        i_data_bus_reg[735]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_734_ ( .D(N769), .CP(clk), .Q(
        i_data_bus_reg[734]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_733_ ( .D(N768), .CP(clk), .Q(
        i_data_bus_reg[733]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_732_ ( .D(N767), .CP(clk), .Q(
        i_data_bus_reg[732]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_731_ ( .D(N766), .CP(clk), .Q(
        i_data_bus_reg[731]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_730_ ( .D(N765), .CP(clk), .Q(
        i_data_bus_reg[730]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_729_ ( .D(N764), .CP(clk), .Q(
        i_data_bus_reg[729]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_728_ ( .D(N763), .CP(clk), .Q(
        i_data_bus_reg[728]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_727_ ( .D(N762), .CP(clk), .Q(
        i_data_bus_reg[727]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_726_ ( .D(N761), .CP(clk), .Q(
        i_data_bus_reg[726]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_725_ ( .D(N760), .CP(clk), .Q(
        i_data_bus_reg[725]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_724_ ( .D(N759), .CP(clk), .Q(
        i_data_bus_reg[724]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_723_ ( .D(N758), .CP(clk), .Q(
        i_data_bus_reg[723]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_722_ ( .D(N757), .CP(clk), .Q(
        i_data_bus_reg[722]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_721_ ( .D(N756), .CP(clk), .Q(
        i_data_bus_reg[721]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_720_ ( .D(N755), .CP(clk), .Q(
        i_data_bus_reg[720]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_719_ ( .D(N754), .CP(clk), .Q(
        i_data_bus_reg[719]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_718_ ( .D(N753), .CP(clk), .Q(
        i_data_bus_reg[718]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_717_ ( .D(N752), .CP(clk), .Q(
        i_data_bus_reg[717]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_716_ ( .D(N751), .CP(clk), .Q(
        i_data_bus_reg[716]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_715_ ( .D(N750), .CP(clk), .Q(
        i_data_bus_reg[715]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_714_ ( .D(N749), .CP(clk), .Q(
        i_data_bus_reg[714]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_713_ ( .D(N748), .CP(clk), .Q(
        i_data_bus_reg[713]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_712_ ( .D(N747), .CP(clk), .Q(
        i_data_bus_reg[712]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_711_ ( .D(N746), .CP(clk), .Q(
        i_data_bus_reg[711]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_710_ ( .D(N745), .CP(clk), .Q(
        i_data_bus_reg[710]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_709_ ( .D(N744), .CP(clk), .Q(
        i_data_bus_reg[709]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_708_ ( .D(N743), .CP(clk), .Q(
        i_data_bus_reg[708]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_707_ ( .D(N742), .CP(clk), .Q(
        i_data_bus_reg[707]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_706_ ( .D(N741), .CP(clk), .Q(
        i_data_bus_reg[706]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_705_ ( .D(N740), .CP(clk), .Q(
        i_data_bus_reg[705]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_704_ ( .D(N739), .CP(clk), .Q(
        i_data_bus_reg[704]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_703_ ( .D(N738), .CP(clk), .Q(
        i_data_bus_reg[703]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_702_ ( .D(N737), .CP(clk), .Q(
        i_data_bus_reg[702]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_701_ ( .D(N736), .CP(clk), .Q(
        i_data_bus_reg[701]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_700_ ( .D(N735), .CP(clk), .Q(
        i_data_bus_reg[700]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_699_ ( .D(N734), .CP(clk), .Q(
        i_data_bus_reg[699]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_698_ ( .D(N733), .CP(clk), .Q(
        i_data_bus_reg[698]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_697_ ( .D(N732), .CP(clk), .Q(
        i_data_bus_reg[697]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_696_ ( .D(N731), .CP(clk), .Q(
        i_data_bus_reg[696]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_695_ ( .D(N730), .CP(clk), .Q(
        i_data_bus_reg[695]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_694_ ( .D(N729), .CP(clk), .Q(
        i_data_bus_reg[694]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_693_ ( .D(N728), .CP(clk), .Q(
        i_data_bus_reg[693]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_692_ ( .D(N727), .CP(clk), .Q(
        i_data_bus_reg[692]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_691_ ( .D(N726), .CP(clk), .Q(
        i_data_bus_reg[691]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_690_ ( .D(N725), .CP(clk), .Q(
        i_data_bus_reg[690]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_689_ ( .D(N724), .CP(clk), .Q(
        i_data_bus_reg[689]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_688_ ( .D(N723), .CP(clk), .Q(
        i_data_bus_reg[688]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_687_ ( .D(N722), .CP(clk), .Q(
        i_data_bus_reg[687]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_686_ ( .D(N721), .CP(clk), .Q(
        i_data_bus_reg[686]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_685_ ( .D(N720), .CP(clk), .Q(
        i_data_bus_reg[685]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_684_ ( .D(N719), .CP(clk), .Q(
        i_data_bus_reg[684]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_683_ ( .D(N718), .CP(clk), .Q(
        i_data_bus_reg[683]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_682_ ( .D(N717), .CP(clk), .Q(
        i_data_bus_reg[682]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_681_ ( .D(N716), .CP(clk), .Q(
        i_data_bus_reg[681]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_680_ ( .D(N715), .CP(clk), .Q(
        i_data_bus_reg[680]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_679_ ( .D(N714), .CP(clk), .Q(
        i_data_bus_reg[679]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_678_ ( .D(N713), .CP(clk), .Q(
        i_data_bus_reg[678]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_677_ ( .D(N712), .CP(clk), .Q(
        i_data_bus_reg[677]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_676_ ( .D(N711), .CP(clk), .Q(
        i_data_bus_reg[676]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_675_ ( .D(N710), .CP(clk), .Q(
        i_data_bus_reg[675]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_674_ ( .D(N709), .CP(clk), .Q(
        i_data_bus_reg[674]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_673_ ( .D(N708), .CP(clk), .Q(
        i_data_bus_reg[673]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_672_ ( .D(N707), .CP(clk), .Q(
        i_data_bus_reg[672]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_671_ ( .D(N706), .CP(clk), .Q(
        i_data_bus_reg[671]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_670_ ( .D(N705), .CP(clk), .Q(
        i_data_bus_reg[670]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_669_ ( .D(N704), .CP(clk), .Q(
        i_data_bus_reg[669]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_668_ ( .D(N703), .CP(clk), .Q(
        i_data_bus_reg[668]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_667_ ( .D(N702), .CP(clk), .Q(
        i_data_bus_reg[667]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_666_ ( .D(N701), .CP(clk), .Q(
        i_data_bus_reg[666]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_665_ ( .D(N700), .CP(clk), .Q(
        i_data_bus_reg[665]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_664_ ( .D(N699), .CP(clk), .Q(
        i_data_bus_reg[664]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_663_ ( .D(N698), .CP(clk), .Q(
        i_data_bus_reg[663]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_662_ ( .D(N697), .CP(clk), .Q(
        i_data_bus_reg[662]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_661_ ( .D(N696), .CP(clk), .Q(
        i_data_bus_reg[661]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_660_ ( .D(N695), .CP(clk), .Q(
        i_data_bus_reg[660]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_659_ ( .D(N694), .CP(clk), .Q(
        i_data_bus_reg[659]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_658_ ( .D(N693), .CP(clk), .Q(
        i_data_bus_reg[658]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_657_ ( .D(N692), .CP(clk), .Q(
        i_data_bus_reg[657]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_656_ ( .D(N691), .CP(clk), .Q(
        i_data_bus_reg[656]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_655_ ( .D(N690), .CP(clk), .Q(
        i_data_bus_reg[655]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_654_ ( .D(N689), .CP(clk), .Q(
        i_data_bus_reg[654]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_653_ ( .D(N688), .CP(clk), .Q(
        i_data_bus_reg[653]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_652_ ( .D(N687), .CP(clk), .Q(
        i_data_bus_reg[652]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_651_ ( .D(N686), .CP(clk), .Q(
        i_data_bus_reg[651]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_650_ ( .D(N685), .CP(clk), .Q(
        i_data_bus_reg[650]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_649_ ( .D(N684), .CP(clk), .Q(
        i_data_bus_reg[649]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_648_ ( .D(N683), .CP(clk), .Q(
        i_data_bus_reg[648]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_647_ ( .D(N682), .CP(clk), .Q(
        i_data_bus_reg[647]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_646_ ( .D(N681), .CP(clk), .Q(
        i_data_bus_reg[646]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_645_ ( .D(N680), .CP(clk), .Q(
        i_data_bus_reg[645]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_644_ ( .D(N679), .CP(clk), .Q(
        i_data_bus_reg[644]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_643_ ( .D(N678), .CP(clk), .Q(
        i_data_bus_reg[643]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_642_ ( .D(N677), .CP(clk), .Q(
        i_data_bus_reg[642]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_641_ ( .D(N676), .CP(clk), .Q(
        i_data_bus_reg[641]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_640_ ( .D(N675), .CP(clk), .Q(
        i_data_bus_reg[640]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_639_ ( .D(N674), .CP(clk), .Q(
        i_data_bus_reg[639]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_638_ ( .D(N673), .CP(clk), .Q(
        i_data_bus_reg[638]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_637_ ( .D(N672), .CP(clk), .Q(
        i_data_bus_reg[637]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_636_ ( .D(N671), .CP(clk), .Q(
        i_data_bus_reg[636]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_635_ ( .D(N670), .CP(clk), .Q(
        i_data_bus_reg[635]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_634_ ( .D(N669), .CP(clk), .Q(
        i_data_bus_reg[634]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_633_ ( .D(N668), .CP(clk), .Q(
        i_data_bus_reg[633]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_632_ ( .D(N667), .CP(clk), .Q(
        i_data_bus_reg[632]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_631_ ( .D(N666), .CP(clk), .Q(
        i_data_bus_reg[631]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_630_ ( .D(N665), .CP(clk), .Q(
        i_data_bus_reg[630]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_629_ ( .D(N664), .CP(clk), .Q(
        i_data_bus_reg[629]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_628_ ( .D(N663), .CP(clk), .Q(
        i_data_bus_reg[628]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_627_ ( .D(N662), .CP(clk), .Q(
        i_data_bus_reg[627]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_626_ ( .D(N661), .CP(clk), .Q(
        i_data_bus_reg[626]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_625_ ( .D(N660), .CP(clk), .Q(
        i_data_bus_reg[625]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_624_ ( .D(N659), .CP(clk), .Q(
        i_data_bus_reg[624]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_623_ ( .D(N658), .CP(clk), .Q(
        i_data_bus_reg[623]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_622_ ( .D(N657), .CP(clk), .Q(
        i_data_bus_reg[622]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_621_ ( .D(N656), .CP(clk), .Q(
        i_data_bus_reg[621]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_620_ ( .D(N655), .CP(clk), .Q(
        i_data_bus_reg[620]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_619_ ( .D(N654), .CP(clk), .Q(
        i_data_bus_reg[619]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_618_ ( .D(N653), .CP(clk), .Q(
        i_data_bus_reg[618]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_617_ ( .D(N652), .CP(clk), .Q(
        i_data_bus_reg[617]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_616_ ( .D(N651), .CP(clk), .Q(
        i_data_bus_reg[616]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_615_ ( .D(N650), .CP(clk), .Q(
        i_data_bus_reg[615]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_614_ ( .D(N649), .CP(clk), .Q(
        i_data_bus_reg[614]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_613_ ( .D(N648), .CP(clk), .Q(
        i_data_bus_reg[613]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_612_ ( .D(N647), .CP(clk), .Q(
        i_data_bus_reg[612]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_611_ ( .D(N646), .CP(clk), .Q(
        i_data_bus_reg[611]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_610_ ( .D(N645), .CP(clk), .Q(
        i_data_bus_reg[610]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_609_ ( .D(N644), .CP(clk), .Q(
        i_data_bus_reg[609]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_608_ ( .D(N643), .CP(clk), .Q(
        i_data_bus_reg[608]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_607_ ( .D(N642), .CP(clk), .Q(
        i_data_bus_reg[607]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_606_ ( .D(N641), .CP(clk), .Q(
        i_data_bus_reg[606]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_605_ ( .D(N640), .CP(clk), .Q(
        i_data_bus_reg[605]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_604_ ( .D(N639), .CP(clk), .Q(
        i_data_bus_reg[604]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_603_ ( .D(N638), .CP(clk), .Q(
        i_data_bus_reg[603]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_602_ ( .D(N637), .CP(clk), .Q(
        i_data_bus_reg[602]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_601_ ( .D(N636), .CP(clk), .Q(
        i_data_bus_reg[601]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_600_ ( .D(N635), .CP(clk), .Q(
        i_data_bus_reg[600]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_599_ ( .D(N634), .CP(clk), .Q(
        i_data_bus_reg[599]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_598_ ( .D(N633), .CP(clk), .Q(
        i_data_bus_reg[598]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_597_ ( .D(N632), .CP(clk), .Q(
        i_data_bus_reg[597]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_596_ ( .D(N631), .CP(clk), .Q(
        i_data_bus_reg[596]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_595_ ( .D(N630), .CP(clk), .Q(
        i_data_bus_reg[595]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_594_ ( .D(N629), .CP(clk), .Q(
        i_data_bus_reg[594]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_593_ ( .D(N628), .CP(clk), .Q(
        i_data_bus_reg[593]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_592_ ( .D(N627), .CP(clk), .Q(
        i_data_bus_reg[592]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_591_ ( .D(N626), .CP(clk), .Q(
        i_data_bus_reg[591]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_590_ ( .D(N625), .CP(clk), .Q(
        i_data_bus_reg[590]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_589_ ( .D(N624), .CP(clk), .Q(
        i_data_bus_reg[589]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_588_ ( .D(N623), .CP(clk), .Q(
        i_data_bus_reg[588]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_587_ ( .D(N622), .CP(clk), .Q(
        i_data_bus_reg[587]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_586_ ( .D(N621), .CP(clk), .Q(
        i_data_bus_reg[586]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_585_ ( .D(N620), .CP(clk), .Q(
        i_data_bus_reg[585]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_584_ ( .D(N619), .CP(clk), .Q(
        i_data_bus_reg[584]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_583_ ( .D(N618), .CP(clk), .Q(
        i_data_bus_reg[583]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_582_ ( .D(N617), .CP(clk), .Q(
        i_data_bus_reg[582]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_581_ ( .D(N616), .CP(clk), .Q(
        i_data_bus_reg[581]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_580_ ( .D(N615), .CP(clk), .Q(
        i_data_bus_reg[580]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_579_ ( .D(N614), .CP(clk), .Q(
        i_data_bus_reg[579]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_578_ ( .D(N613), .CP(clk), .Q(
        i_data_bus_reg[578]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_577_ ( .D(N612), .CP(clk), .Q(
        i_data_bus_reg[577]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_576_ ( .D(N611), .CP(clk), .Q(
        i_data_bus_reg[576]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_575_ ( .D(N610), .CP(clk), .Q(
        i_data_bus_reg[575]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_574_ ( .D(N609), .CP(clk), .Q(
        i_data_bus_reg[574]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_573_ ( .D(N608), .CP(clk), .Q(
        i_data_bus_reg[573]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_572_ ( .D(N607), .CP(clk), .Q(
        i_data_bus_reg[572]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_571_ ( .D(N606), .CP(clk), .Q(
        i_data_bus_reg[571]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_570_ ( .D(N605), .CP(clk), .Q(
        i_data_bus_reg[570]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_569_ ( .D(N604), .CP(clk), .Q(
        i_data_bus_reg[569]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_568_ ( .D(N603), .CP(clk), .Q(
        i_data_bus_reg[568]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_567_ ( .D(N602), .CP(clk), .Q(
        i_data_bus_reg[567]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_566_ ( .D(N601), .CP(clk), .Q(
        i_data_bus_reg[566]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_565_ ( .D(N600), .CP(clk), .Q(
        i_data_bus_reg[565]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_564_ ( .D(N599), .CP(clk), .Q(
        i_data_bus_reg[564]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_563_ ( .D(N598), .CP(clk), .Q(
        i_data_bus_reg[563]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_562_ ( .D(N597), .CP(clk), .Q(
        i_data_bus_reg[562]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_561_ ( .D(N596), .CP(clk), .Q(
        i_data_bus_reg[561]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_560_ ( .D(N595), .CP(clk), .Q(
        i_data_bus_reg[560]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_559_ ( .D(N594), .CP(clk), .Q(
        i_data_bus_reg[559]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_558_ ( .D(N593), .CP(clk), .Q(
        i_data_bus_reg[558]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_557_ ( .D(N592), .CP(clk), .Q(
        i_data_bus_reg[557]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_556_ ( .D(N591), .CP(clk), .Q(
        i_data_bus_reg[556]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_555_ ( .D(N590), .CP(clk), .Q(
        i_data_bus_reg[555]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_554_ ( .D(N589), .CP(clk), .Q(
        i_data_bus_reg[554]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_553_ ( .D(N588), .CP(clk), .Q(
        i_data_bus_reg[553]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_552_ ( .D(N587), .CP(clk), .Q(
        i_data_bus_reg[552]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_551_ ( .D(N586), .CP(clk), .Q(
        i_data_bus_reg[551]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_550_ ( .D(N585), .CP(clk), .Q(
        i_data_bus_reg[550]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_549_ ( .D(N584), .CP(clk), .Q(
        i_data_bus_reg[549]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_548_ ( .D(N583), .CP(clk), .Q(
        i_data_bus_reg[548]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_547_ ( .D(N582), .CP(clk), .Q(
        i_data_bus_reg[547]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_546_ ( .D(N581), .CP(clk), .Q(
        i_data_bus_reg[546]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_545_ ( .D(N580), .CP(clk), .Q(
        i_data_bus_reg[545]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_544_ ( .D(N579), .CP(clk), .Q(
        i_data_bus_reg[544]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_543_ ( .D(N578), .CP(clk), .Q(
        i_data_bus_reg[543]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_542_ ( .D(N577), .CP(clk), .Q(
        i_data_bus_reg[542]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_541_ ( .D(N576), .CP(clk), .Q(
        i_data_bus_reg[541]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_540_ ( .D(N575), .CP(clk), .Q(
        i_data_bus_reg[540]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_539_ ( .D(N574), .CP(clk), .Q(
        i_data_bus_reg[539]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_538_ ( .D(N573), .CP(clk), .Q(
        i_data_bus_reg[538]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_537_ ( .D(N572), .CP(clk), .Q(
        i_data_bus_reg[537]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_536_ ( .D(N571), .CP(clk), .Q(
        i_data_bus_reg[536]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_535_ ( .D(N570), .CP(clk), .Q(
        i_data_bus_reg[535]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_534_ ( .D(N569), .CP(clk), .Q(
        i_data_bus_reg[534]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_533_ ( .D(N568), .CP(clk), .Q(
        i_data_bus_reg[533]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_532_ ( .D(N567), .CP(clk), .Q(
        i_data_bus_reg[532]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_531_ ( .D(N566), .CP(clk), .Q(
        i_data_bus_reg[531]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_530_ ( .D(N565), .CP(clk), .Q(
        i_data_bus_reg[530]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_529_ ( .D(N564), .CP(clk), .Q(
        i_data_bus_reg[529]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_528_ ( .D(N563), .CP(clk), .Q(
        i_data_bus_reg[528]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_527_ ( .D(N562), .CP(clk), .Q(
        i_data_bus_reg[527]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_526_ ( .D(N561), .CP(clk), .Q(
        i_data_bus_reg[526]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_525_ ( .D(N560), .CP(clk), .Q(
        i_data_bus_reg[525]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_524_ ( .D(N559), .CP(clk), .Q(
        i_data_bus_reg[524]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_523_ ( .D(N558), .CP(clk), .Q(
        i_data_bus_reg[523]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_522_ ( .D(N557), .CP(clk), .Q(
        i_data_bus_reg[522]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_521_ ( .D(N556), .CP(clk), .Q(
        i_data_bus_reg[521]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_520_ ( .D(N555), .CP(clk), .Q(
        i_data_bus_reg[520]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_519_ ( .D(N554), .CP(clk), .Q(
        i_data_bus_reg[519]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_518_ ( .D(N553), .CP(clk), .Q(
        i_data_bus_reg[518]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_517_ ( .D(N552), .CP(clk), .Q(
        i_data_bus_reg[517]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_516_ ( .D(N551), .CP(clk), .Q(
        i_data_bus_reg[516]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_515_ ( .D(N550), .CP(clk), .Q(
        i_data_bus_reg[515]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_514_ ( .D(N549), .CP(clk), .Q(
        i_data_bus_reg[514]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_513_ ( .D(N548), .CP(clk), .Q(
        i_data_bus_reg[513]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_512_ ( .D(N547), .CP(clk), .Q(
        i_data_bus_reg[512]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_511_ ( .D(N546), .CP(clk), .Q(
        i_data_bus_reg[511]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_510_ ( .D(N545), .CP(clk), .Q(
        i_data_bus_reg[510]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_509_ ( .D(N544), .CP(clk), .Q(
        i_data_bus_reg[509]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_508_ ( .D(N543), .CP(clk), .Q(
        i_data_bus_reg[508]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_507_ ( .D(N542), .CP(clk), .Q(
        i_data_bus_reg[507]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_506_ ( .D(N541), .CP(clk), .Q(
        i_data_bus_reg[506]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_505_ ( .D(N540), .CP(clk), .Q(
        i_data_bus_reg[505]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_504_ ( .D(N539), .CP(clk), .Q(
        i_data_bus_reg[504]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_503_ ( .D(N538), .CP(clk), .Q(
        i_data_bus_reg[503]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_502_ ( .D(N537), .CP(clk), .Q(
        i_data_bus_reg[502]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_501_ ( .D(N536), .CP(clk), .Q(
        i_data_bus_reg[501]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_500_ ( .D(N535), .CP(clk), .Q(
        i_data_bus_reg[500]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_499_ ( .D(N534), .CP(clk), .Q(
        i_data_bus_reg[499]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_498_ ( .D(N533), .CP(clk), .Q(
        i_data_bus_reg[498]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_497_ ( .D(N532), .CP(clk), .Q(
        i_data_bus_reg[497]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_496_ ( .D(N531), .CP(clk), .Q(
        i_data_bus_reg[496]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_495_ ( .D(N530), .CP(clk), .Q(
        i_data_bus_reg[495]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_494_ ( .D(N529), .CP(clk), .Q(
        i_data_bus_reg[494]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_493_ ( .D(N528), .CP(clk), .Q(
        i_data_bus_reg[493]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_492_ ( .D(N527), .CP(clk), .Q(
        i_data_bus_reg[492]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_491_ ( .D(N526), .CP(clk), .Q(
        i_data_bus_reg[491]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_490_ ( .D(N525), .CP(clk), .Q(
        i_data_bus_reg[490]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_489_ ( .D(N524), .CP(clk), .Q(
        i_data_bus_reg[489]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_488_ ( .D(N523), .CP(clk), .Q(
        i_data_bus_reg[488]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_487_ ( .D(N522), .CP(clk), .Q(
        i_data_bus_reg[487]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_486_ ( .D(N521), .CP(clk), .Q(
        i_data_bus_reg[486]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_485_ ( .D(N520), .CP(clk), .Q(
        i_data_bus_reg[485]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_484_ ( .D(N519), .CP(clk), .Q(
        i_data_bus_reg[484]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_483_ ( .D(N518), .CP(clk), .Q(
        i_data_bus_reg[483]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_482_ ( .D(N517), .CP(clk), .Q(
        i_data_bus_reg[482]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_481_ ( .D(N516), .CP(clk), .Q(
        i_data_bus_reg[481]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_480_ ( .D(N515), .CP(clk), .Q(
        i_data_bus_reg[480]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_479_ ( .D(N514), .CP(clk), .Q(
        i_data_bus_reg[479]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_478_ ( .D(N513), .CP(clk), .Q(
        i_data_bus_reg[478]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_477_ ( .D(N512), .CP(clk), .Q(
        i_data_bus_reg[477]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_476_ ( .D(N511), .CP(clk), .Q(
        i_data_bus_reg[476]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_475_ ( .D(N510), .CP(clk), .Q(
        i_data_bus_reg[475]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_474_ ( .D(N509), .CP(clk), .Q(
        i_data_bus_reg[474]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_473_ ( .D(N508), .CP(clk), .Q(
        i_data_bus_reg[473]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_472_ ( .D(N507), .CP(clk), .Q(
        i_data_bus_reg[472]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_471_ ( .D(N506), .CP(clk), .Q(
        i_data_bus_reg[471]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_470_ ( .D(N505), .CP(clk), .Q(
        i_data_bus_reg[470]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_469_ ( .D(N504), .CP(clk), .Q(
        i_data_bus_reg[469]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_468_ ( .D(N503), .CP(clk), .Q(
        i_data_bus_reg[468]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_467_ ( .D(N502), .CP(clk), .Q(
        i_data_bus_reg[467]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_466_ ( .D(N501), .CP(clk), .Q(
        i_data_bus_reg[466]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_465_ ( .D(N500), .CP(clk), .Q(
        i_data_bus_reg[465]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_464_ ( .D(N499), .CP(clk), .Q(
        i_data_bus_reg[464]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_463_ ( .D(N498), .CP(clk), .Q(
        i_data_bus_reg[463]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_462_ ( .D(N497), .CP(clk), .Q(
        i_data_bus_reg[462]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_461_ ( .D(N496), .CP(clk), .Q(
        i_data_bus_reg[461]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_460_ ( .D(N495), .CP(clk), .Q(
        i_data_bus_reg[460]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_459_ ( .D(N494), .CP(clk), .Q(
        i_data_bus_reg[459]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_458_ ( .D(N493), .CP(clk), .Q(
        i_data_bus_reg[458]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_457_ ( .D(N492), .CP(clk), .Q(
        i_data_bus_reg[457]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_456_ ( .D(N491), .CP(clk), .Q(
        i_data_bus_reg[456]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_455_ ( .D(N490), .CP(clk), .Q(
        i_data_bus_reg[455]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_454_ ( .D(N489), .CP(clk), .Q(
        i_data_bus_reg[454]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_453_ ( .D(N488), .CP(clk), .Q(
        i_data_bus_reg[453]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_452_ ( .D(N487), .CP(clk), .Q(
        i_data_bus_reg[452]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_451_ ( .D(N486), .CP(clk), .Q(
        i_data_bus_reg[451]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_450_ ( .D(N485), .CP(clk), .Q(
        i_data_bus_reg[450]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_449_ ( .D(N484), .CP(clk), .Q(
        i_data_bus_reg[449]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_448_ ( .D(N483), .CP(clk), .Q(
        i_data_bus_reg[448]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_447_ ( .D(N482), .CP(clk), .Q(
        i_data_bus_reg[447]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_446_ ( .D(N481), .CP(clk), .Q(
        i_data_bus_reg[446]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_445_ ( .D(N480), .CP(clk), .Q(
        i_data_bus_reg[445]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_444_ ( .D(N479), .CP(clk), .Q(
        i_data_bus_reg[444]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_443_ ( .D(N478), .CP(clk), .Q(
        i_data_bus_reg[443]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_442_ ( .D(N477), .CP(clk), .Q(
        i_data_bus_reg[442]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_441_ ( .D(N476), .CP(clk), .Q(
        i_data_bus_reg[441]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_440_ ( .D(N475), .CP(clk), .Q(
        i_data_bus_reg[440]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_439_ ( .D(N474), .CP(clk), .Q(
        i_data_bus_reg[439]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_438_ ( .D(N473), .CP(clk), .Q(
        i_data_bus_reg[438]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_437_ ( .D(N472), .CP(clk), .Q(
        i_data_bus_reg[437]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_436_ ( .D(N471), .CP(clk), .Q(
        i_data_bus_reg[436]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_435_ ( .D(N470), .CP(clk), .Q(
        i_data_bus_reg[435]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_434_ ( .D(N469), .CP(clk), .Q(
        i_data_bus_reg[434]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_433_ ( .D(N468), .CP(clk), .Q(
        i_data_bus_reg[433]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_432_ ( .D(N467), .CP(clk), .Q(
        i_data_bus_reg[432]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_431_ ( .D(N466), .CP(clk), .Q(
        i_data_bus_reg[431]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_430_ ( .D(N465), .CP(clk), .Q(
        i_data_bus_reg[430]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_429_ ( .D(N464), .CP(clk), .Q(
        i_data_bus_reg[429]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_428_ ( .D(N463), .CP(clk), .Q(
        i_data_bus_reg[428]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_427_ ( .D(N462), .CP(clk), .Q(
        i_data_bus_reg[427]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_426_ ( .D(N461), .CP(clk), .Q(
        i_data_bus_reg[426]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_425_ ( .D(N460), .CP(clk), .Q(
        i_data_bus_reg[425]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_424_ ( .D(N459), .CP(clk), .Q(
        i_data_bus_reg[424]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_423_ ( .D(N458), .CP(clk), .Q(
        i_data_bus_reg[423]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_422_ ( .D(N457), .CP(clk), .Q(
        i_data_bus_reg[422]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_421_ ( .D(N456), .CP(clk), .Q(
        i_data_bus_reg[421]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_420_ ( .D(N455), .CP(clk), .Q(
        i_data_bus_reg[420]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_419_ ( .D(N454), .CP(clk), .Q(
        i_data_bus_reg[419]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_418_ ( .D(N453), .CP(clk), .Q(
        i_data_bus_reg[418]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_417_ ( .D(N452), .CP(clk), .Q(
        i_data_bus_reg[417]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_416_ ( .D(N451), .CP(clk), .Q(
        i_data_bus_reg[416]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_415_ ( .D(N450), .CP(clk), .Q(
        i_data_bus_reg[415]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_414_ ( .D(N449), .CP(clk), .Q(
        i_data_bus_reg[414]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_413_ ( .D(N448), .CP(clk), .Q(
        i_data_bus_reg[413]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_412_ ( .D(N447), .CP(clk), .Q(
        i_data_bus_reg[412]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_411_ ( .D(N446), .CP(clk), .Q(
        i_data_bus_reg[411]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_410_ ( .D(N445), .CP(clk), .Q(
        i_data_bus_reg[410]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_409_ ( .D(N444), .CP(clk), .Q(
        i_data_bus_reg[409]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_408_ ( .D(N443), .CP(clk), .Q(
        i_data_bus_reg[408]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_407_ ( .D(N442), .CP(clk), .Q(
        i_data_bus_reg[407]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_406_ ( .D(N441), .CP(clk), .Q(
        i_data_bus_reg[406]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_405_ ( .D(N440), .CP(clk), .Q(
        i_data_bus_reg[405]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_404_ ( .D(N439), .CP(clk), .Q(
        i_data_bus_reg[404]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_403_ ( .D(N438), .CP(clk), .Q(
        i_data_bus_reg[403]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_402_ ( .D(N437), .CP(clk), .Q(
        i_data_bus_reg[402]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_401_ ( .D(N436), .CP(clk), .Q(
        i_data_bus_reg[401]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_400_ ( .D(N435), .CP(clk), .Q(
        i_data_bus_reg[400]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_399_ ( .D(N434), .CP(clk), .Q(
        i_data_bus_reg[399]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_398_ ( .D(N433), .CP(clk), .Q(
        i_data_bus_reg[398]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_397_ ( .D(N432), .CP(clk), .Q(
        i_data_bus_reg[397]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_396_ ( .D(N431), .CP(clk), .Q(
        i_data_bus_reg[396]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_395_ ( .D(N430), .CP(clk), .Q(
        i_data_bus_reg[395]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_394_ ( .D(N429), .CP(clk), .Q(
        i_data_bus_reg[394]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_393_ ( .D(N428), .CP(clk), .Q(
        i_data_bus_reg[393]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_392_ ( .D(N427), .CP(clk), .Q(
        i_data_bus_reg[392]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_391_ ( .D(N426), .CP(clk), .Q(
        i_data_bus_reg[391]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_390_ ( .D(N425), .CP(clk), .Q(
        i_data_bus_reg[390]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_389_ ( .D(N424), .CP(clk), .Q(
        i_data_bus_reg[389]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_388_ ( .D(N423), .CP(clk), .Q(
        i_data_bus_reg[388]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_387_ ( .D(N422), .CP(clk), .Q(
        i_data_bus_reg[387]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_386_ ( .D(N421), .CP(clk), .Q(
        i_data_bus_reg[386]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_385_ ( .D(N420), .CP(clk), .Q(
        i_data_bus_reg[385]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_384_ ( .D(N419), .CP(clk), .Q(
        i_data_bus_reg[384]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_383_ ( .D(N418), .CP(clk), .Q(
        i_data_bus_reg[383]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_382_ ( .D(N417), .CP(clk), .Q(
        i_data_bus_reg[382]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_381_ ( .D(N416), .CP(clk), .Q(
        i_data_bus_reg[381]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_380_ ( .D(N415), .CP(clk), .Q(
        i_data_bus_reg[380]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_379_ ( .D(N414), .CP(clk), .Q(
        i_data_bus_reg[379]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_378_ ( .D(N413), .CP(clk), .Q(
        i_data_bus_reg[378]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_377_ ( .D(N412), .CP(clk), .Q(
        i_data_bus_reg[377]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_376_ ( .D(N411), .CP(clk), .Q(
        i_data_bus_reg[376]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_375_ ( .D(N410), .CP(clk), .Q(
        i_data_bus_reg[375]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_374_ ( .D(N409), .CP(clk), .Q(
        i_data_bus_reg[374]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_373_ ( .D(N408), .CP(clk), .Q(
        i_data_bus_reg[373]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_372_ ( .D(N407), .CP(clk), .Q(
        i_data_bus_reg[372]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_371_ ( .D(N406), .CP(clk), .Q(
        i_data_bus_reg[371]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_370_ ( .D(N405), .CP(clk), .Q(
        i_data_bus_reg[370]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_369_ ( .D(N404), .CP(clk), .Q(
        i_data_bus_reg[369]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_368_ ( .D(N403), .CP(clk), .Q(
        i_data_bus_reg[368]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_367_ ( .D(N402), .CP(clk), .Q(
        i_data_bus_reg[367]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_366_ ( .D(N401), .CP(clk), .Q(
        i_data_bus_reg[366]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_365_ ( .D(N400), .CP(clk), .Q(
        i_data_bus_reg[365]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_364_ ( .D(N399), .CP(clk), .Q(
        i_data_bus_reg[364]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_363_ ( .D(N398), .CP(clk), .Q(
        i_data_bus_reg[363]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_362_ ( .D(N397), .CP(clk), .Q(
        i_data_bus_reg[362]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_361_ ( .D(N396), .CP(clk), .Q(
        i_data_bus_reg[361]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_360_ ( .D(N395), .CP(clk), .Q(
        i_data_bus_reg[360]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_359_ ( .D(N394), .CP(clk), .Q(
        i_data_bus_reg[359]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_358_ ( .D(N393), .CP(clk), .Q(
        i_data_bus_reg[358]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_357_ ( .D(N392), .CP(clk), .Q(
        i_data_bus_reg[357]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_356_ ( .D(N391), .CP(clk), .Q(
        i_data_bus_reg[356]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_355_ ( .D(N390), .CP(clk), .Q(
        i_data_bus_reg[355]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_354_ ( .D(N389), .CP(clk), .Q(
        i_data_bus_reg[354]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_353_ ( .D(N388), .CP(clk), .Q(
        i_data_bus_reg[353]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_352_ ( .D(N387), .CP(clk), .Q(
        i_data_bus_reg[352]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_351_ ( .D(N386), .CP(clk), .Q(
        i_data_bus_reg[351]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_350_ ( .D(N385), .CP(clk), .Q(
        i_data_bus_reg[350]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_349_ ( .D(N384), .CP(clk), .Q(
        i_data_bus_reg[349]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_348_ ( .D(N383), .CP(clk), .Q(
        i_data_bus_reg[348]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_347_ ( .D(N382), .CP(clk), .Q(
        i_data_bus_reg[347]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_346_ ( .D(N381), .CP(clk), .Q(
        i_data_bus_reg[346]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_345_ ( .D(N380), .CP(clk), .Q(
        i_data_bus_reg[345]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_344_ ( .D(N379), .CP(clk), .Q(
        i_data_bus_reg[344]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_343_ ( .D(N378), .CP(clk), .Q(
        i_data_bus_reg[343]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_342_ ( .D(N377), .CP(clk), .Q(
        i_data_bus_reg[342]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_341_ ( .D(N376), .CP(clk), .Q(
        i_data_bus_reg[341]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_340_ ( .D(N375), .CP(clk), .Q(
        i_data_bus_reg[340]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_339_ ( .D(N374), .CP(clk), .Q(
        i_data_bus_reg[339]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_338_ ( .D(N373), .CP(clk), .Q(
        i_data_bus_reg[338]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_337_ ( .D(N372), .CP(clk), .Q(
        i_data_bus_reg[337]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_336_ ( .D(N371), .CP(clk), .Q(
        i_data_bus_reg[336]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_335_ ( .D(N370), .CP(clk), .Q(
        i_data_bus_reg[335]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_334_ ( .D(N369), .CP(clk), .Q(
        i_data_bus_reg[334]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_333_ ( .D(N368), .CP(clk), .Q(
        i_data_bus_reg[333]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_332_ ( .D(N367), .CP(clk), .Q(
        i_data_bus_reg[332]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_331_ ( .D(N366), .CP(clk), .Q(
        i_data_bus_reg[331]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_330_ ( .D(N365), .CP(clk), .Q(
        i_data_bus_reg[330]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_329_ ( .D(N364), .CP(clk), .Q(
        i_data_bus_reg[329]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_328_ ( .D(N363), .CP(clk), .Q(
        i_data_bus_reg[328]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_327_ ( .D(N362), .CP(clk), .Q(
        i_data_bus_reg[327]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_326_ ( .D(N361), .CP(clk), .Q(
        i_data_bus_reg[326]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_325_ ( .D(N360), .CP(clk), .Q(
        i_data_bus_reg[325]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_324_ ( .D(N359), .CP(clk), .Q(
        i_data_bus_reg[324]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_323_ ( .D(N358), .CP(clk), .Q(
        i_data_bus_reg[323]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_322_ ( .D(N357), .CP(clk), .Q(
        i_data_bus_reg[322]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_321_ ( .D(N356), .CP(clk), .Q(
        i_data_bus_reg[321]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_320_ ( .D(N355), .CP(clk), .Q(
        i_data_bus_reg[320]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_319_ ( .D(N354), .CP(clk), .Q(
        i_data_bus_reg[319]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_318_ ( .D(N353), .CP(clk), .Q(
        i_data_bus_reg[318]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_317_ ( .D(N352), .CP(clk), .Q(
        i_data_bus_reg[317]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_316_ ( .D(N351), .CP(clk), .Q(
        i_data_bus_reg[316]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_315_ ( .D(N350), .CP(clk), .Q(
        i_data_bus_reg[315]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_314_ ( .D(N349), .CP(clk), .Q(
        i_data_bus_reg[314]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_313_ ( .D(N348), .CP(clk), .Q(
        i_data_bus_reg[313]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_312_ ( .D(N347), .CP(clk), .Q(
        i_data_bus_reg[312]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_311_ ( .D(N346), .CP(clk), .Q(
        i_data_bus_reg[311]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_310_ ( .D(N345), .CP(clk), .Q(
        i_data_bus_reg[310]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_309_ ( .D(N344), .CP(clk), .Q(
        i_data_bus_reg[309]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_308_ ( .D(N343), .CP(clk), .Q(
        i_data_bus_reg[308]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_300_ ( .D(N335), .CP(clk), .Q(
        i_data_bus_reg[300]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_299_ ( .D(N334), .CP(clk), .Q(
        i_data_bus_reg[299]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_298_ ( .D(N333), .CP(clk), .Q(
        i_data_bus_reg[298]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_297_ ( .D(N332), .CP(clk), .Q(
        i_data_bus_reg[297]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_296_ ( .D(N331), .CP(clk), .Q(
        i_data_bus_reg[296]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_291_ ( .D(N326), .CP(clk), .Q(
        i_data_bus_reg[291]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_290_ ( .D(N325), .CP(clk), .Q(
        i_data_bus_reg[290]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_289_ ( .D(N324), .CP(clk), .Q(
        i_data_bus_reg[289]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_288_ ( .D(N323), .CP(clk), .Q(
        i_data_bus_reg[288]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_287_ ( .D(N322), .CP(clk), .Q(
        i_data_bus_reg[287]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_286_ ( .D(N321), .CP(clk), .Q(
        i_data_bus_reg[286]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_285_ ( .D(N320), .CP(clk), .Q(
        i_data_bus_reg[285]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_284_ ( .D(N319), .CP(clk), .Q(
        i_data_bus_reg[284]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_228_ ( .D(N263), .CP(clk), .Q(
        i_data_bus_reg[228]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_227_ ( .D(N262), .CP(clk), .Q(
        i_data_bus_reg[227]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_226_ ( .D(N261), .CP(clk), .Q(
        i_data_bus_reg[226]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_225_ ( .D(N260), .CP(clk), .Q(
        i_data_bus_reg[225]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_224_ ( .D(N259), .CP(clk), .Q(
        i_data_bus_reg[224]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_219_ ( .D(N254), .CP(clk), .Q(
        i_data_bus_reg[219]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_218_ ( .D(N253), .CP(clk), .Q(
        i_data_bus_reg[218]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_217_ ( .D(N252), .CP(clk), .Q(
        i_data_bus_reg[217]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_216_ ( .D(N251), .CP(clk), .Q(
        i_data_bus_reg[216]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_215_ ( .D(N250), .CP(clk), .Q(
        i_data_bus_reg[215]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_214_ ( .D(N249), .CP(clk), .Q(
        i_data_bus_reg[214]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_213_ ( .D(N248), .CP(clk), .Q(
        i_data_bus_reg[213]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_212_ ( .D(N247), .CP(clk), .Q(
        i_data_bus_reg[212]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_156_ ( .D(N191), .CP(clk), .Q(
        i_data_bus_reg[156]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_155_ ( .D(N190), .CP(clk), .Q(
        i_data_bus_reg[155]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_154_ ( .D(N189), .CP(clk), .Q(
        i_data_bus_reg[154]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_153_ ( .D(N188), .CP(clk), .Q(
        i_data_bus_reg[153]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_152_ ( .D(N187), .CP(clk), .Q(
        i_data_bus_reg[152]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_147_ ( .D(N182), .CP(clk), .Q(
        i_data_bus_reg[147]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_146_ ( .D(N181), .CP(clk), .Q(
        i_data_bus_reg[146]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_145_ ( .D(N180), .CP(clk), .Q(
        i_data_bus_reg[145]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_144_ ( .D(N179), .CP(clk), .Q(
        i_data_bus_reg[144]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_143_ ( .D(N178), .CP(clk), .Q(
        i_data_bus_reg[143]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_142_ ( .D(N177), .CP(clk), .Q(
        i_data_bus_reg[142]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_141_ ( .D(N176), .CP(clk), .Q(
        i_data_bus_reg[141]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_140_ ( .D(N175), .CP(clk), .Q(
        i_data_bus_reg[140]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_127_ ( .D(N162), .CP(clk), .Q(
        i_data_bus_reg[127]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_126_ ( .D(N161), .CP(clk), .Q(
        i_data_bus_reg[126]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_125_ ( .D(N160), .CP(clk), .Q(
        i_data_bus_reg[125]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_124_ ( .D(N159), .CP(clk), .Q(
        i_data_bus_reg[124]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_123_ ( .D(N158), .CP(clk), .Q(
        i_data_bus_reg[123]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_122_ ( .D(N157), .CP(clk), .Q(
        i_data_bus_reg[122]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_121_ ( .D(N156), .CP(clk), .Q(
        i_data_bus_reg[121]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_120_ ( .D(N155), .CP(clk), .Q(
        i_data_bus_reg[120]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_119_ ( .D(N154), .CP(clk), .Q(
        i_data_bus_reg[119]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_118_ ( .D(N153), .CP(clk), .Q(
        i_data_bus_reg[118]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_117_ ( .D(N152), .CP(clk), .Q(
        i_data_bus_reg[117]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_116_ ( .D(N151), .CP(clk), .Q(
        i_data_bus_reg[116]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_110_ ( .D(N145), .CP(clk), .Q(
        i_data_bus_reg[110]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_109_ ( .D(N144), .CP(clk), .Q(
        i_data_bus_reg[109]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_108_ ( .D(N143), .CP(clk), .Q(
        i_data_bus_reg[108]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_107_ ( .D(N142), .CP(clk), .Q(
        i_data_bus_reg[107]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_106_ ( .D(N141), .CP(clk), .Q(
        i_data_bus_reg[106]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_105_ ( .D(N140), .CP(clk), .Q(
        i_data_bus_reg[105]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_104_ ( .D(N139), .CP(clk), .Q(
        i_data_bus_reg[104]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_103_ ( .D(N138), .CP(clk), .Q(
        i_data_bus_reg[103]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_102_ ( .D(N137), .CP(clk), .Q(
        i_data_bus_reg[102]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_101_ ( .D(N136), .CP(clk), .Q(
        i_data_bus_reg[101]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_100_ ( .D(N135), .CP(clk), .Q(
        i_data_bus_reg[100]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_99_ ( .D(N134), .CP(clk), .Q(
        i_data_bus_reg[99]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_98_ ( .D(N133), .CP(clk), .Q(
        i_data_bus_reg[98]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_97_ ( .D(N132), .CP(clk), .Q(
        i_data_bus_reg[97]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_96_ ( .D(N131), .CP(clk), .Q(
        i_data_bus_reg[96]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_95_ ( .D(N130), .CP(clk), .Q(
        i_data_bus_reg[95]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_94_ ( .D(N129), .CP(clk), .Q(
        i_data_bus_reg[94]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_93_ ( .D(N128), .CP(clk), .Q(
        i_data_bus_reg[93]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_92_ ( .D(N127), .CP(clk), .Q(
        i_data_bus_reg[92]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_84_ ( .D(N119), .CP(clk), .Q(
        i_data_bus_reg[84]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_83_ ( .D(N118), .CP(clk), .Q(
        i_data_bus_reg[83]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_82_ ( .D(N117), .CP(clk), .Q(
        i_data_bus_reg[82]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_81_ ( .D(N116), .CP(clk), .Q(
        i_data_bus_reg[81]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_80_ ( .D(N115), .CP(clk), .Q(
        i_data_bus_reg[80]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_75_ ( .D(N110), .CP(clk), .Q(
        i_data_bus_reg[75]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_74_ ( .D(N109), .CP(clk), .Q(
        i_data_bus_reg[74]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_73_ ( .D(N108), .CP(clk), .Q(
        i_data_bus_reg[73]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_72_ ( .D(N107), .CP(clk), .Q(
        i_data_bus_reg[72]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_71_ ( .D(N106), .CP(clk), .Q(
        i_data_bus_reg[71]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_70_ ( .D(N105), .CP(clk), .Q(
        i_data_bus_reg[70]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_69_ ( .D(N104), .CP(clk), .Q(
        i_data_bus_reg[69]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_68_ ( .D(N103), .CP(clk), .Q(
        i_data_bus_reg[68]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_32_ ( .D(N67), .CP(clk), .Q(
        i_data_bus_reg[32]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_31_ ( .D(N66), .CP(clk), .Q(
        i_data_bus_reg[31]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_30_ ( .D(N65), .CP(clk), .Q(
        i_data_bus_reg[30]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_29_ ( .D(N64), .CP(clk), .Q(
        i_data_bus_reg[29]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_28_ ( .D(N63), .CP(clk), .Q(
        i_data_bus_reg[28]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_27_ ( .D(N62), .CP(clk), .Q(
        i_data_bus_reg[27]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_26_ ( .D(N61), .CP(clk), .Q(
        i_data_bus_reg[26]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_24_ ( .D(N59), .CP(clk), .Q(
        i_data_bus_reg[24]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_23_ ( .D(N58), .CP(clk), .Q(
        i_data_bus_reg[23]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_22_ ( .D(N57), .CP(clk), .Q(
        i_data_bus_reg[22]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_21_ ( .D(N56), .CP(clk), .Q(
        i_data_bus_reg[21]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_20_ ( .D(N55), .CP(clk), .Q(
        i_data_bus_reg[20]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_19_ ( .D(N54), .CP(clk), .Q(
        i_data_bus_reg[19]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_18_ ( .D(N53), .CP(clk), .Q(
        i_data_bus_reg[18]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_17_ ( .D(N52), .CP(clk), .Q(
        i_data_bus_reg[17]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_16_ ( .D(N51), .CP(clk), .Q(
        i_data_bus_reg[16]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_15_ ( .D(N50), .CP(clk), .Q(
        i_data_bus_reg[15]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_14_ ( .D(N49), .CP(clk), .Q(
        i_data_bus_reg[14]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_13_ ( .D(N48), .CP(clk), .Q(
        i_data_bus_reg[13]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_12_ ( .D(N47), .CP(clk), .Q(
        i_data_bus_reg[12]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_11_ ( .D(N46), .CP(clk), .Q(
        i_data_bus_reg[11]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_10_ ( .D(N45), .CP(clk), .Q(
        i_data_bus_reg[10]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_9_ ( .D(N44), .CP(clk), .Q(
        i_data_bus_reg[9]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_8_ ( .D(N43), .CP(clk), .Q(
        i_data_bus_reg[8]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_7_ ( .D(N42), .CP(clk), .Q(
        i_data_bus_reg[7]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_6_ ( .D(N41), .CP(clk), .Q(
        i_data_bus_reg[6]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_5_ ( .D(N40), .CP(clk), .Q(
        i_data_bus_reg[5]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_4_ ( .D(N39), .CP(clk), .Q(
        i_data_bus_reg[4]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_3_ ( .D(N38), .CP(clk), .Q(
        i_data_bus_reg[3]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_2_ ( .D(N37), .CP(clk), .Q(
        i_data_bus_reg[2]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_1_ ( .D(N36), .CP(clk), .Q(
        i_data_bus_reg[1]) );
  DFQD1BWP30P140LVT i_data_bus_reg_reg_0_ ( .D(N35), .CP(clk), .Q(
        i_data_bus_reg[0]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_7_ ( .D(o_valid_wire[7]), .CP(clk), .Q(
        o_valid[7]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_6_ ( .D(o_valid_wire[6]), .CP(clk), .Q(
        o_valid[6]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_5_ ( .D(o_valid_wire[5]), .CP(clk), .Q(
        o_valid[5]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_4_ ( .D(o_valid_wire[4]), .CP(clk), .Q(
        o_valid[4]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_3_ ( .D(o_valid_wire[3]), .CP(clk), .Q(
        o_valid[3]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_2_ ( .D(o_valid_wire[2]), .CP(clk), .Q(
        o_valid[2]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_1_ ( .D(o_valid_wire[1]), .CP(clk), .Q(
        o_valid[1]) );
  DFQD2BWP30P140LVT o_valid_reg_reg_0_ ( .D(o_valid_wire[0]), .CP(clk), .Q(
        o_valid[0]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(o_data_bus_wire[255]), .CP(
        clk), .Q(o_data_bus[255]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(o_data_bus_wire[254]), .CP(
        clk), .Q(o_data_bus[254]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(o_data_bus_wire[253]), .CP(
        clk), .Q(o_data_bus[253]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(o_data_bus_wire[252]), .CP(
        clk), .Q(o_data_bus[252]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(o_data_bus_wire[251]), .CP(
        clk), .Q(o_data_bus[251]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(o_data_bus_wire[250]), .CP(
        clk), .Q(o_data_bus[250]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(o_data_bus_wire[249]), .CP(
        clk), .Q(o_data_bus[249]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(o_data_bus_wire[248]), .CP(
        clk), .Q(o_data_bus[248]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(o_data_bus_wire[247]), .CP(
        clk), .Q(o_data_bus[247]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(o_data_bus_wire[246]), .CP(
        clk), .Q(o_data_bus[246]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(o_data_bus_wire[245]), .CP(
        clk), .Q(o_data_bus[245]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(o_data_bus_wire[244]), .CP(
        clk), .Q(o_data_bus[244]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(o_data_bus_wire[243]), .CP(
        clk), .Q(o_data_bus[243]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(o_data_bus_wire[242]), .CP(
        clk), .Q(o_data_bus[242]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(o_data_bus_wire[241]), .CP(
        clk), .Q(o_data_bus[241]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(o_data_bus_wire[240]), .CP(
        clk), .Q(o_data_bus[240]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(o_data_bus_wire[239]), .CP(
        clk), .Q(o_data_bus[239]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(o_data_bus_wire[238]), .CP(
        clk), .Q(o_data_bus[238]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(o_data_bus_wire[237]), .CP(
        clk), .Q(o_data_bus[237]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(o_data_bus_wire[236]), .CP(
        clk), .Q(o_data_bus[236]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(o_data_bus_wire[235]), .CP(
        clk), .Q(o_data_bus[235]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(o_data_bus_wire[234]), .CP(
        clk), .Q(o_data_bus[234]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(o_data_bus_wire[233]), .CP(
        clk), .Q(o_data_bus[233]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(o_data_bus_wire[232]), .CP(
        clk), .Q(o_data_bus[232]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(o_data_bus_wire[231]), .CP(
        clk), .Q(o_data_bus[231]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(o_data_bus_wire[230]), .CP(
        clk), .Q(o_data_bus[230]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(o_data_bus_wire[229]), .CP(
        clk), .Q(o_data_bus[229]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(o_data_bus_wire[228]), .CP(
        clk), .Q(o_data_bus[228]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(o_data_bus_wire[227]), .CP(
        clk), .Q(o_data_bus[227]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(o_data_bus_wire[226]), .CP(
        clk), .Q(o_data_bus[226]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(o_data_bus_wire[225]), .CP(
        clk), .Q(o_data_bus[225]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(o_data_bus_wire[224]), .CP(
        clk), .Q(o_data_bus[224]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(o_data_bus_wire[223]), .CP(
        clk), .Q(o_data_bus[223]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(o_data_bus_wire[222]), .CP(
        clk), .Q(o_data_bus[222]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(o_data_bus_wire[221]), .CP(
        clk), .Q(o_data_bus[221]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(o_data_bus_wire[220]), .CP(
        clk), .Q(o_data_bus[220]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(o_data_bus_wire[219]), .CP(
        clk), .Q(o_data_bus[219]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(o_data_bus_wire[218]), .CP(
        clk), .Q(o_data_bus[218]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(o_data_bus_wire[217]), .CP(
        clk), .Q(o_data_bus[217]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(o_data_bus_wire[216]), .CP(
        clk), .Q(o_data_bus[216]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(o_data_bus_wire[215]), .CP(
        clk), .Q(o_data_bus[215]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(o_data_bus_wire[214]), .CP(
        clk), .Q(o_data_bus[214]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(o_data_bus_wire[213]), .CP(
        clk), .Q(o_data_bus[213]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(o_data_bus_wire[212]), .CP(
        clk), .Q(o_data_bus[212]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(o_data_bus_wire[211]), .CP(
        clk), .Q(o_data_bus[211]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(o_data_bus_wire[210]), .CP(
        clk), .Q(o_data_bus[210]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(o_data_bus_wire[209]), .CP(
        clk), .Q(o_data_bus[209]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(o_data_bus_wire[208]), .CP(
        clk), .Q(o_data_bus[208]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(o_data_bus_wire[207]), .CP(
        clk), .Q(o_data_bus[207]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(o_data_bus_wire[206]), .CP(
        clk), .Q(o_data_bus[206]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(o_data_bus_wire[205]), .CP(
        clk), .Q(o_data_bus[205]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(o_data_bus_wire[204]), .CP(
        clk), .Q(o_data_bus[204]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(o_data_bus_wire[203]), .CP(
        clk), .Q(o_data_bus[203]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(o_data_bus_wire[202]), .CP(
        clk), .Q(o_data_bus[202]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(o_data_bus_wire[201]), .CP(
        clk), .Q(o_data_bus[201]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(o_data_bus_wire[200]), .CP(
        clk), .Q(o_data_bus[200]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(o_data_bus_wire[199]), .CP(
        clk), .Q(o_data_bus[199]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(o_data_bus_wire[198]), .CP(
        clk), .Q(o_data_bus[198]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(o_data_bus_wire[197]), .CP(
        clk), .Q(o_data_bus[197]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(o_data_bus_wire[196]), .CP(
        clk), .Q(o_data_bus[196]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(o_data_bus_wire[195]), .CP(
        clk), .Q(o_data_bus[195]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(o_data_bus_wire[194]), .CP(
        clk), .Q(o_data_bus[194]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(o_data_bus_wire[193]), .CP(
        clk), .Q(o_data_bus[193]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(o_data_bus_wire[192]), .CP(
        clk), .Q(o_data_bus[192]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(o_data_bus_wire[191]), .CP(
        clk), .Q(o_data_bus[191]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(o_data_bus_wire[190]), .CP(
        clk), .Q(o_data_bus[190]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(o_data_bus_wire[189]), .CP(
        clk), .Q(o_data_bus[189]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(o_data_bus_wire[188]), .CP(
        clk), .Q(o_data_bus[188]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(o_data_bus_wire[187]), .CP(
        clk), .Q(o_data_bus[187]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(o_data_bus_wire[186]), .CP(
        clk), .Q(o_data_bus[186]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(o_data_bus_wire[185]), .CP(
        clk), .Q(o_data_bus[185]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(o_data_bus_wire[184]), .CP(
        clk), .Q(o_data_bus[184]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(o_data_bus_wire[183]), .CP(
        clk), .Q(o_data_bus[183]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(o_data_bus_wire[182]), .CP(
        clk), .Q(o_data_bus[182]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(o_data_bus_wire[181]), .CP(
        clk), .Q(o_data_bus[181]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(o_data_bus_wire[180]), .CP(
        clk), .Q(o_data_bus[180]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(o_data_bus_wire[179]), .CP(
        clk), .Q(o_data_bus[179]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(o_data_bus_wire[177]), .CP(
        clk), .Q(o_data_bus[177]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(o_data_bus_wire[176]), .CP(
        clk), .Q(o_data_bus[176]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(o_data_bus_wire[175]), .CP(
        clk), .Q(o_data_bus[175]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(o_data_bus_wire[174]), .CP(
        clk), .Q(o_data_bus[174]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(o_data_bus_wire[173]), .CP(
        clk), .Q(o_data_bus[173]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(o_data_bus_wire[172]), .CP(
        clk), .Q(o_data_bus[172]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(o_data_bus_wire[171]), .CP(
        clk), .Q(o_data_bus[171]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(o_data_bus_wire[170]), .CP(
        clk), .Q(o_data_bus[170]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(o_data_bus_wire[169]), .CP(
        clk), .Q(o_data_bus[169]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(o_data_bus_wire[168]), .CP(
        clk), .Q(o_data_bus[168]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(o_data_bus_wire[167]), .CP(
        clk), .Q(o_data_bus[167]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(o_data_bus_wire[166]), .CP(
        clk), .Q(o_data_bus[166]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(o_data_bus_wire[165]), .CP(
        clk), .Q(o_data_bus[165]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(o_data_bus_wire[164]), .CP(
        clk), .Q(o_data_bus[164]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(o_data_bus_wire[163]), .CP(
        clk), .Q(o_data_bus[163]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(o_data_bus_wire[162]), .CP(
        clk), .Q(o_data_bus[162]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(o_data_bus_wire[161]), .CP(
        clk), .Q(o_data_bus[161]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(o_data_bus_wire[160]), .CP(
        clk), .Q(o_data_bus[160]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(o_data_bus_wire[159]), .CP(
        clk), .Q(o_data_bus[159]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(o_data_bus_wire[158]), .CP(
        clk), .Q(o_data_bus[158]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(o_data_bus_wire[157]), .CP(
        clk), .Q(o_data_bus[157]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(o_data_bus_wire[156]), .CP(
        clk), .Q(o_data_bus[156]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(o_data_bus_wire[155]), .CP(
        clk), .Q(o_data_bus[155]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(o_data_bus_wire[154]), .CP(
        clk), .Q(o_data_bus[154]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(o_data_bus_wire[153]), .CP(
        clk), .Q(o_data_bus[153]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(o_data_bus_wire[152]), .CP(
        clk), .Q(o_data_bus[152]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(o_data_bus_wire[151]), .CP(
        clk), .Q(o_data_bus[151]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(o_data_bus_wire[150]), .CP(
        clk), .Q(o_data_bus[150]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(o_data_bus_wire[149]), .CP(
        clk), .Q(o_data_bus[149]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(o_data_bus_wire[148]), .CP(
        clk), .Q(o_data_bus[148]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(o_data_bus_wire[147]), .CP(
        clk), .Q(o_data_bus[147]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(o_data_bus_wire[146]), .CP(
        clk), .Q(o_data_bus[146]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(o_data_bus_wire[145]), .CP(
        clk), .Q(o_data_bus[145]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(o_data_bus_wire[144]), .CP(
        clk), .Q(o_data_bus[144]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(o_data_bus_wire[143]), .CP(
        clk), .Q(o_data_bus[143]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(o_data_bus_wire[142]), .CP(
        clk), .Q(o_data_bus[142]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(o_data_bus_wire[141]), .CP(
        clk), .Q(o_data_bus[141]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(o_data_bus_wire[140]), .CP(
        clk), .Q(o_data_bus[140]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(o_data_bus_wire[139]), .CP(
        clk), .Q(o_data_bus[139]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(o_data_bus_wire[138]), .CP(
        clk), .Q(o_data_bus[138]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(o_data_bus_wire[137]), .CP(
        clk), .Q(o_data_bus[137]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(o_data_bus_wire[136]), .CP(
        clk), .Q(o_data_bus[136]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(o_data_bus_wire[135]), .CP(
        clk), .Q(o_data_bus[135]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(o_data_bus_wire[134]), .CP(
        clk), .Q(o_data_bus[134]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(o_data_bus_wire[133]), .CP(
        clk), .Q(o_data_bus[133]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(o_data_bus_wire[132]), .CP(
        clk), .Q(o_data_bus[132]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(o_data_bus_wire[131]), .CP(
        clk), .Q(o_data_bus[131]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(o_data_bus_wire[130]), .CP(
        clk), .Q(o_data_bus[130]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(o_data_bus_wire[129]), .CP(
        clk), .Q(o_data_bus[129]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(o_data_bus_wire[128]), .CP(
        clk), .Q(o_data_bus[128]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(o_data_bus_wire[127]), .CP(
        clk), .Q(o_data_bus[127]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(o_data_bus_wire[126]), .CP(
        clk), .Q(o_data_bus[126]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(o_data_bus_wire[125]), .CP(
        clk), .Q(o_data_bus[125]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(o_data_bus_wire[124]), .CP(
        clk), .Q(o_data_bus[124]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(o_data_bus_wire[123]), .CP(
        clk), .Q(o_data_bus[123]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(o_data_bus_wire[122]), .CP(
        clk), .Q(o_data_bus[122]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(o_data_bus_wire[121]), .CP(
        clk), .Q(o_data_bus[121]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(o_data_bus_wire[120]), .CP(
        clk), .Q(o_data_bus[120]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(o_data_bus_wire[119]), .CP(
        clk), .Q(o_data_bus[119]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(o_data_bus_wire[118]), .CP(
        clk), .Q(o_data_bus[118]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(o_data_bus_wire[117]), .CP(
        clk), .Q(o_data_bus[117]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(o_data_bus_wire[116]), .CP(
        clk), .Q(o_data_bus[116]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(o_data_bus_wire[115]), .CP(
        clk), .Q(o_data_bus[115]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(o_data_bus_wire[114]), .CP(
        clk), .Q(o_data_bus[114]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(o_data_bus_wire[113]), .CP(
        clk), .Q(o_data_bus[113]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(o_data_bus_wire[112]), .CP(
        clk), .Q(o_data_bus[112]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(o_data_bus_wire[110]), .CP(
        clk), .Q(o_data_bus[110]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(o_data_bus_wire[109]), .CP(
        clk), .Q(o_data_bus[109]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(o_data_bus_wire[108]), .CP(
        clk), .Q(o_data_bus[108]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(o_data_bus_wire[107]), .CP(
        clk), .Q(o_data_bus[107]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(o_data_bus_wire[106]), .CP(
        clk), .Q(o_data_bus[106]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(o_data_bus_wire[105]), .CP(
        clk), .Q(o_data_bus[105]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(o_data_bus_wire[104]), .CP(
        clk), .Q(o_data_bus[104]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(o_data_bus_wire[103]), .CP(
        clk), .Q(o_data_bus[103]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(o_data_bus_wire[101]), .CP(
        clk), .Q(o_data_bus[101]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(o_data_bus_wire[100]), .CP(
        clk), .Q(o_data_bus[100]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(o_data_bus_wire[99]), .CP(clk), 
        .Q(o_data_bus[99]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(o_data_bus_wire[98]), .CP(clk), 
        .Q(o_data_bus[98]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(o_data_bus_wire[97]), .CP(clk), 
        .Q(o_data_bus[97]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(o_data_bus_wire[96]), .CP(clk), 
        .Q(o_data_bus[96]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(o_data_bus_wire[95]), .CP(clk), 
        .Q(o_data_bus[95]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(o_data_bus_wire[94]), .CP(clk), 
        .Q(o_data_bus[94]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(o_data_bus_wire[93]), .CP(clk), 
        .Q(o_data_bus[93]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(o_data_bus_wire[92]), .CP(clk), 
        .Q(o_data_bus[92]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(o_data_bus_wire[91]), .CP(clk), 
        .Q(o_data_bus[91]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(o_data_bus_wire[89]), .CP(clk), 
        .Q(o_data_bus[89]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(o_data_bus_wire[88]), .CP(clk), 
        .Q(o_data_bus[88]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(o_data_bus_wire[87]), .CP(clk), 
        .Q(o_data_bus[87]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(o_data_bus_wire[86]), .CP(clk), 
        .Q(o_data_bus[86]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(o_data_bus_wire[85]), .CP(clk), 
        .Q(o_data_bus[85]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(o_data_bus_wire[84]), .CP(clk), 
        .Q(o_data_bus[84]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(o_data_bus_wire[83]), .CP(clk), 
        .Q(o_data_bus[83]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(o_data_bus_wire[82]), .CP(clk), 
        .Q(o_data_bus[82]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(o_data_bus_wire[81]), .CP(clk), 
        .Q(o_data_bus[81]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(o_data_bus_wire[80]), .CP(clk), 
        .Q(o_data_bus[80]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(o_data_bus_wire[79]), .CP(clk), 
        .Q(o_data_bus[79]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(o_data_bus_wire[78]), .CP(clk), 
        .Q(o_data_bus[78]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(o_data_bus_wire[77]), .CP(clk), 
        .Q(o_data_bus[77]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(o_data_bus_wire[76]), .CP(clk), 
        .Q(o_data_bus[76]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(o_data_bus_wire[75]), .CP(clk), 
        .Q(o_data_bus[75]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(o_data_bus_wire[74]), .CP(clk), 
        .Q(o_data_bus[74]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(o_data_bus_wire[73]), .CP(clk), 
        .Q(o_data_bus[73]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(o_data_bus_wire[72]), .CP(clk), 
        .Q(o_data_bus[72]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(o_data_bus_wire[71]), .CP(clk), 
        .Q(o_data_bus[71]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(o_data_bus_wire[70]), .CP(clk), 
        .Q(o_data_bus[70]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(o_data_bus_wire[69]), .CP(clk), 
        .Q(o_data_bus[69]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(o_data_bus_wire[67]), .CP(clk), 
        .Q(o_data_bus[67]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(o_data_bus_wire[66]), .CP(clk), 
        .Q(o_data_bus[66]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(o_data_bus_wire[65]), .CP(clk), 
        .Q(o_data_bus[65]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(o_data_bus_wire[64]), .CP(clk), 
        .Q(o_data_bus[64]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(o_data_bus_wire[63]), .CP(clk), 
        .Q(o_data_bus[63]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(o_data_bus_wire[62]), .CP(clk), 
        .Q(o_data_bus[62]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(o_data_bus_wire[61]), .CP(clk), 
        .Q(o_data_bus[61]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(o_data_bus_wire[60]), .CP(clk), 
        .Q(o_data_bus[60]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(o_data_bus_wire[59]), .CP(clk), 
        .Q(o_data_bus[59]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(o_data_bus_wire[58]), .CP(clk), 
        .Q(o_data_bus[58]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(o_data_bus_wire[57]), .CP(clk), 
        .Q(o_data_bus[57]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(o_data_bus_wire[56]), .CP(clk), 
        .Q(o_data_bus[56]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(o_data_bus_wire[55]), .CP(clk), 
        .Q(o_data_bus[55]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(o_data_bus_wire[54]), .CP(clk), 
        .Q(o_data_bus[54]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(o_data_bus_wire[53]), .CP(clk), 
        .Q(o_data_bus[53]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(o_data_bus_wire[52]), .CP(clk), 
        .Q(o_data_bus[52]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(o_data_bus_wire[51]), .CP(clk), 
        .Q(o_data_bus[51]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(o_data_bus_wire[50]), .CP(clk), 
        .Q(o_data_bus[50]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(o_data_bus_wire[49]), .CP(clk), 
        .Q(o_data_bus[49]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(o_data_bus_wire[48]), .CP(clk), 
        .Q(o_data_bus[48]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(o_data_bus_wire[47]), .CP(clk), 
        .Q(o_data_bus[47]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(o_data_bus_wire[46]), .CP(clk), 
        .Q(o_data_bus[46]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(o_data_bus_wire[45]), .CP(clk), 
        .Q(o_data_bus[45]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(o_data_bus_wire[44]), .CP(clk), 
        .Q(o_data_bus[44]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(o_data_bus_wire[43]), .CP(clk), 
        .Q(o_data_bus[43]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(o_data_bus_wire[42]), .CP(clk), 
        .Q(o_data_bus[42]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(o_data_bus_wire[41]), .CP(clk), 
        .Q(o_data_bus[41]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(o_data_bus_wire[40]), .CP(clk), 
        .Q(o_data_bus[40]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(o_data_bus_wire[39]), .CP(clk), 
        .Q(o_data_bus[39]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(o_data_bus_wire[38]), .CP(clk), 
        .Q(o_data_bus[38]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(o_data_bus_wire[37]), .CP(clk), 
        .Q(o_data_bus[37]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(o_data_bus_wire[36]), .CP(clk), 
        .Q(o_data_bus[36]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(o_data_bus_wire[35]), .CP(clk), 
        .Q(o_data_bus[35]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(o_data_bus_wire[34]), .CP(clk), 
        .Q(o_data_bus[34]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(o_data_bus_wire[33]), .CP(clk), 
        .Q(o_data_bus[33]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(o_data_bus_wire[32]), .CP(clk), 
        .Q(o_data_bus[32]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(o_data_bus_wire[31]), .CP(clk), 
        .Q(o_data_bus[31]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(o_data_bus_wire[30]), .CP(clk), 
        .Q(o_data_bus[30]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(o_data_bus_wire[29]), .CP(clk), 
        .Q(o_data_bus[29]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(o_data_bus_wire[28]), .CP(clk), 
        .Q(o_data_bus[28]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(o_data_bus_wire[27]), .CP(clk), 
        .Q(o_data_bus[27]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(o_data_bus_wire[26]), .CP(clk), 
        .Q(o_data_bus[26]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(o_data_bus_wire[25]), .CP(clk), 
        .Q(o_data_bus[25]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(o_data_bus_wire[24]), .CP(clk), 
        .Q(o_data_bus[24]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(o_data_bus_wire[23]), .CP(clk), 
        .Q(o_data_bus[23]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(o_data_bus_wire[22]), .CP(clk), 
        .Q(o_data_bus[22]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(o_data_bus_wire[21]), .CP(clk), 
        .Q(o_data_bus[21]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(o_data_bus_wire[20]), .CP(clk), 
        .Q(o_data_bus[20]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(o_data_bus_wire[19]), .CP(clk), 
        .Q(o_data_bus[19]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(o_data_bus_wire[18]), .CP(clk), 
        .Q(o_data_bus[18]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(o_data_bus_wire[17]), .CP(clk), 
        .Q(o_data_bus[17]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(o_data_bus_wire[16]), .CP(clk), 
        .Q(o_data_bus[16]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(o_data_bus_wire[15]), .CP(clk), 
        .Q(o_data_bus[15]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(o_data_bus_wire[14]), .CP(clk), 
        .Q(o_data_bus[14]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(o_data_bus_wire[13]), .CP(clk), 
        .Q(o_data_bus[13]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(o_data_bus_wire[12]), .CP(clk), 
        .Q(o_data_bus[12]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(o_data_bus_wire[11]), .CP(clk), 
        .Q(o_data_bus[11]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(o_data_bus_wire[10]), .CP(clk), 
        .Q(o_data_bus[10]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(o_data_bus_wire[9]), .CP(clk), 
        .Q(o_data_bus[9]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(o_data_bus_wire[8]), .CP(clk), 
        .Q(o_data_bus[8]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(o_data_bus_wire[7]), .CP(clk), 
        .Q(o_data_bus[7]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(o_data_bus_wire[6]), .CP(clk), 
        .Q(o_data_bus[6]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(o_data_bus_wire[5]), .CP(clk), 
        .Q(o_data_bus[5]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(o_data_bus_wire[4]), .CP(clk), 
        .Q(o_data_bus[4]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(o_data_bus_wire[3]), .CP(clk), 
        .Q(o_data_bus[3]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(o_data_bus_wire[2]), .CP(clk), 
        .Q(o_data_bus[2]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(o_data_bus_wire[1]), .CP(clk), 
        .Q(o_data_bus[1]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(o_data_bus_wire[0]), .CP(clk), 
        .Q(o_data_bus[0]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_307_ ( .CN(i_data_bus[307]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[307]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_306_ ( .CN(i_data_bus[306]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[306]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_305_ ( .CN(i_data_bus[305]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[305]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_304_ ( .CN(i_data_bus[304]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[304]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_303_ ( .CN(i_data_bus[303]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[303]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_302_ ( .CN(i_data_bus[302]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[302]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_301_ ( .CN(i_data_bus[301]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[301]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_295_ ( .CN(i_data_bus[295]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[295]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_294_ ( .CN(i_data_bus[294]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[294]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_293_ ( .CN(i_data_bus[293]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[293]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_292_ ( .CN(i_data_bus[292]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[292]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_283_ ( .CN(i_data_bus[283]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[283]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_282_ ( .CN(i_data_bus[282]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[282]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_281_ ( .CN(i_data_bus[281]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[281]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_280_ ( .CN(i_data_bus[280]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[280]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_279_ ( .CN(i_data_bus[279]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[279]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_278_ ( .CN(i_data_bus[278]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[278]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_277_ ( .CN(i_data_bus[277]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[277]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_276_ ( .CN(i_data_bus[276]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[276]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_275_ ( .CN(i_data_bus[275]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[275]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_274_ ( .CN(i_data_bus[274]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[274]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_273_ ( .CN(i_data_bus[273]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[273]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_272_ ( .CN(i_data_bus[272]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[272]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_271_ ( .CN(i_data_bus[271]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[271]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_270_ ( .CN(i_data_bus[270]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[270]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_269_ ( .CN(i_data_bus[269]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[269]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_268_ ( .CN(i_data_bus[268]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[268]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_267_ ( .CN(i_data_bus[267]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[267]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_266_ ( .CN(i_data_bus[266]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[266]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_265_ ( .CN(i_data_bus[265]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[265]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_264_ ( .CN(i_data_bus[264]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[264]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_263_ ( .CN(i_data_bus[263]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[263]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_262_ ( .CN(i_data_bus[262]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[262]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_261_ ( .CN(i_data_bus[261]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[261]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_260_ ( .CN(i_data_bus[260]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[260]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_259_ ( .CN(i_data_bus[259]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[259]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_258_ ( .CN(i_data_bus[258]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[258]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_257_ ( .CN(i_data_bus[257]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[257]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_256_ ( .CN(i_data_bus[256]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[256]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_255_ ( .CN(i_data_bus[255]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[255]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_254_ ( .CN(i_data_bus[254]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[254]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_253_ ( .CN(i_data_bus[253]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[253]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_252_ ( .CN(i_data_bus[252]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[252]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_251_ ( .CN(i_data_bus[251]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[251]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_250_ ( .CN(i_data_bus[250]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[250]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_249_ ( .CN(i_data_bus[249]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[249]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_248_ ( .CN(i_data_bus[248]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[248]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_247_ ( .CN(i_data_bus[247]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[247]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_246_ ( .CN(i_data_bus[246]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[246]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_245_ ( .CN(i_data_bus[245]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[245]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_244_ ( .CN(i_data_bus[244]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[244]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_243_ ( .CN(i_data_bus[243]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[243]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_242_ ( .CN(i_data_bus[242]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[242]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_241_ ( .CN(i_data_bus[241]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[241]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_240_ ( .CN(i_data_bus[240]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[240]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_239_ ( .CN(i_data_bus[239]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[239]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_238_ ( .CN(i_data_bus[238]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[238]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_237_ ( .CN(i_data_bus[237]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[237]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_236_ ( .CN(i_data_bus[236]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[236]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_235_ ( .CN(i_data_bus[235]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[235]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_234_ ( .CN(i_data_bus[234]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[234]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_233_ ( .CN(i_data_bus[233]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[233]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_232_ ( .CN(i_data_bus[232]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[232]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_231_ ( .CN(i_data_bus[231]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[231]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_230_ ( .CN(i_data_bus[230]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[230]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_229_ ( .CN(i_data_bus[229]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[229]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_223_ ( .CN(i_data_bus[223]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[223]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_222_ ( .CN(i_data_bus[222]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[222]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_221_ ( .CN(i_data_bus[221]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[221]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_220_ ( .CN(i_data_bus[220]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[220]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_211_ ( .CN(i_data_bus[211]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[211]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_210_ ( .CN(i_data_bus[210]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[210]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_209_ ( .CN(i_data_bus[209]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[209]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_208_ ( .CN(i_data_bus[208]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[208]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_207_ ( .CN(i_data_bus[207]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[207]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_206_ ( .CN(i_data_bus[206]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[206]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_205_ ( .CN(i_data_bus[205]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[205]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_204_ ( .CN(i_data_bus[204]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[204]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_203_ ( .CN(i_data_bus[203]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[203]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_202_ ( .CN(i_data_bus[202]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[202]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_201_ ( .CN(i_data_bus[201]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[201]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_200_ ( .CN(i_data_bus[200]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[200]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_199_ ( .CN(i_data_bus[199]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[199]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_198_ ( .CN(i_data_bus[198]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[198]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_197_ ( .CN(i_data_bus[197]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[197]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_196_ ( .CN(i_data_bus[196]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[196]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_195_ ( .CN(i_data_bus[195]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[195]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_194_ ( .CN(i_data_bus[194]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[194]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_193_ ( .CN(i_data_bus[193]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[193]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_192_ ( .CN(i_data_bus[192]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[192]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_191_ ( .CN(i_data_bus[191]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[191]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_190_ ( .CN(i_data_bus[190]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[190]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_189_ ( .CN(i_data_bus[189]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[189]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_188_ ( .CN(i_data_bus[188]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[188]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_187_ ( .CN(i_data_bus[187]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[187]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_186_ ( .CN(i_data_bus[186]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[186]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_185_ ( .CN(i_data_bus[185]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[185]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_184_ ( .CN(i_data_bus[184]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[184]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_183_ ( .CN(i_data_bus[183]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[183]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_182_ ( .CN(i_data_bus[182]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[182]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_181_ ( .CN(i_data_bus[181]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[181]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_180_ ( .CN(i_data_bus[180]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[180]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_179_ ( .CN(i_data_bus[179]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[179]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_178_ ( .CN(i_data_bus[178]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[178]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_177_ ( .CN(i_data_bus[177]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[177]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_176_ ( .CN(i_data_bus[176]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[176]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_175_ ( .CN(i_data_bus[175]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[175]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_174_ ( .CN(i_data_bus[174]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[174]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_173_ ( .CN(i_data_bus[173]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[173]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_172_ ( .CN(i_data_bus[172]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[172]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_171_ ( .CN(i_data_bus[171]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[171]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_170_ ( .CN(i_data_bus[170]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[170]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_169_ ( .CN(i_data_bus[169]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[169]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_168_ ( .CN(i_data_bus[168]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[168]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_167_ ( .CN(i_data_bus[167]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[167]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_166_ ( .CN(i_data_bus[166]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[166]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_165_ ( .CN(i_data_bus[165]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[165]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_164_ ( .CN(i_data_bus[164]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[164]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_163_ ( .CN(i_data_bus[163]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[163]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_162_ ( .CN(i_data_bus[162]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[162]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_161_ ( .CN(i_data_bus[161]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[161]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_160_ ( .CN(i_data_bus[160]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[160]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_159_ ( .CN(i_data_bus[159]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[159]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_158_ ( .CN(i_data_bus[158]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[158]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_157_ ( .CN(i_data_bus[157]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[157]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_151_ ( .CN(i_data_bus[151]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[151]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_150_ ( .CN(i_data_bus[150]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[150]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_149_ ( .CN(i_data_bus[149]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[149]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_148_ ( .CN(i_data_bus[148]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[148]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_139_ ( .CN(i_data_bus[139]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[139]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_138_ ( .CN(i_data_bus[138]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[138]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_137_ ( .CN(i_data_bus[137]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[137]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_136_ ( .CN(i_data_bus[136]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[136]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_135_ ( .CN(i_data_bus[135]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[135]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_134_ ( .CN(i_data_bus[134]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[134]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_133_ ( .CN(i_data_bus[133]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[133]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_132_ ( .CN(i_data_bus[132]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[132]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_131_ ( .CN(i_data_bus[131]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[131]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_130_ ( .CN(i_data_bus[130]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[130]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_129_ ( .CN(i_data_bus[129]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[129]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_128_ ( .CN(i_data_bus[128]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[128]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_115_ ( .CN(i_data_bus[115]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[115]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_114_ ( .CN(i_data_bus[114]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[114]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_113_ ( .CN(i_data_bus[113]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[113]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_112_ ( .CN(i_data_bus[112]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[112]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_111_ ( .CN(i_data_bus[111]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[111]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_91_ ( .CN(i_data_bus[91]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[91]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_90_ ( .CN(i_data_bus[90]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[90]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_89_ ( .CN(i_data_bus[89]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[89]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_88_ ( .CN(i_data_bus[88]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[88]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_87_ ( .CN(i_data_bus[87]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[87]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_86_ ( .CN(i_data_bus[86]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[86]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_85_ ( .CN(i_data_bus[85]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[85]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_79_ ( .CN(i_data_bus[79]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[79]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_78_ ( .CN(i_data_bus[78]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[78]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_77_ ( .CN(i_data_bus[77]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[77]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_76_ ( .CN(i_data_bus[76]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[76]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_67_ ( .CN(i_data_bus[67]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[67]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_66_ ( .CN(i_data_bus[66]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[66]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_65_ ( .CN(i_data_bus[65]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[65]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_64_ ( .CN(i_data_bus[64]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[64]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_63_ ( .CN(i_data_bus[63]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[63]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_62_ ( .CN(i_data_bus[62]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[62]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_61_ ( .CN(i_data_bus[61]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[61]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_60_ ( .CN(i_data_bus[60]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[60]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_59_ ( .CN(i_data_bus[59]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[59]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_58_ ( .CN(i_data_bus[58]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[58]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_57_ ( .CN(i_data_bus[57]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[57]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_56_ ( .CN(i_data_bus[56]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[56]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_55_ ( .CN(i_data_bus[55]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[55]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_54_ ( .CN(i_data_bus[54]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[54]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_53_ ( .CN(i_data_bus[53]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[53]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_52_ ( .CN(i_data_bus[52]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[52]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_51_ ( .CN(i_data_bus[51]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[51]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_50_ ( .CN(i_data_bus[50]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[50]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_49_ ( .CN(i_data_bus[49]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[49]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_48_ ( .CN(i_data_bus[48]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[48]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_47_ ( .CN(i_data_bus[47]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[47]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_46_ ( .CN(i_data_bus[46]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[46]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_45_ ( .CN(i_data_bus[45]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[45]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_44_ ( .CN(i_data_bus[44]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[44]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_43_ ( .CN(i_data_bus[43]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[43]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_42_ ( .CN(i_data_bus[42]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[42]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_41_ ( .CN(i_data_bus[41]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[41]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_40_ ( .CN(i_data_bus[40]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[40]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_39_ ( .CN(i_data_bus[39]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[39]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_38_ ( .CN(i_data_bus[38]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[38]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_37_ ( .CN(i_data_bus[37]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[37]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_36_ ( .CN(i_data_bus[36]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[36]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_35_ ( .CN(i_data_bus[35]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[35]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_34_ ( .CN(i_data_bus[34]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[34]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_33_ ( .CN(i_data_bus[33]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[33]) );
  DFKCNQD1BWP30P140LVT i_data_bus_reg_reg_25_ ( .CN(i_data_bus[25]), .D(n15), 
        .CP(clk), .Q(i_data_bus_reg[25]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_139_ ( .D(N1198), .CP(clk), .Q(
        i_cmd_reg[139]) );
  DFQD1BWP30P140LVT i_cmd_reg_reg_221_ ( .D(N1280), .CP(clk), .Q(
        i_cmd_reg[221]) );
  DFQD2BWP30P140LVT i_cmd_reg_reg_147_ ( .D(N1206), .CP(clk), .Q(
        i_cmd_reg[147]) );
  DFD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(o_data_bus_wire[68]), .CP(clk), 
        .Q(o_data_bus[68]) );
  DFD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(o_data_bus_wire[178]), .CP(clk), .Q(o_data_bus[178]) );
  DFD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(o_data_bus_wire[90]), .CP(clk), 
        .Q(o_data_bus[90]) );
  DFD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(o_data_bus_wire[111]), .CP(clk), .Q(o_data_bus[111]) );
  DFD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(o_data_bus_wire[102]), .CP(clk), .Q(o_data_bus[102]) );
  BUFFD4BWP30P140LVT U1316 ( .I(n15), .Z(n14) );
  CKBD1BWP30P140LVT U1317 ( .I(n15), .Z(n12) );
  INR2D6BWP30P140LVT U1318 ( .A1(i_en), .B1(rst), .ZN(n15) );
  CKAN2D1BWP30P140LVT U1319 ( .A1(n15), .A2(i_data_bus[4]), .Z(N39) );
  CKAN2D1BWP30P140LVT U1320 ( .A1(n15), .A2(i_data_bus[5]), .Z(N40) );
  CKAN2D1BWP30P140LVT U1321 ( .A1(n15), .A2(i_data_bus[6]), .Z(N41) );
  CKAN2D1BWP30P140LVT U1322 ( .A1(n15), .A2(i_data_bus[7]), .Z(N42) );
  CKAN2D1BWP30P140LVT U1323 ( .A1(n15), .A2(i_data_bus[13]), .Z(N48) );
  CKAN2D1BWP30P140LVT U1324 ( .A1(n15), .A2(i_data_bus[14]), .Z(N49) );
  CKAN2D1BWP30P140LVT U1325 ( .A1(n15), .A2(i_data_bus[15]), .Z(N50) );
  CKAN2D1BWP30P140LVT U1326 ( .A1(n15), .A2(i_data_bus[16]), .Z(N51) );
  CKAN2D1BWP30P140LVT U1327 ( .A1(n15), .A2(i_data_bus[17]), .Z(N52) );
  CKAN2D1BWP30P140LVT U1328 ( .A1(n15), .A2(i_data_bus[18]), .Z(N53) );
  CKAN2D1BWP30P140LVT U1329 ( .A1(n15), .A2(i_data_bus[19]), .Z(N54) );
  CKAN2D1BWP30P140LVT U1330 ( .A1(n14), .A2(i_data_bus[321]), .Z(N356) );
  CKAN2D1BWP30P140LVT U1331 ( .A1(n14), .A2(i_data_bus[322]), .Z(N357) );
  CKAN2D1BWP30P140LVT U1332 ( .A1(n14), .A2(i_data_bus[323]), .Z(N358) );
  CKAN2D1BWP30P140LVT U1333 ( .A1(n14), .A2(i_data_bus[324]), .Z(N359) );
  CKAN2D1BWP30P140LVT U1334 ( .A1(n14), .A2(i_data_bus[325]), .Z(N360) );
  CKAN2D1BWP30P140LVT U1335 ( .A1(n14), .A2(i_data_bus[326]), .Z(N361) );
  CKAN2D1BWP30P140LVT U1336 ( .A1(n14), .A2(i_data_bus[327]), .Z(N362) );
  CKAN2D1BWP30P140LVT U1337 ( .A1(n14), .A2(i_data_bus[328]), .Z(N363) );
  CKAN2D1BWP30P140LVT U1338 ( .A1(n14), .A2(i_data_bus[329]), .Z(N364) );
  CKAN2D1BWP30P140LVT U1339 ( .A1(n14), .A2(i_data_bus[330]), .Z(N365) );
  CKAN2D1BWP30P140LVT U1340 ( .A1(n14), .A2(i_data_bus[331]), .Z(N366) );
  CKAN2D1BWP30P140LVT U1341 ( .A1(n14), .A2(i_data_bus[332]), .Z(N367) );
  CKAN2D1BWP30P140LVT U1342 ( .A1(n14), .A2(i_data_bus[333]), .Z(N368) );
  CKAN2D1BWP30P140LVT U1343 ( .A1(n14), .A2(i_data_bus[334]), .Z(N369) );
  CKAN2D1BWP30P140LVT U1344 ( .A1(n14), .A2(i_data_bus[335]), .Z(N370) );
  CKAN2D1BWP30P140LVT U1345 ( .A1(n14), .A2(i_data_bus[336]), .Z(N371) );
  CKAN2D1BWP30P140LVT U1346 ( .A1(n14), .A2(i_data_bus[337]), .Z(N372) );
  CKAN2D1BWP30P140LVT U1347 ( .A1(n14), .A2(i_data_bus[338]), .Z(N373) );
  CKAN2D1BWP30P140LVT U1348 ( .A1(n14), .A2(i_data_bus[339]), .Z(N374) );
  CKAN2D1BWP30P140LVT U1349 ( .A1(n14), .A2(i_data_bus[340]), .Z(N375) );
  CKAN2D1BWP30P140LVT U1350 ( .A1(n14), .A2(i_data_bus[341]), .Z(N376) );
  CKAN2D1BWP30P140LVT U1351 ( .A1(n14), .A2(i_data_bus[342]), .Z(N377) );
  CKAN2D1BWP30P140LVT U1352 ( .A1(n14), .A2(i_data_bus[343]), .Z(N378) );
  CKAN2D1BWP30P140LVT U1353 ( .A1(n14), .A2(i_data_bus[344]), .Z(N379) );
  CKAN2D1BWP30P140LVT U1354 ( .A1(n14), .A2(i_data_bus[345]), .Z(N380) );
  CKAN2D1BWP30P140LVT U1355 ( .A1(n14), .A2(i_data_bus[346]), .Z(N381) );
  CKAN2D1BWP30P140LVT U1356 ( .A1(n14), .A2(i_data_bus[347]), .Z(N382) );
  CKAN2D1BWP30P140LVT U1357 ( .A1(n14), .A2(i_data_bus[348]), .Z(N383) );
  CKAN2D1BWP30P140LVT U1358 ( .A1(n14), .A2(i_data_bus[349]), .Z(N384) );
  CKAN2D1BWP30P140LVT U1359 ( .A1(n14), .A2(i_data_bus[350]), .Z(N385) );
  CKAN2D1BWP30P140LVT U1360 ( .A1(n14), .A2(i_data_bus[351]), .Z(N386) );
  CKAN2D1BWP30P140LVT U1361 ( .A1(n14), .A2(i_data_bus[352]), .Z(N387) );
  CKAN2D1BWP30P140LVT U1362 ( .A1(n14), .A2(i_data_bus[353]), .Z(N388) );
  CKAN2D1BWP30P140LVT U1363 ( .A1(n14), .A2(i_data_bus[354]), .Z(N389) );
  CKAN2D1BWP30P140LVT U1364 ( .A1(n14), .A2(i_data_bus[355]), .Z(N390) );
  CKAN2D1BWP30P140LVT U1365 ( .A1(n14), .A2(i_data_bus[364]), .Z(N399) );
  CKAN2D1BWP30P140LVT U1366 ( .A1(n14), .A2(i_data_bus[365]), .Z(N400) );
  CKAN2D1BWP30P140LVT U1367 ( .A1(n14), .A2(i_data_bus[366]), .Z(N401) );
  CKAN2D1BWP30P140LVT U1368 ( .A1(n14), .A2(i_data_bus[367]), .Z(N402) );
  CKAN2D1BWP30P140LVT U1369 ( .A1(n14), .A2(i_data_bus[373]), .Z(N408) );
  CKAN2D1BWP30P140LVT U1370 ( .A1(n14), .A2(i_data_bus[374]), .Z(N409) );
  CKAN2D1BWP30P140LVT U1371 ( .A1(n14), .A2(i_data_bus[375]), .Z(N410) );
  CKAN2D1BWP30P140LVT U1372 ( .A1(n14), .A2(i_data_bus[376]), .Z(N411) );
  CKAN2D1BWP30P140LVT U1373 ( .A1(n14), .A2(i_data_bus[377]), .Z(N412) );
  CKAN2D1BWP30P140LVT U1374 ( .A1(n14), .A2(i_data_bus[378]), .Z(N413) );
  CKAN2D1BWP30P140LVT U1375 ( .A1(n14), .A2(i_data_bus[379]), .Z(N414) );
  CKAN2D1BWP30P140LVT U1376 ( .A1(n14), .A2(i_data_bus[393]), .Z(N428) );
  CKAN2D1BWP30P140LVT U1377 ( .A1(n14), .A2(i_data_bus[394]), .Z(N429) );
  CKAN2D1BWP30P140LVT U1378 ( .A1(n14), .A2(i_data_bus[395]), .Z(N430) );
  CKAN2D1BWP30P140LVT U1379 ( .A1(n14), .A2(i_data_bus[396]), .Z(N431) );
  CKAN2D1BWP30P140LVT U1380 ( .A1(n14), .A2(i_data_bus[397]), .Z(N432) );
  CKAN2D1BWP30P140LVT U1381 ( .A1(n14), .A2(i_data_bus[398]), .Z(N433) );
  CKAN2D1BWP30P140LVT U1382 ( .A1(n14), .A2(i_data_bus[399]), .Z(N434) );
  CKAN2D1BWP30P140LVT U1383 ( .A1(n14), .A2(i_data_bus[400]), .Z(N435) );
  CKAN2D1BWP30P140LVT U1384 ( .A1(n14), .A2(i_data_bus[401]), .Z(N436) );
  CKAN2D1BWP30P140LVT U1385 ( .A1(n14), .A2(i_data_bus[402]), .Z(N437) );
  CKAN2D1BWP30P140LVT U1386 ( .A1(n14), .A2(i_data_bus[403]), .Z(N438) );
  CKAN2D1BWP30P140LVT U1387 ( .A1(n14), .A2(i_data_bus[404]), .Z(N439) );
  CKAN2D1BWP30P140LVT U1388 ( .A1(n14), .A2(i_data_bus[405]), .Z(N440) );
  CKAN2D1BWP30P140LVT U1389 ( .A1(n14), .A2(i_data_bus[406]), .Z(N441) );
  CKAN2D1BWP30P140LVT U1390 ( .A1(n14), .A2(i_data_bus[407]), .Z(N442) );
  CKAN2D1BWP30P140LVT U1391 ( .A1(n14), .A2(i_data_bus[408]), .Z(N443) );
  CKAN2D1BWP30P140LVT U1392 ( .A1(n14), .A2(i_data_bus[409]), .Z(N444) );
  CKAN2D1BWP30P140LVT U1393 ( .A1(n14), .A2(i_data_bus[410]), .Z(N445) );
  CKAN2D1BWP30P140LVT U1394 ( .A1(n14), .A2(i_data_bus[411]), .Z(N446) );
  CKAN2D1BWP30P140LVT U1395 ( .A1(n14), .A2(i_data_bus[412]), .Z(N447) );
  CKAN2D1BWP30P140LVT U1396 ( .A1(n14), .A2(i_data_bus[413]), .Z(N448) );
  CKAN2D1BWP30P140LVT U1397 ( .A1(n14), .A2(i_data_bus[414]), .Z(N449) );
  CKAN2D1BWP30P140LVT U1398 ( .A1(n14), .A2(i_data_bus[415]), .Z(N450) );
  CKAN2D1BWP30P140LVT U1399 ( .A1(n14), .A2(i_data_bus[416]), .Z(N451) );
  CKAN2D1BWP30P140LVT U1400 ( .A1(n14), .A2(i_data_bus[417]), .Z(N452) );
  CKAN2D1BWP30P140LVT U1401 ( .A1(n14), .A2(i_data_bus[418]), .Z(N453) );
  CKAN2D1BWP30P140LVT U1402 ( .A1(n14), .A2(i_data_bus[419]), .Z(N454) );
  CKAN2D1BWP30P140LVT U1403 ( .A1(n14), .A2(i_data_bus[420]), .Z(N455) );
  CKAN2D1BWP30P140LVT U1404 ( .A1(n14), .A2(i_data_bus[421]), .Z(N456) );
  CKAN2D1BWP30P140LVT U1405 ( .A1(n14), .A2(i_data_bus[422]), .Z(N457) );
  CKAN2D1BWP30P140LVT U1406 ( .A1(n14), .A2(i_data_bus[423]), .Z(N458) );
  CKAN2D1BWP30P140LVT U1407 ( .A1(n14), .A2(i_data_bus[424]), .Z(N459) );
  CKAN2D1BWP30P140LVT U1408 ( .A1(n14), .A2(i_data_bus[425]), .Z(N460) );
  CKAN2D1BWP30P140LVT U1409 ( .A1(n14), .A2(i_data_bus[426]), .Z(N461) );
  CKAN2D1BWP30P140LVT U1410 ( .A1(n14), .A2(i_data_bus[427]), .Z(N462) );
  CKAN2D1BWP30P140LVT U1411 ( .A1(n14), .A2(i_data_bus[436]), .Z(N471) );
  CKAN2D1BWP30P140LVT U1412 ( .A1(n14), .A2(i_data_bus[437]), .Z(N472) );
  CKAN2D1BWP30P140LVT U1413 ( .A1(n14), .A2(i_data_bus[438]), .Z(N473) );
  CKAN2D1BWP30P140LVT U1414 ( .A1(n14), .A2(i_data_bus[439]), .Z(N474) );
  CKAN2D1BWP30P140LVT U1415 ( .A1(n14), .A2(i_data_bus[445]), .Z(N480) );
  CKAN2D1BWP30P140LVT U1416 ( .A1(n14), .A2(i_data_bus[446]), .Z(N481) );
  CKAN2D1BWP30P140LVT U1417 ( .A1(n14), .A2(i_data_bus[447]), .Z(N482) );
  CKAN2D1BWP30P140LVT U1418 ( .A1(n14), .A2(i_data_bus[448]), .Z(N483) );
  CKAN2D1BWP30P140LVT U1419 ( .A1(n14), .A2(i_data_bus[449]), .Z(N484) );
  CKAN2D1BWP30P140LVT U1420 ( .A1(n14), .A2(i_data_bus[450]), .Z(N485) );
  CKAN2D1BWP30P140LVT U1421 ( .A1(n14), .A2(i_data_bus[451]), .Z(N486) );
  CKAN2D1BWP30P140LVT U1422 ( .A1(n14), .A2(i_data_bus[457]), .Z(N492) );
  CKAN2D1BWP30P140LVT U1423 ( .A1(n14), .A2(i_data_bus[465]), .Z(N500) );
  CKAN2D1BWP30P140LVT U1424 ( .A1(n14), .A2(i_data_bus[466]), .Z(N501) );
  CKAN2D1BWP30P140LVT U1425 ( .A1(n14), .A2(i_data_bus[467]), .Z(N502) );
  CKAN2D1BWP30P140LVT U1426 ( .A1(n14), .A2(i_data_bus[468]), .Z(N503) );
  CKAN2D1BWP30P140LVT U1427 ( .A1(n14), .A2(i_data_bus[469]), .Z(N504) );
  CKAN2D1BWP30P140LVT U1428 ( .A1(n14), .A2(i_data_bus[470]), .Z(N505) );
  CKAN2D1BWP30P140LVT U1429 ( .A1(n14), .A2(i_data_bus[471]), .Z(N506) );
  CKAN2D1BWP30P140LVT U1430 ( .A1(n14), .A2(i_data_bus[472]), .Z(N507) );
  CKAN2D1BWP30P140LVT U1431 ( .A1(n14), .A2(i_data_bus[473]), .Z(N508) );
  CKAN2D1BWP30P140LVT U1432 ( .A1(n14), .A2(i_data_bus[474]), .Z(N509) );
  CKAN2D1BWP30P140LVT U1433 ( .A1(n14), .A2(i_data_bus[475]), .Z(N510) );
  CKAN2D1BWP30P140LVT U1434 ( .A1(n14), .A2(i_data_bus[476]), .Z(N511) );
  CKAN2D1BWP30P140LVT U1435 ( .A1(n14), .A2(i_data_bus[477]), .Z(N512) );
  CKAN2D1BWP30P140LVT U1436 ( .A1(n14), .A2(i_data_bus[478]), .Z(N513) );
  CKAN2D1BWP30P140LVT U1437 ( .A1(n14), .A2(i_data_bus[479]), .Z(N514) );
  CKAN2D1BWP30P140LVT U1438 ( .A1(n14), .A2(i_data_bus[480]), .Z(N515) );
  CKAN2D1BWP30P140LVT U1439 ( .A1(n14), .A2(i_data_bus[481]), .Z(N516) );
  CKAN2D1BWP30P140LVT U1440 ( .A1(n14), .A2(i_data_bus[482]), .Z(N517) );
  CKAN2D1BWP30P140LVT U1441 ( .A1(n14), .A2(i_data_bus[483]), .Z(N518) );
  CKAN2D1BWP30P140LVT U1442 ( .A1(n14), .A2(i_data_bus[484]), .Z(N519) );
  CKAN2D1BWP30P140LVT U1443 ( .A1(n14), .A2(i_data_bus[485]), .Z(N520) );
  CKAN2D1BWP30P140LVT U1444 ( .A1(n14), .A2(i_data_bus[486]), .Z(N521) );
  CKAN2D1BWP30P140LVT U1445 ( .A1(n14), .A2(i_data_bus[487]), .Z(N522) );
  CKAN2D1BWP30P140LVT U1446 ( .A1(n14), .A2(i_data_bus[488]), .Z(N523) );
  CKAN2D1BWP30P140LVT U1447 ( .A1(n14), .A2(i_data_bus[489]), .Z(N524) );
  CKAN2D1BWP30P140LVT U1448 ( .A1(n14), .A2(i_data_bus[490]), .Z(N525) );
  CKAN2D1BWP30P140LVT U1449 ( .A1(n14), .A2(i_data_bus[491]), .Z(N526) );
  CKAN2D1BWP30P140LVT U1450 ( .A1(n14), .A2(i_data_bus[492]), .Z(N527) );
  CKAN2D1BWP30P140LVT U1451 ( .A1(n14), .A2(i_data_bus[493]), .Z(N528) );
  CKAN2D1BWP30P140LVT U1452 ( .A1(n14), .A2(i_data_bus[494]), .Z(N529) );
  CKAN2D1BWP30P140LVT U1453 ( .A1(n14), .A2(i_data_bus[495]), .Z(N530) );
  CKAN2D1BWP30P140LVT U1454 ( .A1(n14), .A2(i_data_bus[496]), .Z(N531) );
  CKAN2D1BWP30P140LVT U1455 ( .A1(n14), .A2(i_data_bus[497]), .Z(N532) );
  CKAN2D1BWP30P140LVT U1456 ( .A1(n14), .A2(i_data_bus[498]), .Z(N533) );
  CKAN2D1BWP30P140LVT U1457 ( .A1(n14), .A2(i_data_bus[499]), .Z(N534) );
  CKAN2D1BWP30P140LVT U1458 ( .A1(n14), .A2(i_data_bus[508]), .Z(N543) );
  CKAN2D1BWP30P140LVT U1459 ( .A1(n14), .A2(i_data_bus[509]), .Z(N544) );
  CKAN2D1BWP30P140LVT U1460 ( .A1(n14), .A2(i_data_bus[510]), .Z(N545) );
  CKAN2D1BWP30P140LVT U1461 ( .A1(n14), .A2(i_data_bus[511]), .Z(N546) );
  CKAN2D1BWP30P140LVT U1462 ( .A1(n14), .A2(i_data_bus[517]), .Z(N552) );
  CKAN2D1BWP30P140LVT U1463 ( .A1(n14), .A2(i_data_bus[518]), .Z(N553) );
  CKAN2D1BWP30P140LVT U1464 ( .A1(n14), .A2(i_data_bus[519]), .Z(N554) );
  CKAN2D1BWP30P140LVT U1465 ( .A1(n14), .A2(i_data_bus[520]), .Z(N555) );
  CKAN2D1BWP30P140LVT U1466 ( .A1(n14), .A2(i_data_bus[521]), .Z(N556) );
  CKAN2D1BWP30P140LVT U1467 ( .A1(n14), .A2(i_data_bus[522]), .Z(N557) );
  CKAN2D1BWP30P140LVT U1468 ( .A1(n14), .A2(i_data_bus[523]), .Z(N558) );
  CKAN2D1BWP30P140LVT U1469 ( .A1(n14), .A2(i_data_bus[543]), .Z(N578) );
  CKAN2D1BWP30P140LVT U1470 ( .A1(n14), .A2(i_data_bus[544]), .Z(N579) );
  CKAN2D1BWP30P140LVT U1471 ( .A1(n14), .A2(i_data_bus[545]), .Z(N580) );
  CKAN2D1BWP30P140LVT U1472 ( .A1(n14), .A2(i_data_bus[546]), .Z(N581) );
  CKAN2D1BWP30P140LVT U1473 ( .A1(n14), .A2(i_data_bus[547]), .Z(N582) );
  CKAN2D1BWP30P140LVT U1474 ( .A1(n14), .A2(i_data_bus[560]), .Z(N595) );
  CKAN2D1BWP30P140LVT U1475 ( .A1(n14), .A2(i_data_bus[561]), .Z(N596) );
  CKAN2D1BWP30P140LVT U1476 ( .A1(n14), .A2(i_data_bus[562]), .Z(N597) );
  CKAN2D1BWP30P140LVT U1477 ( .A1(n14), .A2(i_data_bus[563]), .Z(N598) );
  CKAN2D1BWP30P140LVT U1478 ( .A1(n14), .A2(i_data_bus[564]), .Z(N599) );
  CKAN2D1BWP30P140LVT U1479 ( .A1(n14), .A2(i_data_bus[565]), .Z(N600) );
  CKAN2D1BWP30P140LVT U1480 ( .A1(n14), .A2(i_data_bus[566]), .Z(N601) );
  CKAN2D1BWP30P140LVT U1481 ( .A1(n14), .A2(i_data_bus[567]), .Z(N602) );
  CKAN2D1BWP30P140LVT U1482 ( .A1(n14), .A2(i_data_bus[568]), .Z(N603) );
  CKAN2D1BWP30P140LVT U1483 ( .A1(n14), .A2(i_data_bus[569]), .Z(N604) );
  CKAN2D1BWP30P140LVT U1484 ( .A1(n14), .A2(i_data_bus[570]), .Z(N605) );
  CKAN2D1BWP30P140LVT U1485 ( .A1(n14), .A2(i_data_bus[571]), .Z(N606) );
  CKAN2D1BWP30P140LVT U1486 ( .A1(n14), .A2(i_data_bus[580]), .Z(N615) );
  CKAN2D1BWP30P140LVT U1487 ( .A1(n14), .A2(i_data_bus[581]), .Z(N616) );
  CKAN2D1BWP30P140LVT U1488 ( .A1(n14), .A2(i_data_bus[582]), .Z(N617) );
  CKAN2D1BWP30P140LVT U1489 ( .A1(n14), .A2(i_data_bus[583]), .Z(N618) );
  CKAN2D1BWP30P140LVT U1490 ( .A1(n14), .A2(i_data_bus[589]), .Z(N624) );
  CKAN2D1BWP30P140LVT U1491 ( .A1(n14), .A2(i_data_bus[590]), .Z(N625) );
  CKAN2D1BWP30P140LVT U1492 ( .A1(n14), .A2(i_data_bus[591]), .Z(N626) );
  CKAN2D1BWP30P140LVT U1493 ( .A1(n14), .A2(i_data_bus[592]), .Z(N627) );
  CKAN2D1BWP30P140LVT U1494 ( .A1(n14), .A2(i_data_bus[593]), .Z(N628) );
  CKAN2D1BWP30P140LVT U1495 ( .A1(n14), .A2(i_data_bus[594]), .Z(N629) );
  CKAN2D1BWP30P140LVT U1496 ( .A1(n14), .A2(i_data_bus[595]), .Z(N630) );
  CKAN2D1BWP30P140LVT U1497 ( .A1(n14), .A2(i_data_bus[596]), .Z(N631) );
  CKAN2D1BWP30P140LVT U1498 ( .A1(n14), .A2(i_data_bus[597]), .Z(N632) );
  CKAN2D1BWP30P140LVT U1499 ( .A1(n14), .A2(i_data_bus[598]), .Z(N633) );
  CKAN2D1BWP30P140LVT U1500 ( .A1(n14), .A2(i_data_bus[599]), .Z(N634) );
  CKAN2D1BWP30P140LVT U1501 ( .A1(n14), .A2(i_data_bus[600]), .Z(N635) );
  CKAN2D1BWP30P140LVT U1502 ( .A1(n14), .A2(i_data_bus[601]), .Z(N636) );
  CKAN2D1BWP30P140LVT U1503 ( .A1(n14), .A2(i_data_bus[608]), .Z(N643) );
  CKAN2D1BWP30P140LVT U1504 ( .A1(n14), .A2(i_data_bus[609]), .Z(N644) );
  CKAN2D1BWP30P140LVT U1505 ( .A1(n14), .A2(i_data_bus[610]), .Z(N645) );
  CKAN2D1BWP30P140LVT U1506 ( .A1(n14), .A2(i_data_bus[611]), .Z(N646) );
  CKAN2D1BWP30P140LVT U1507 ( .A1(n14), .A2(i_data_bus[612]), .Z(N647) );
  CKAN2D1BWP30P140LVT U1508 ( .A1(n14), .A2(i_data_bus[613]), .Z(N648) );
  CKAN2D1BWP30P140LVT U1509 ( .A1(n14), .A2(i_data_bus[614]), .Z(N649) );
  CKAN2D1BWP30P140LVT U1510 ( .A1(n14), .A2(i_data_bus[615]), .Z(N650) );
  CKAN2D1BWP30P140LVT U1511 ( .A1(n14), .A2(i_data_bus[616]), .Z(N651) );
  CKAN2D1BWP30P140LVT U1512 ( .A1(n14), .A2(i_data_bus[617]), .Z(N652) );
  CKAN2D1BWP30P140LVT U1513 ( .A1(n14), .A2(i_data_bus[618]), .Z(N653) );
  CKAN2D1BWP30P140LVT U1514 ( .A1(n14), .A2(i_data_bus[619]), .Z(N654) );
  CKAN2D1BWP30P140LVT U1515 ( .A1(n14), .A2(i_data_bus[620]), .Z(N655) );
  CKAN2D1BWP30P140LVT U1516 ( .A1(n14), .A2(i_data_bus[621]), .Z(N656) );
  CKAN2D1BWP30P140LVT U1517 ( .A1(n14), .A2(i_data_bus[622]), .Z(N657) );
  CKAN2D1BWP30P140LVT U1518 ( .A1(n14), .A2(i_data_bus[623]), .Z(N658) );
  CKAN2D1BWP30P140LVT U1519 ( .A1(n14), .A2(i_data_bus[624]), .Z(N659) );
  CKAN2D1BWP30P140LVT U1520 ( .A1(n14), .A2(i_data_bus[625]), .Z(N660) );
  CKAN2D1BWP30P140LVT U1521 ( .A1(n14), .A2(i_data_bus[626]), .Z(N661) );
  CKAN2D1BWP30P140LVT U1522 ( .A1(n14), .A2(i_data_bus[627]), .Z(N662) );
  CKAN2D1BWP30P140LVT U1523 ( .A1(n14), .A2(i_data_bus[628]), .Z(N663) );
  CKAN2D1BWP30P140LVT U1524 ( .A1(n14), .A2(i_data_bus[629]), .Z(N664) );
  CKAN2D1BWP30P140LVT U1525 ( .A1(n14), .A2(i_data_bus[630]), .Z(N665) );
  CKAN2D1BWP30P140LVT U1526 ( .A1(n14), .A2(i_data_bus[631]), .Z(N666) );
  CKAN2D1BWP30P140LVT U1527 ( .A1(n14), .A2(i_data_bus[632]), .Z(N667) );
  CKAN2D1BWP30P140LVT U1528 ( .A1(n14), .A2(i_data_bus[633]), .Z(N668) );
  CKAN2D1BWP30P140LVT U1529 ( .A1(n14), .A2(i_data_bus[634]), .Z(N669) );
  CKAN2D1BWP30P140LVT U1530 ( .A1(n14), .A2(i_data_bus[635]), .Z(N670) );
  CKAN2D1BWP30P140LVT U1531 ( .A1(n14), .A2(i_data_bus[636]), .Z(N671) );
  CKAN2D1BWP30P140LVT U1532 ( .A1(n14), .A2(i_data_bus[637]), .Z(N672) );
  CKAN2D1BWP30P140LVT U1533 ( .A1(n14), .A2(i_data_bus[638]), .Z(N673) );
  CKAN2D1BWP30P140LVT U1534 ( .A1(n14), .A2(i_data_bus[639]), .Z(N674) );
  CKAN2D1BWP30P140LVT U1535 ( .A1(n14), .A2(i_data_bus[640]), .Z(N675) );
  CKAN2D1BWP30P140LVT U1536 ( .A1(n14), .A2(i_data_bus[641]), .Z(N676) );
  CKAN2D1BWP30P140LVT U1537 ( .A1(n14), .A2(i_data_bus[642]), .Z(N677) );
  CKAN2D1BWP30P140LVT U1538 ( .A1(n14), .A2(i_data_bus[643]), .Z(N678) );
  CKAN2D1BWP30P140LVT U1539 ( .A1(n14), .A2(i_data_bus[652]), .Z(N687) );
  CKAN2D1BWP30P140LVT U1540 ( .A1(n14), .A2(i_data_bus[653]), .Z(N688) );
  CKAN2D1BWP30P140LVT U1541 ( .A1(n14), .A2(i_data_bus[654]), .Z(N689) );
  CKAN2D1BWP30P140LVT U1542 ( .A1(n14), .A2(i_data_bus[655]), .Z(N690) );
  CKAN2D1BWP30P140LVT U1543 ( .A1(n14), .A2(i_data_bus[661]), .Z(N696) );
  CKAN2D1BWP30P140LVT U1544 ( .A1(n14), .A2(i_data_bus[662]), .Z(N697) );
  CKAN2D1BWP30P140LVT U1545 ( .A1(n14), .A2(i_data_bus[663]), .Z(N698) );
  CKAN2D1BWP30P140LVT U1546 ( .A1(n14), .A2(i_data_bus[664]), .Z(N699) );
  CKAN2D1BWP30P140LVT U1547 ( .A1(n14), .A2(i_data_bus[665]), .Z(N700) );
  CKAN2D1BWP30P140LVT U1548 ( .A1(n14), .A2(i_data_bus[666]), .Z(N701) );
  CKAN2D1BWP30P140LVT U1549 ( .A1(n14), .A2(i_data_bus[667]), .Z(N702) );
  CKAN2D1BWP30P140LVT U1550 ( .A1(n14), .A2(i_data_bus[673]), .Z(N708) );
  CKAN2D1BWP30P140LVT U1551 ( .A1(n14), .A2(i_data_bus[674]), .Z(N709) );
  CKAN2D1BWP30P140LVT U1552 ( .A1(n14), .A2(i_data_bus[675]), .Z(N710) );
  CKAN2D1BWP30P140LVT U1553 ( .A1(n14), .A2(i_data_bus[676]), .Z(N711) );
  CKAN2D1BWP30P140LVT U1554 ( .A1(n14), .A2(i_data_bus[677]), .Z(N712) );
  CKAN2D1BWP30P140LVT U1555 ( .A1(n14), .A2(i_data_bus[678]), .Z(N713) );
  CKAN2D1BWP30P140LVT U1556 ( .A1(n14), .A2(i_data_bus[679]), .Z(N714) );
  CKAN2D1BWP30P140LVT U1557 ( .A1(n14), .A2(i_data_bus[681]), .Z(N716) );
  CKAN2D1BWP30P140LVT U1558 ( .A1(n14), .A2(i_data_bus[682]), .Z(N717) );
  CKAN2D1BWP30P140LVT U1559 ( .A1(n14), .A2(i_data_bus[683]), .Z(N718) );
  CKAN2D1BWP30P140LVT U1560 ( .A1(n14), .A2(i_data_bus[684]), .Z(N719) );
  CKAN2D1BWP30P140LVT U1561 ( .A1(n14), .A2(i_data_bus[685]), .Z(N720) );
  CKAN2D1BWP30P140LVT U1562 ( .A1(n14), .A2(i_data_bus[686]), .Z(N721) );
  CKAN2D1BWP30P140LVT U1563 ( .A1(n14), .A2(i_data_bus[687]), .Z(N722) );
  CKAN2D1BWP30P140LVT U1564 ( .A1(n14), .A2(i_data_bus[688]), .Z(N723) );
  CKAN2D1BWP30P140LVT U1565 ( .A1(n14), .A2(i_data_bus[689]), .Z(N724) );
  CKAN2D1BWP30P140LVT U1566 ( .A1(n14), .A2(i_data_bus[690]), .Z(N725) );
  CKAN2D1BWP30P140LVT U1567 ( .A1(n14), .A2(i_data_bus[691]), .Z(N726) );
  CKAN2D1BWP30P140LVT U1568 ( .A1(n14), .A2(i_data_bus[692]), .Z(N727) );
  CKAN2D1BWP30P140LVT U1569 ( .A1(n14), .A2(i_data_bus[693]), .Z(N728) );
  CKAN2D1BWP30P140LVT U1570 ( .A1(n14), .A2(i_data_bus[694]), .Z(N729) );
  CKAN2D1BWP30P140LVT U1571 ( .A1(n14), .A2(i_data_bus[695]), .Z(N730) );
  CKAN2D1BWP30P140LVT U1572 ( .A1(n14), .A2(i_data_bus[696]), .Z(N731) );
  CKAN2D1BWP30P140LVT U1573 ( .A1(n14), .A2(i_data_bus[697]), .Z(N732) );
  CKAN2D1BWP30P140LVT U1574 ( .A1(n14), .A2(i_data_bus[698]), .Z(N733) );
  CKAN2D1BWP30P140LVT U1575 ( .A1(n14), .A2(i_data_bus[699]), .Z(N734) );
  CKAN2D1BWP30P140LVT U1576 ( .A1(n14), .A2(i_data_bus[700]), .Z(N735) );
  CKAN2D1BWP30P140LVT U1577 ( .A1(n14), .A2(i_data_bus[701]), .Z(N736) );
  CKAN2D1BWP30P140LVT U1578 ( .A1(n14), .A2(i_data_bus[702]), .Z(N737) );
  CKAN2D1BWP30P140LVT U1579 ( .A1(n14), .A2(i_data_bus[703]), .Z(N738) );
  CKAN2D1BWP30P140LVT U1580 ( .A1(n14), .A2(i_data_bus[704]), .Z(N739) );
  CKAN2D1BWP30P140LVT U1581 ( .A1(n14), .A2(i_data_bus[705]), .Z(N740) );
  CKAN2D1BWP30P140LVT U1582 ( .A1(n14), .A2(i_data_bus[706]), .Z(N741) );
  CKAN2D1BWP30P140LVT U1583 ( .A1(n14), .A2(i_data_bus[707]), .Z(N742) );
  CKAN2D1BWP30P140LVT U1584 ( .A1(n14), .A2(i_data_bus[708]), .Z(N743) );
  CKAN2D1BWP30P140LVT U1585 ( .A1(n14), .A2(i_data_bus[709]), .Z(N744) );
  CKAN2D1BWP30P140LVT U1586 ( .A1(n14), .A2(i_data_bus[710]), .Z(N745) );
  CKAN2D1BWP30P140LVT U1587 ( .A1(n14), .A2(i_data_bus[711]), .Z(N746) );
  CKAN2D1BWP30P140LVT U1588 ( .A1(n14), .A2(i_data_bus[712]), .Z(N747) );
  CKAN2D1BWP30P140LVT U1589 ( .A1(n14), .A2(i_data_bus[713]), .Z(N748) );
  CKAN2D1BWP30P140LVT U1590 ( .A1(n14), .A2(i_data_bus[714]), .Z(N749) );
  CKAN2D1BWP30P140LVT U1591 ( .A1(n14), .A2(i_data_bus[715]), .Z(N750) );
  CKAN2D1BWP30P140LVT U1592 ( .A1(n14), .A2(i_data_bus[724]), .Z(N759) );
  CKAN2D1BWP30P140LVT U1593 ( .A1(n14), .A2(i_data_bus[725]), .Z(N760) );
  CKAN2D1BWP30P140LVT U1594 ( .A1(n14), .A2(i_data_bus[726]), .Z(N761) );
  CKAN2D1BWP30P140LVT U1595 ( .A1(n14), .A2(i_data_bus[727]), .Z(N762) );
  CKAN2D1BWP30P140LVT U1596 ( .A1(n14), .A2(i_data_bus[733]), .Z(N768) );
  CKAN2D1BWP30P140LVT U1597 ( .A1(n14), .A2(i_data_bus[734]), .Z(N769) );
  CKAN2D1BWP30P140LVT U1598 ( .A1(n14), .A2(i_data_bus[735]), .Z(N770) );
  CKAN2D1BWP30P140LVT U1599 ( .A1(n14), .A2(i_data_bus[736]), .Z(N771) );
  CKAN2D1BWP30P140LVT U1600 ( .A1(n14), .A2(i_data_bus[737]), .Z(N772) );
  CKAN2D1BWP30P140LVT U1601 ( .A1(n14), .A2(i_data_bus[738]), .Z(N773) );
  CKAN2D1BWP30P140LVT U1602 ( .A1(n14), .A2(i_data_bus[739]), .Z(N774) );
  CKAN2D1BWP30P140LVT U1603 ( .A1(n14), .A2(i_data_bus[890]), .Z(N925) );
  CKAN2D1BWP30P140LVT U1604 ( .A1(n14), .A2(i_data_bus[891]), .Z(N926) );
  CKAN2D1BWP30P140LVT U1605 ( .A1(n14), .A2(i_data_bus[892]), .Z(N927) );
  CKAN2D1BWP30P140LVT U1606 ( .A1(n14), .A2(i_data_bus[893]), .Z(N928) );
  CKAN2D1BWP30P140LVT U1607 ( .A1(n14), .A2(i_data_bus[894]), .Z(N929) );
  CKAN2D1BWP30P140LVT U1608 ( .A1(n14), .A2(i_data_bus[895]), .Z(N930) );
  CKAN2D1BWP30P140LVT U1609 ( .A1(n14), .A2(i_data_bus[956]), .Z(N991) );
  CKAN2D1BWP30P140LVT U1610 ( .A1(n14), .A2(i_data_bus[957]), .Z(N992) );
  CKAN2D1BWP30P140LVT U1611 ( .A1(n14), .A2(i_data_bus[958]), .Z(N993) );
  CKAN2D1BWP30P140LVT U1612 ( .A1(n14), .A2(i_data_bus[959]), .Z(N994) );
  CKAN2D1BWP30P140LVT U1613 ( .A1(n14), .A2(i_data_bus[960]), .Z(N995) );
  CKAN2D1BWP30P140LVT U1614 ( .A1(n14), .A2(i_data_bus[968]), .Z(N1003) );
  CKAN2D1BWP30P140LVT U1615 ( .A1(n15), .A2(i_cmd[145]), .Z(N1204) );
  CKAN2D1BWP30P140LVT U1616 ( .A1(n15), .A2(i_cmd[146]), .Z(N1205) );
  CKAN2D1BWP30P140LVT U1617 ( .A1(n15), .A2(i_cmd[147]), .Z(N1206) );
  CKAN2D1BWP30P140LVT U1618 ( .A1(n15), .A2(i_cmd[148]), .Z(N1207) );
  CKAN2D1BWP30P140LVT U1619 ( .A1(n15), .A2(i_cmd[149]), .Z(N1208) );
  CKAN2D1BWP30P140LVT U1620 ( .A1(n15), .A2(i_cmd[150]), .Z(N1209) );
  CKAN2D1BWP30P140LVT U1621 ( .A1(n15), .A2(i_cmd[151]), .Z(N1210) );
  CKAN2D1BWP30P140LVT U1622 ( .A1(n15), .A2(i_cmd[152]), .Z(N1211) );
  CKAN2D1BWP30P140LVT U1623 ( .A1(n15), .A2(i_cmd[153]), .Z(N1212) );
  CKAN2D1BWP30P140LVT U1624 ( .A1(n15), .A2(i_cmd[154]), .Z(N1213) );
  CKAN2D1BWP30P140LVT U1625 ( .A1(n15), .A2(i_cmd[155]), .Z(N1214) );
  CKAN2D1BWP30P140LVT U1626 ( .A1(n15), .A2(i_cmd[156]), .Z(N1215) );
  CKAN2D1BWP30P140LVT U1627 ( .A1(n15), .A2(i_cmd[157]), .Z(N1216) );
  CKAN2D1BWP30P140LVT U1628 ( .A1(n15), .A2(i_cmd[158]), .Z(N1217) );
  CKAN2D1BWP30P140LVT U1629 ( .A1(n15), .A2(i_cmd[159]), .Z(N1218) );
  CKAN2D1BWP30P140LVT U1630 ( .A1(n15), .A2(i_cmd[160]), .Z(N1219) );
  CKAN2D1BWP30P140LVT U1631 ( .A1(n15), .A2(i_cmd[161]), .Z(N1220) );
  CKAN2D1BWP30P140LVT U1632 ( .A1(n15), .A2(i_cmd[162]), .Z(N1221) );
  CKAN2D1BWP30P140LVT U1633 ( .A1(n15), .A2(i_cmd[163]), .Z(N1222) );
  CKAN2D1BWP30P140LVT U1634 ( .A1(n15), .A2(i_cmd[164]), .Z(N1223) );
  CKAN2D1BWP30P140LVT U1635 ( .A1(n15), .A2(i_cmd[165]), .Z(N1224) );
  CKAN2D1BWP30P140LVT U1636 ( .A1(n15), .A2(i_cmd[166]), .Z(N1225) );
  CKAN2D1BWP30P140LVT U1637 ( .A1(n15), .A2(i_cmd[167]), .Z(N1226) );
  CKAN2D1BWP30P140LVT U1638 ( .A1(n15), .A2(i_cmd[168]), .Z(N1227) );
  CKAN2D1BWP30P140LVT U1639 ( .A1(n15), .A2(i_cmd[169]), .Z(N1228) );
  CKAN2D1BWP30P140LVT U1640 ( .A1(n15), .A2(i_cmd[170]), .Z(N1229) );
  CKAN2D1BWP30P140LVT U1641 ( .A1(n15), .A2(i_cmd[171]), .Z(N1230) );
  CKAN2D1BWP30P140LVT U1642 ( .A1(n15), .A2(i_cmd[172]), .Z(N1231) );
  CKAN2D1BWP30P140LVT U1643 ( .A1(n15), .A2(i_cmd[173]), .Z(N1232) );
  CKAN2D1BWP30P140LVT U1644 ( .A1(n15), .A2(i_cmd[174]), .Z(N1233) );
  CKAN2D1BWP30P140LVT U1645 ( .A1(n15), .A2(i_cmd[175]), .Z(N1234) );
  CKAN2D1BWP30P140LVT U1646 ( .A1(n15), .A2(i_cmd[176]), .Z(N1235) );
  CKAN2D1BWP30P140LVT U1647 ( .A1(n15), .A2(i_cmd[177]), .Z(N1236) );
  CKAN2D1BWP30P140LVT U1648 ( .A1(n15), .A2(i_cmd[178]), .Z(N1237) );
  CKAN2D1BWP30P140LVT U1649 ( .A1(n15), .A2(i_cmd[179]), .Z(N1238) );
  CKAN2D1BWP30P140LVT U1650 ( .A1(n15), .A2(i_cmd[188]), .Z(N1247) );
  CKAN2D1BWP30P140LVT U1651 ( .A1(n15), .A2(i_cmd[189]), .Z(N1248) );
  CKAN2D1BWP30P140LVT U1652 ( .A1(n15), .A2(i_cmd[190]), .Z(N1249) );
  CKAN2D1BWP30P140LVT U1653 ( .A1(n15), .A2(i_cmd[191]), .Z(N1250) );
  CKAN2D1BWP30P140LVT U1654 ( .A1(n15), .A2(i_cmd[197]), .Z(N1256) );
  CKAN2D1BWP30P140LVT U1655 ( .A1(n15), .A2(i_cmd[198]), .Z(N1257) );
  CKAN2D1BWP30P140LVT U1656 ( .A1(n15), .A2(i_cmd[199]), .Z(N1258) );
  CKAN2D1BWP30P140LVT U1657 ( .A1(n15), .A2(i_cmd[200]), .Z(N1259) );
  CKAN2D1BWP30P140LVT U1658 ( .A1(n15), .A2(i_cmd[201]), .Z(N1260) );
  CKAN2D1BWP30P140LVT U1659 ( .A1(n15), .A2(i_cmd[202]), .Z(N1261) );
  CKAN2D1BWP30P140LVT U1660 ( .A1(n15), .A2(i_cmd[203]), .Z(N1262) );
  CKAN2D1BWP30P140LVT U1661 ( .A1(n15), .A2(i_cmd[217]), .Z(N1276) );
  CKAN2D1BWP30P140LVT U1662 ( .A1(n15), .A2(i_cmd[218]), .Z(N1277) );
  CKAN2D1BWP30P140LVT U1663 ( .A1(n15), .A2(i_cmd[219]), .Z(N1278) );
  CKAN2D1BWP30P140LVT U1664 ( .A1(n15), .A2(i_cmd[220]), .Z(N1279) );
  CKAN2D1BWP30P140LVT U1665 ( .A1(n15), .A2(i_cmd[221]), .Z(N1280) );
  CKAN2D1BWP30P140LVT U1666 ( .A1(n15), .A2(i_cmd[222]), .Z(N1281) );
  CKAN2D1BWP30P140LVT U1667 ( .A1(n15), .A2(i_cmd[223]), .Z(N1282) );
  CKAN2D1BWP30P140LVT U1668 ( .A1(n15), .A2(i_cmd[224]), .Z(N1283) );
  CKAN2D1BWP30P140LVT U1669 ( .A1(n15), .A2(i_cmd[225]), .Z(N1284) );
  CKAN2D1BWP30P140LVT U1670 ( .A1(n15), .A2(i_cmd[226]), .Z(N1285) );
  CKAN2D1BWP30P140LVT U1671 ( .A1(n15), .A2(i_cmd[227]), .Z(N1286) );
  CKAN2D1BWP30P140LVT U1672 ( .A1(n15), .A2(i_cmd[228]), .Z(N1287) );
  CKAN2D1BWP30P140LVT U1673 ( .A1(n15), .A2(i_cmd[229]), .Z(N1288) );
  CKAN2D1BWP30P140LVT U1674 ( .A1(n15), .A2(i_cmd[230]), .Z(N1289) );
  CKAN2D1BWP30P140LVT U1675 ( .A1(n15), .A2(i_cmd[231]), .Z(N1290) );
  CKAN2D1BWP30P140LVT U1676 ( .A1(n15), .A2(i_cmd[232]), .Z(N1291) );
  CKAN2D1BWP30P140LVT U1677 ( .A1(n15), .A2(i_cmd[233]), .Z(N1292) );
  CKAN2D1BWP30P140LVT U1678 ( .A1(n15), .A2(i_cmd[234]), .Z(N1293) );
  CKAN2D1BWP30P140LVT U1679 ( .A1(n15), .A2(i_cmd[235]), .Z(N1294) );
  CKAN2D1BWP30P140LVT U1680 ( .A1(n15), .A2(i_cmd[236]), .Z(N1295) );
  CKAN2D1BWP30P140LVT U1681 ( .A1(n15), .A2(i_cmd[237]), .Z(N1296) );
  CKAN2D1BWP30P140LVT U1682 ( .A1(n15), .A2(i_cmd[238]), .Z(N1297) );
  CKAN2D1BWP30P140LVT U1683 ( .A1(n15), .A2(i_cmd[239]), .Z(N1298) );
  CKAN2D1BWP30P140LVT U1684 ( .A1(n15), .A2(i_cmd[240]), .Z(N1299) );
  CKAN2D1BWP30P140LVT U1685 ( .A1(n15), .A2(i_cmd[241]), .Z(N1300) );
  CKAN2D1BWP30P140LVT U1686 ( .A1(n15), .A2(i_cmd[242]), .Z(N1301) );
  CKAN2D1BWP30P140LVT U1687 ( .A1(n15), .A2(i_cmd[243]), .Z(N1302) );
  CKAN2D1BWP30P140LVT U1688 ( .A1(n15), .A2(i_cmd[244]), .Z(N1303) );
  CKAN2D1BWP30P140LVT U1689 ( .A1(n15), .A2(i_cmd[245]), .Z(N1304) );
  CKAN2D1BWP30P140LVT U1690 ( .A1(n15), .A2(i_cmd[246]), .Z(N1305) );
  CKAN2D1BWP30P140LVT U1691 ( .A1(n15), .A2(i_cmd[247]), .Z(N1306) );
  CKAN2D1BWP30P140LVT U1692 ( .A1(n15), .A2(i_cmd[248]), .Z(N1307) );
  CKAN2D1BWP30P140LVT U1693 ( .A1(n15), .A2(i_cmd[249]), .Z(N1308) );
  CKAN2D1BWP30P140LVT U1694 ( .A1(n15), .A2(i_cmd[250]), .Z(N1309) );
  CKAN2D1BWP30P140LVT U1695 ( .A1(n15), .A2(i_cmd[251]), .Z(N1310) );
  CKBD1BWP30P140LVT U1696 ( .I(n15), .Z(n8) );
  CKBD1BWP30P140LVT U1697 ( .I(n15), .Z(n9) );
  CKBD1BWP30P140LVT U1698 ( .I(n15), .Z(n10) );
  CKBD1BWP30P140LVT U1699 ( .I(n15), .Z(n7) );
  CKBD1BWP30P140LVT U1700 ( .I(n15), .Z(n13) );
  CKBD1BWP30P140LVT U1701 ( .I(n15), .Z(n11) );
  CKAN2D1BWP30P140LVT U1702 ( .A1(n12), .A2(i_data_bus[789]), .Z(N824) );
  CKAN2D1BWP30P140LVT U1703 ( .A1(n12), .A2(i_data_bus[847]), .Z(N882) );
  CKAN2D1BWP30P140LVT U1704 ( .A1(n12), .A2(i_data_bus[803]), .Z(N838) );
  CKAN2D1BWP30P140LVT U1705 ( .A1(n12), .A2(i_cmd[112]), .Z(N1171) );
  CKAN2D1BWP30P140LVT U1706 ( .A1(n12), .A2(i_data_bus[790]), .Z(N825) );
  CKAN2D1BWP30P140LVT U1707 ( .A1(n13), .A2(i_data_bus[801]), .Z(N836) );
  CKAN2D1BWP30P140LVT U1708 ( .A1(n14), .A2(i_data_bus[793]), .Z(N828) );
  CKAN2D1BWP30P140LVT U1709 ( .A1(n12), .A2(i_data_bus[788]), .Z(N823) );
  CKAN2D1BWP30P140LVT U1710 ( .A1(n12), .A2(i_cmd[69]), .Z(N1128) );
  CKAN2D1BWP30P140LVT U1711 ( .A1(n13), .A2(i_data_bus[841]), .Z(N876) );
  CKAN2D1BWP30P140LVT U1712 ( .A1(n14), .A2(i_data_bus[839]), .Z(N874) );
  CKAN2D1BWP30P140LVT U1713 ( .A1(n12), .A2(i_data_bus[802]), .Z(N837) );
  CKAN2D1BWP30P140LVT U1714 ( .A1(n12), .A2(i_cmd[40]), .Z(N1099) );
  CKAN2D1BWP30P140LVT U1715 ( .A1(n13), .A2(i_data_bus[804]), .Z(N839) );
  CKAN2D1BWP30P140LVT U1716 ( .A1(n14), .A2(i_cmd[12]), .Z(N1071) );
  CKAN2D1BWP30P140LVT U1717 ( .A1(n12), .A2(i_data_bus[792]), .Z(N827) );
  CKAN2D1BWP30P140LVT U1718 ( .A1(n12), .A2(i_data_bus[837]), .Z(N872) );
  CKAN2D1BWP30P140LVT U1719 ( .A1(n13), .A2(i_data_bus[843]), .Z(N878) );
  CKAN2D1BWP30P140LVT U1720 ( .A1(n12), .A2(i_data_bus[826]), .Z(N861) );
  CKAN2D1BWP30P140LVT U1721 ( .A1(n12), .A2(i_data_bus[791]), .Z(N826) );
  CKAN2D1BWP30P140LVT U1722 ( .A1(n12), .A2(i_cmd[0]), .Z(N1059) );
  CKAN2D1BWP30P140LVT U1723 ( .A1(n13), .A2(i_data_bus[800]), .Z(N835) );
  CKAN2D1BWP30P140LVT U1724 ( .A1(n14), .A2(i_data_bus[830]), .Z(N865) );
  CKAN2D1BWP30P140LVT U1725 ( .A1(n12), .A2(i_data_bus[795]), .Z(N830) );
  CKAN2D1BWP30P140LVT U1726 ( .A1(n12), .A2(i_data_bus[845]), .Z(N880) );
  CKAN2D1BWP30P140LVT U1727 ( .A1(n13), .A2(i_data_bus[828]), .Z(N863) );
  CKAN2D1BWP30P140LVT U1728 ( .A1(n14), .A2(i_cmd[59]), .Z(N1118) );
  CKAN2D1BWP30P140LVT U1729 ( .A1(n12), .A2(i_data_bus[794]), .Z(N829) );
  CKAN2D1BWP30P140LVT U1730 ( .A1(n9), .A2(i_data_bus[817]), .Z(N852) );
  CKAN2D1BWP30P140LVT U1731 ( .A1(n13), .A2(i_data_bus[844]), .Z(N879) );
  CKAN2D1BWP30P140LVT U1732 ( .A1(n11), .A2(i_data_bus[821]), .Z(N856) );
  CKAN2D1BWP30P140LVT U1733 ( .A1(n7), .A2(i_data_bus[752]), .Z(N787) );
  CKAN2D1BWP30P140LVT U1734 ( .A1(n10), .A2(i_data_bus[820]), .Z(N855) );
  CKAN2D1BWP30P140LVT U1735 ( .A1(n8), .A2(i_data_bus[819]), .Z(N854) );
  CKAN2D1BWP30P140LVT U1736 ( .A1(n9), .A2(i_data_bus[825]), .Z(N860) );
  CKAN2D1BWP30P140LVT U1737 ( .A1(n13), .A2(i_data_bus[842]), .Z(N877) );
  CKAN2D1BWP30P140LVT U1738 ( .A1(n11), .A2(i_data_bus[846]), .Z(N881) );
  CKAN2D1BWP30P140LVT U1739 ( .A1(n7), .A2(i_data_bus[840]), .Z(N875) );
  CKAN2D1BWP30P140LVT U1740 ( .A1(n10), .A2(i_data_bus[829]), .Z(N864) );
  CKAN2D1BWP30P140LVT U1741 ( .A1(n8), .A2(i_data_bus[822]), .Z(N857) );
  CKAN2D1BWP30P140LVT U1742 ( .A1(n9), .A2(i_data_bus[823]), .Z(N858) );
  CKAN2D1BWP30P140LVT U1743 ( .A1(n13), .A2(i_data_bus[838]), .Z(N873) );
  CKAN2D1BWP30P140LVT U1744 ( .A1(n11), .A2(i_data_bus[818]), .Z(N853) );
  CKAN2D1BWP30P140LVT U1745 ( .A1(n7), .A2(i_data_bus[740]), .Z(N775) );
  CKAN2D1BWP30P140LVT U1746 ( .A1(n10), .A2(i_data_bus[741]), .Z(N776) );
  CKAN2D1BWP30P140LVT U1747 ( .A1(n8), .A2(i_data_bus[742]), .Z(N777) );
  CKAN2D1BWP30P140LVT U1748 ( .A1(n9), .A2(i_data_bus[743]), .Z(N778) );
  CKAN2D1BWP30P140LVT U1749 ( .A1(n13), .A2(i_data_bus[744]), .Z(N779) );
  CKAN2D1BWP30P140LVT U1750 ( .A1(n11), .A2(i_data_bus[827]), .Z(N862) );
  CKAN2D1BWP30P140LVT U1751 ( .A1(n7), .A2(i_cmd[58]), .Z(N1117) );
  CKAN2D1BWP30P140LVT U1752 ( .A1(n10), .A2(i_data_bus[836]), .Z(N871) );
  CKAN2D1BWP30P140LVT U1753 ( .A1(n8), .A2(i_cmd[41]), .Z(N1100) );
  CKAN2D1BWP30P140LVT U1754 ( .A1(n9), .A2(i_cmd[24]), .Z(N1083) );
  CKAN2D1BWP30P140LVT U1755 ( .A1(n13), .A2(i_cmd[68]), .Z(N1127) );
  CKAN2D1BWP30P140LVT U1756 ( .A1(n11), .A2(i_cmd[64]), .Z(N1123) );
  CKAN2D1BWP30P140LVT U1757 ( .A1(n7), .A2(i_cmd[113]), .Z(N1172) );
  CKAN2D1BWP30P140LVT U1758 ( .A1(n7), .A2(i_cmd[23]), .Z(N1082) );
  CKAN2D1BWP30P140LVT U1759 ( .A1(n7), .A2(i_cmd[54]), .Z(N1113) );
  CKAN2D1BWP30P140LVT U1760 ( .A1(n7), .A2(i_cmd[28]), .Z(N1087) );
  CKAN2D1BWP30P140LVT U1761 ( .A1(n7), .A2(i_cmd[11]), .Z(N1070) );
  CKAN2D1BWP30P140LVT U1762 ( .A1(n7), .A2(i_cmd[94]), .Z(N1153) );
  CKAN2D1BWP30P140LVT U1763 ( .A1(n7), .A2(i_data_bus[812]), .Z(N847) );
  CKAN2D1BWP30P140LVT U1764 ( .A1(n7), .A2(i_data_bus[750]), .Z(N785) );
  CKAN2D1BWP30P140LVT U1765 ( .A1(n7), .A2(i_data_bus[815]), .Z(N850) );
  CKAN2D1BWP30P140LVT U1766 ( .A1(n7), .A2(i_cmd[70]), .Z(N1129) );
  CKAN2D1BWP30P140LVT U1767 ( .A1(n7), .A2(i_data_bus[814]), .Z(N849) );
  CKAN2D1BWP30P140LVT U1768 ( .A1(n7), .A2(i_cmd[104]), .Z(N1163) );
  CKAN2D1BWP30P140LVT U1769 ( .A1(n7), .A2(i_data_bus[751]), .Z(N786) );
  CKAN2D1BWP30P140LVT U1770 ( .A1(n7), .A2(i_cmd[126]), .Z(N1185) );
  CKAN2D1BWP30P140LVT U1771 ( .A1(n7), .A2(i_data_bus[749]), .Z(N784) );
  CKAN2D1BWP30P140LVT U1772 ( .A1(n7), .A2(i_cmd[60]), .Z(N1119) );
  CKAN2D1BWP30P140LVT U1773 ( .A1(n7), .A2(i_cmd[106]), .Z(N1165) );
  CKAN2D1BWP30P140LVT U1774 ( .A1(n7), .A2(i_data_bus[813]), .Z(N848) );
  CKAN2D1BWP30P140LVT U1775 ( .A1(n7), .A2(i_data_bus[747]), .Z(N782) );
  CKAN2D1BWP30P140LVT U1776 ( .A1(n7), .A2(i_data_bus[746]), .Z(N781) );
  CKAN2D1BWP30P140LVT U1777 ( .A1(n7), .A2(i_cmd[100]), .Z(N1159) );
  CKAN2D1BWP30P140LVT U1778 ( .A1(n7), .A2(i_cmd[118]), .Z(N1177) );
  CKAN2D1BWP30P140LVT U1779 ( .A1(n7), .A2(i_data_bus[816]), .Z(N851) );
  CKAN2D1BWP30P140LVT U1780 ( .A1(n7), .A2(i_cmd[98]), .Z(N1157) );
  CKAN2D1BWP30P140LVT U1781 ( .A1(n7), .A2(i_data_bus[824]), .Z(N859) );
  CKAN2D1BWP30P140LVT U1782 ( .A1(n7), .A2(i_cmd[96]), .Z(N1155) );
  CKAN2D1BWP30P140LVT U1783 ( .A1(n7), .A2(i_data_bus[748]), .Z(N783) );
  CKAN2D1BWP30P140LVT U1784 ( .A1(n7), .A2(i_cmd[130]), .Z(N1189) );
  CKAN2D1BWP30P140LVT U1785 ( .A1(n7), .A2(i_cmd[102]), .Z(N1161) );
  CKAN2D1BWP30P140LVT U1786 ( .A1(n7), .A2(i_cmd[116]), .Z(N1175) );
  CKAN2D1BWP30P140LVT U1787 ( .A1(n7), .A2(i_cmd[119]), .Z(N1178) );
  CKAN2D1BWP30P140LVT U1788 ( .A1(n9), .A2(i_cmd[55]), .Z(N1114) );
  CKAN2D1BWP30P140LVT U1789 ( .A1(n13), .A2(i_cmd[44]), .Z(N1103) );
  CKAN2D1BWP30P140LVT U1790 ( .A1(n11), .A2(i_cmd[93]), .Z(N1152) );
  CKAN2D1BWP30P140LVT U1791 ( .A1(n7), .A2(i_cmd[61]), .Z(N1120) );
  CKAN2D1BWP30P140LVT U1792 ( .A1(n10), .A2(i_cmd[27]), .Z(N1086) );
  CKAN2D1BWP30P140LVT U1793 ( .A1(n8), .A2(i_cmd[97]), .Z(N1156) );
  CKAN2D1BWP30P140LVT U1794 ( .A1(n9), .A2(i_cmd[107]), .Z(N1166) );
  CKAN2D1BWP30P140LVT U1795 ( .A1(n13), .A2(i_cmd[71]), .Z(N1130) );
  CKAN2D1BWP30P140LVT U1796 ( .A1(n11), .A2(i_cmd[99]), .Z(N1158) );
  CKAN2D1BWP30P140LVT U1797 ( .A1(n7), .A2(i_cmd[117]), .Z(N1176) );
  CKAN2D1BWP30P140LVT U1798 ( .A1(n10), .A2(i_cmd[101]), .Z(N1160) );
  CKAN2D1BWP30P140LVT U1799 ( .A1(n8), .A2(i_cmd[82]), .Z(N1141) );
  CKAN2D1BWP30P140LVT U1800 ( .A1(n9), .A2(i_cmd[103]), .Z(N1162) );
  CKAN2D1BWP30P140LVT U1801 ( .A1(n13), .A2(i_cmd[127]), .Z(N1186) );
  CKAN2D1BWP30P140LVT U1802 ( .A1(n11), .A2(i_cmd[105]), .Z(N1164) );
  CKAN2D1BWP30P140LVT U1803 ( .A1(n7), .A2(i_cmd[131]), .Z(N1190) );
  CKAN2D1BWP30P140LVT U1804 ( .A1(n10), .A2(i_data_bus[864]), .Z(N899) );
  CKAN2D1BWP30P140LVT U1805 ( .A1(n8), .A2(i_data_bus[861]), .Z(N896) );
  CKAN2D1BWP30P140LVT U1806 ( .A1(n9), .A2(i_data_bus[866]), .Z(N901) );
  CKAN2D1BWP30P140LVT U1807 ( .A1(n13), .A2(i_data_bus[867]), .Z(N902) );
  CKAN2D1BWP30P140LVT U1808 ( .A1(n11), .A2(i_data_bus[875]), .Z(N910) );
  CKAN2D1BWP30P140LVT U1809 ( .A1(n7), .A2(i_data_bus[863]), .Z(N898) );
  CKAN2D1BWP30P140LVT U1810 ( .A1(n10), .A2(i_data_bus[862]), .Z(N897) );
  CKAN2D1BWP30P140LVT U1811 ( .A1(n8), .A2(i_data_bus[873]), .Z(N908) );
  CKAN2D1BWP30P140LVT U1812 ( .A1(n9), .A2(i_data_bus[874]), .Z(N909) );
  CKAN2D1BWP30P140LVT U1813 ( .A1(n13), .A2(i_data_bus[860]), .Z(N895) );
  CKAN2D1BWP30P140LVT U1814 ( .A1(n11), .A2(i_data_bus[876]), .Z(N911) );
  CKAN2D1BWP30P140LVT U1815 ( .A1(n7), .A2(i_data_bus[865]), .Z(N900) );
  CKAN2D1BWP30P140LVT U1816 ( .A1(n10), .A2(i_data_bus[872]), .Z(N907) );
  CKAN2D1BWP30P140LVT U1817 ( .A1(n11), .A2(i_valid[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U1818 ( .A1(n13), .A2(i_valid[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U1819 ( .A1(n8), .A2(i_valid[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U1820 ( .A1(n11), .A2(i_valid[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U1821 ( .A1(n10), .A2(i_cmd[2]), .Z(N1061) );
  CKAN2D1BWP30P140LVT U1822 ( .A1(n14), .A2(i_valid[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U1823 ( .A1(n9), .A2(i_valid[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U1824 ( .A1(n8), .A2(i_cmd[5]), .Z(N1064) );
  CKAN2D1BWP30P140LVT U1825 ( .A1(n10), .A2(i_valid[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U1826 ( .A1(n10), .A2(i_cmd[143]), .Z(N1202) );
  CKAN2D1BWP30P140LVT U1827 ( .A1(n9), .A2(i_cmd[15]), .Z(N1074) );
  CKAN2D1BWP30P140LVT U1828 ( .A1(n11), .A2(i_cmd[4]), .Z(N1063) );
  CKAN2D1BWP30P140LVT U1829 ( .A1(n8), .A2(i_cmd[17]), .Z(N1076) );
  CKAN2D1BWP30P140LVT U1830 ( .A1(n10), .A2(i_valid[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U1831 ( .A1(n14), .A2(i_valid[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U1832 ( .A1(n7), .A2(i_valid[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U1833 ( .A1(n9), .A2(i_cmd[3]), .Z(N1062) );
  CKAN2D1BWP30P140LVT U1834 ( .A1(n8), .A2(i_valid[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U1835 ( .A1(n8), .A2(i_cmd[34]), .Z(N1093) );
  CKAN2D1BWP30P140LVT U1836 ( .A1(n11), .A2(i_cmd[35]), .Z(N1094) );
  CKAN2D1BWP30P140LVT U1837 ( .A1(n11), .A2(i_cmd[36]), .Z(N1095) );
  CKAN2D1BWP30P140LVT U1838 ( .A1(n9), .A2(i_cmd[37]), .Z(N1096) );
  CKAN2D1BWP30P140LVT U1839 ( .A1(n10), .A2(i_cmd[38]), .Z(N1097) );
  CKAN2D1BWP30P140LVT U1840 ( .A1(n9), .A2(i_valid[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U1841 ( .A1(n8), .A2(i_cmd[43]), .Z(N1102) );
  CKAN2D1BWP30P140LVT U1842 ( .A1(n8), .A2(i_valid[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U1843 ( .A1(n9), .A2(i_cmd[45]), .Z(N1104) );
  CKAN2D1BWP30P140LVT U1844 ( .A1(n10), .A2(i_cmd[46]), .Z(N1105) );
  CKAN2D1BWP30P140LVT U1845 ( .A1(n8), .A2(i_cmd[48]), .Z(N1107) );
  CKAN2D1BWP30P140LVT U1846 ( .A1(n8), .A2(i_data_bus[859]), .Z(N894) );
  CKAN2D1BWP30P140LVT U1847 ( .A1(n10), .A2(i_data_bus[757]), .Z(N792) );
  CKAN2D1BWP30P140LVT U1848 ( .A1(n7), .A2(i_cmd[56]), .Z(N1115) );
  CKAN2D1BWP30P140LVT U1849 ( .A1(n8), .A2(i_data_bus[756]), .Z(N791) );
  CKAN2D1BWP30P140LVT U1850 ( .A1(n11), .A2(i_data_bus[755]), .Z(N790) );
  CKAN2D1BWP30P140LVT U1851 ( .A1(n10), .A2(i_cmd[14]), .Z(N1073) );
  CKAN2D1BWP30P140LVT U1852 ( .A1(n9), .A2(i_data_bus[754]), .Z(N789) );
  CKAN2D1BWP30P140LVT U1853 ( .A1(n11), .A2(i_cmd[16]), .Z(N1075) );
  CKAN2D1BWP30P140LVT U1854 ( .A1(n11), .A2(i_cmd[62]), .Z(N1121) );
  CKAN2D1BWP30P140LVT U1855 ( .A1(n11), .A2(i_data_bus[1015]), .Z(N1050) );
  CKAN2D1BWP30P140LVT U1856 ( .A1(n14), .A2(i_data_bus[1023]), .Z(N1058) );
  CKAN2D1BWP30P140LVT U1857 ( .A1(n13), .A2(i_cmd[26]), .Z(N1085) );
  CKAN2D1BWP30P140LVT U1858 ( .A1(n9), .A2(i_valid[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U1859 ( .A1(n10), .A2(i_data_bus[753]), .Z(N788) );
  CKAN2D1BWP30P140LVT U1860 ( .A1(n8), .A2(i_cmd[77]), .Z(N1136) );
  CKAN2D1BWP30P140LVT U1861 ( .A1(n8), .A2(i_data_bus[1014]), .Z(N1049) );
  CKAN2D1BWP30P140LVT U1862 ( .A1(n11), .A2(i_cmd[78]), .Z(N1137) );
  CKAN2D1BWP30P140LVT U1863 ( .A1(n9), .A2(i_cmd[79]), .Z(N1138) );
  CKAN2D1BWP30P140LVT U1864 ( .A1(n10), .A2(i_cmd[80]), .Z(N1139) );
  CKAN2D1BWP30P140LVT U1865 ( .A1(n8), .A2(i_cmd[86]), .Z(N1145) );
  CKAN2D1BWP30P140LVT U1866 ( .A1(n11), .A2(i_cmd[87]), .Z(N1146) );
  CKAN2D1BWP30P140LVT U1867 ( .A1(n9), .A2(i_cmd[88]), .Z(N1147) );
  CKAN2D1BWP30P140LVT U1868 ( .A1(n8), .A2(i_data_bus[745]), .Z(N780) );
  CKAN2D1BWP30P140LVT U1869 ( .A1(n10), .A2(i_cmd[216]), .Z(N1275) );
  CKAN2D1BWP30P140LVT U1870 ( .A1(n9), .A2(i_cmd[215]), .Z(N1274) );
  CKAN2D1BWP30P140LVT U1871 ( .A1(n10), .A2(i_cmd[89]), .Z(N1148) );
  CKAN2D1BWP30P140LVT U1872 ( .A1(n8), .A2(i_cmd[92]), .Z(N1151) );
  CKAN2D1BWP30P140LVT U1873 ( .A1(n9), .A2(i_cmd[214]), .Z(N1273) );
  CKAN2D1BWP30P140LVT U1874 ( .A1(n9), .A2(i_cmd[213]), .Z(N1272) );
  CKAN2D1BWP30P140LVT U1875 ( .A1(n9), .A2(i_cmd[212]), .Z(N1271) );
  CKAN2D1BWP30P140LVT U1876 ( .A1(n9), .A2(i_cmd[211]), .Z(N1270) );
  CKAN2D1BWP30P140LVT U1877 ( .A1(n9), .A2(i_cmd[210]), .Z(N1269) );
  CKAN2D1BWP30P140LVT U1878 ( .A1(n9), .A2(i_cmd[209]), .Z(N1268) );
  CKAN2D1BWP30P140LVT U1879 ( .A1(n10), .A2(i_cmd[208]), .Z(N1267) );
  CKAN2D1BWP30P140LVT U1880 ( .A1(n10), .A2(i_cmd[207]), .Z(N1266) );
  CKAN2D1BWP30P140LVT U1881 ( .A1(n10), .A2(i_cmd[206]), .Z(N1265) );
  CKAN2D1BWP30P140LVT U1882 ( .A1(n10), .A2(i_cmd[205]), .Z(N1264) );
  CKAN2D1BWP30P140LVT U1883 ( .A1(n10), .A2(i_cmd[204]), .Z(N1263) );
  CKAN2D1BWP30P140LVT U1884 ( .A1(n11), .A2(i_cmd[196]), .Z(N1255) );
  CKAN2D1BWP30P140LVT U1885 ( .A1(n11), .A2(i_cmd[195]), .Z(N1254) );
  CKAN2D1BWP30P140LVT U1886 ( .A1(n11), .A2(i_cmd[194]), .Z(N1253) );
  CKAN2D1BWP30P140LVT U1887 ( .A1(n11), .A2(i_cmd[193]), .Z(N1252) );
  CKAN2D1BWP30P140LVT U1888 ( .A1(n11), .A2(i_cmd[108]), .Z(N1167) );
  CKAN2D1BWP30P140LVT U1889 ( .A1(n9), .A2(i_cmd[109]), .Z(N1168) );
  CKAN2D1BWP30P140LVT U1890 ( .A1(n10), .A2(i_cmd[110]), .Z(N1169) );
  CKAN2D1BWP30P140LVT U1891 ( .A1(n11), .A2(i_cmd[192]), .Z(N1251) );
  CKAN2D1BWP30P140LVT U1892 ( .A1(n10), .A2(i_cmd[115]), .Z(N1174) );
  CKAN2D1BWP30P140LVT U1893 ( .A1(n11), .A2(i_cmd[187]), .Z(N1246) );
  CKAN2D1BWP30P140LVT U1894 ( .A1(n11), .A2(i_cmd[186]), .Z(N1245) );
  CKAN2D1BWP30P140LVT U1895 ( .A1(n11), .A2(i_cmd[185]), .Z(N1244) );
  CKAN2D1BWP30P140LVT U1896 ( .A1(n11), .A2(i_cmd[184]), .Z(N1243) );
  CKAN2D1BWP30P140LVT U1897 ( .A1(n8), .A2(i_cmd[124]), .Z(N1183) );
  CKAN2D1BWP30P140LVT U1898 ( .A1(n7), .A2(i_cmd[125]), .Z(N1184) );
  CKAN2D1BWP30P140LVT U1899 ( .A1(n11), .A2(i_cmd[182]), .Z(N1241) );
  CKAN2D1BWP30P140LVT U1900 ( .A1(n11), .A2(i_cmd[181]), .Z(N1240) );
  CKAN2D1BWP30P140LVT U1901 ( .A1(n11), .A2(i_cmd[129]), .Z(N1188) );
  CKAN2D1BWP30P140LVT U1902 ( .A1(n11), .A2(i_cmd[180]), .Z(N1239) );
  CKAN2D1BWP30P140LVT U1903 ( .A1(n9), .A2(i_cmd[144]), .Z(N1203) );
  CKAN2D1BWP30P140LVT U1904 ( .A1(n9), .A2(i_cmd[132]), .Z(N1191) );
  CKAN2D1BWP30P140LVT U1905 ( .A1(n9), .A2(i_cmd[133]), .Z(N1192) );
  CKAN2D1BWP30P140LVT U1906 ( .A1(n9), .A2(i_cmd[134]), .Z(N1193) );
  CKAN2D1BWP30P140LVT U1907 ( .A1(n9), .A2(i_cmd[135]), .Z(N1194) );
  CKAN2D1BWP30P140LVT U1908 ( .A1(n9), .A2(i_cmd[136]), .Z(N1195) );
  CKAN2D1BWP30P140LVT U1909 ( .A1(n10), .A2(i_cmd[137]), .Z(N1196) );
  CKAN2D1BWP30P140LVT U1910 ( .A1(n10), .A2(i_cmd[138]), .Z(N1197) );
  CKAN2D1BWP30P140LVT U1911 ( .A1(n10), .A2(i_cmd[139]), .Z(N1198) );
  CKAN2D1BWP30P140LVT U1912 ( .A1(n10), .A2(i_cmd[140]), .Z(N1199) );
  CKAN2D1BWP30P140LVT U1913 ( .A1(n10), .A2(i_cmd[141]), .Z(N1200) );
  CKAN2D1BWP30P140LVT U1914 ( .A1(n10), .A2(i_cmd[142]), .Z(N1201) );
  CKAN2D1BWP30P140LVT U1915 ( .A1(n11), .A2(i_cmd[183]), .Z(N1242) );
  CKAN2D1BWP30P140LVT U1916 ( .A1(n9), .A2(i_data_bus[869]), .Z(N904) );
  CKAN2D1BWP30P140LVT U1917 ( .A1(n10), .A2(i_data_bus[870]), .Z(N905) );
  CKAN2D1BWP30P140LVT U1918 ( .A1(n13), .A2(i_data_bus[858]), .Z(N893) );
  CKAN2D1BWP30P140LVT U1919 ( .A1(n10), .A2(i_data_bus[850]), .Z(N885) );
  CKAN2D1BWP30P140LVT U1920 ( .A1(n9), .A2(i_data_bus[849]), .Z(N884) );
  CKAN2D1BWP30P140LVT U1921 ( .A1(n11), .A2(i_data_bus[848]), .Z(N883) );
  CKAN2D1BWP30P140LVT U1922 ( .A1(n9), .A2(i_data_bus[882]), .Z(N917) );
  CKAN2D1BWP30P140LVT U1923 ( .A1(n8), .A2(i_data_bus[883]), .Z(N918) );
  CKAN2D1BWP30P140LVT U1924 ( .A1(n11), .A2(i_data_bus[889]), .Z(N924) );
  CKAN2D1BWP30P140LVT U1925 ( .A1(n11), .A2(i_data_bus[897]), .Z(N932) );
  CKAN2D1BWP30P140LVT U1926 ( .A1(n8), .A2(i_data_bus[898]), .Z(N933) );
  CKAN2D1BWP30P140LVT U1927 ( .A1(n8), .A2(i_data_bus[899]), .Z(N934) );
  CKAN2D1BWP30P140LVT U1928 ( .A1(n13), .A2(i_data_bus[900]), .Z(N935) );
  CKAN2D1BWP30P140LVT U1929 ( .A1(n11), .A2(i_data_bus[868]), .Z(N903) );
  CKAN2D1BWP30P140LVT U1930 ( .A1(n14), .A2(i_data_bus[908]), .Z(N943) );
  CKAN2D1BWP30P140LVT U1931 ( .A1(n10), .A2(i_data_bus[918]), .Z(N953) );
  CKAN2D1BWP30P140LVT U1932 ( .A1(n9), .A2(i_data_bus[919]), .Z(N954) );
  CKAN2D1BWP30P140LVT U1933 ( .A1(n10), .A2(i_data_bus[920]), .Z(N955) );
  CKAN2D1BWP30P140LVT U1934 ( .A1(n9), .A2(i_data_bus[921]), .Z(N956) );
  CKAN2D1BWP30P140LVT U1935 ( .A1(n14), .A2(i_data_bus[922]), .Z(N957) );
  CKAN2D1BWP30P140LVT U1936 ( .A1(n10), .A2(i_data_bus[940]), .Z(N975) );
  CKAN2D1BWP30P140LVT U1937 ( .A1(n9), .A2(i_data_bus[941]), .Z(N976) );
  CKAN2D1BWP30P140LVT U1938 ( .A1(n11), .A2(i_data_bus[942]), .Z(N977) );
  CKAN2D1BWP30P140LVT U1939 ( .A1(n8), .A2(i_data_bus[943]), .Z(N978) );
  CKAN2D1BWP30P140LVT U1940 ( .A1(n10), .A2(i_data_bus[952]), .Z(N987) );
  CKAN2D1BWP30P140LVT U1941 ( .A1(n8), .A2(i_data_bus[156]), .Z(N191) );
  CKAN2D1BWP30P140LVT U1942 ( .A1(n8), .A2(i_data_bus[155]), .Z(N190) );
  CKAN2D1BWP30P140LVT U1943 ( .A1(n8), .A2(i_data_bus[154]), .Z(N189) );
  CKAN2D1BWP30P140LVT U1944 ( .A1(n8), .A2(i_data_bus[153]), .Z(N188) );
  CKAN2D1BWP30P140LVT U1945 ( .A1(n8), .A2(i_data_bus[152]), .Z(N187) );
  CKAN2D1BWP30P140LVT U1946 ( .A1(n8), .A2(i_data_bus[147]), .Z(N182) );
  CKAN2D1BWP30P140LVT U1947 ( .A1(n8), .A2(i_data_bus[146]), .Z(N181) );
  CKAN2D1BWP30P140LVT U1948 ( .A1(n8), .A2(i_data_bus[145]), .Z(N180) );
  CKAN2D1BWP30P140LVT U1949 ( .A1(n8), .A2(i_data_bus[144]), .Z(N179) );
  CKAN2D1BWP30P140LVT U1950 ( .A1(n8), .A2(i_data_bus[143]), .Z(N178) );
  CKAN2D1BWP30P140LVT U1951 ( .A1(n8), .A2(i_data_bus[142]), .Z(N177) );
  CKAN2D1BWP30P140LVT U1952 ( .A1(n8), .A2(i_data_bus[141]), .Z(N176) );
  CKAN2D1BWP30P140LVT U1953 ( .A1(n8), .A2(i_data_bus[140]), .Z(N175) );
  CKAN2D1BWP30P140LVT U1954 ( .A1(n14), .A2(i_data_bus[127]), .Z(N162) );
  CKAN2D1BWP30P140LVT U1955 ( .A1(n8), .A2(i_data_bus[126]), .Z(N161) );
  CKAN2D1BWP30P140LVT U1956 ( .A1(n14), .A2(i_data_bus[125]), .Z(N160) );
  CKAN2D1BWP30P140LVT U1957 ( .A1(n10), .A2(i_data_bus[124]), .Z(N159) );
  CKAN2D1BWP30P140LVT U1958 ( .A1(n14), .A2(i_data_bus[123]), .Z(N158) );
  CKAN2D1BWP30P140LVT U1959 ( .A1(n7), .A2(i_data_bus[122]), .Z(N157) );
  CKAN2D1BWP30P140LVT U1960 ( .A1(n14), .A2(i_data_bus[121]), .Z(N156) );
  CKAN2D1BWP30P140LVT U1961 ( .A1(n11), .A2(i_data_bus[120]), .Z(N155) );
  CKAN2D1BWP30P140LVT U1962 ( .A1(n14), .A2(i_data_bus[119]), .Z(N154) );
  CKAN2D1BWP30P140LVT U1963 ( .A1(n13), .A2(i_data_bus[118]), .Z(N153) );
  CKAN2D1BWP30P140LVT U1964 ( .A1(n9), .A2(i_data_bus[758]), .Z(N793) );
  CKAN2D1BWP30P140LVT U1965 ( .A1(n10), .A2(i_data_bus[833]), .Z(N868) );
  CKAN2D1BWP30P140LVT U1966 ( .A1(n9), .A2(i_data_bus[832]), .Z(N867) );
  CKAN2D1BWP30P140LVT U1967 ( .A1(n13), .A2(i_data_bus[117]), .Z(N152) );
  CKAN2D1BWP30P140LVT U1968 ( .A1(n8), .A2(i_data_bus[116]), .Z(N151) );
  CKAN2D1BWP30P140LVT U1969 ( .A1(n14), .A2(i_data_bus[110]), .Z(N145) );
  CKAN2D1BWP30P140LVT U1970 ( .A1(n10), .A2(i_data_bus[109]), .Z(N144) );
  CKAN2D1BWP30P140LVT U1971 ( .A1(n11), .A2(i_data_bus[831]), .Z(N866) );
  CKAN2D1BWP30P140LVT U1972 ( .A1(n12), .A2(i_data_bus[108]), .Z(N143) );
  CKAN2D1BWP30P140LVT U1973 ( .A1(n12), .A2(i_data_bus[107]), .Z(N142) );
  CKAN2D1BWP30P140LVT U1974 ( .A1(n14), .A2(i_data_bus[106]), .Z(N141) );
  CKAN2D1BWP30P140LVT U1975 ( .A1(n7), .A2(i_data_bus[105]), .Z(N140) );
  CKAN2D1BWP30P140LVT U1976 ( .A1(n7), .A2(i_data_bus[104]), .Z(N139) );
  CKAN2D1BWP30P140LVT U1977 ( .A1(n11), .A2(i_data_bus[103]), .Z(N138) );
  CKAN2D1BWP30P140LVT U1978 ( .A1(n13), .A2(i_data_bus[102]), .Z(N137) );
  CKAN2D1BWP30P140LVT U1979 ( .A1(n9), .A2(i_data_bus[101]), .Z(N136) );
  CKAN2D1BWP30P140LVT U1980 ( .A1(n8), .A2(i_data_bus[100]), .Z(N135) );
  CKAN2D1BWP30P140LVT U1981 ( .A1(n10), .A2(i_data_bus[99]), .Z(N134) );
  CKAN2D1BWP30P140LVT U1982 ( .A1(n12), .A2(i_data_bus[98]), .Z(N133) );
  CKAN2D1BWP30P140LVT U1983 ( .A1(n7), .A2(i_data_bus[97]), .Z(N132) );
  CKAN2D1BWP30P140LVT U1984 ( .A1(n11), .A2(i_data_bus[96]), .Z(N131) );
  CKAN2D1BWP30P140LVT U1985 ( .A1(n13), .A2(i_data_bus[95]), .Z(N130) );
  CKAN2D1BWP30P140LVT U1986 ( .A1(n9), .A2(i_data_bus[94]), .Z(N129) );
  CKAN2D1BWP30P140LVT U1987 ( .A1(n8), .A2(i_data_bus[93]), .Z(N128) );
  CKAN2D1BWP30P140LVT U1988 ( .A1(n10), .A2(i_data_bus[92]), .Z(N127) );
  CKAN2D1BWP30P140LVT U1989 ( .A1(n12), .A2(i_data_bus[901]), .Z(N936) );
  CKAN2D1BWP30P140LVT U1990 ( .A1(n13), .A2(i_data_bus[84]), .Z(N119) );
  CKAN2D1BWP30P140LVT U1991 ( .A1(n14), .A2(i_data_bus[83]), .Z(N118) );
  CKAN2D1BWP30P140LVT U1992 ( .A1(n11), .A2(i_data_bus[82]), .Z(N117) );
  CKAN2D1BWP30P140LVT U1993 ( .A1(n9), .A2(i_data_bus[962]), .Z(N997) );
  CKAN2D1BWP30P140LVT U1994 ( .A1(n9), .A2(i_data_bus[811]), .Z(N846) );
  CKAN2D1BWP30P140LVT U1995 ( .A1(n10), .A2(i_data_bus[810]), .Z(N845) );
  CKAN2D1BWP30P140LVT U1996 ( .A1(n8), .A2(i_data_bus[964]), .Z(N999) );
  CKAN2D1BWP30P140LVT U1997 ( .A1(n12), .A2(i_data_bus[81]), .Z(N116) );
  CKAN2D1BWP30P140LVT U1998 ( .A1(n14), .A2(i_data_bus[80]), .Z(N115) );
  CKAN2D1BWP30P140LVT U1999 ( .A1(n7), .A2(i_data_bus[780]), .Z(N815) );
  CKAN2D1BWP30P140LVT U2000 ( .A1(n7), .A2(i_data_bus[75]), .Z(N110) );
  CKAN2D1BWP30P140LVT U2001 ( .A1(n12), .A2(i_data_bus[74]), .Z(N109) );
  CKAN2D1BWP30P140LVT U2002 ( .A1(n7), .A2(i_data_bus[73]), .Z(N108) );
  CKAN2D1BWP30P140LVT U2003 ( .A1(n7), .A2(i_data_bus[26]), .Z(N61) );
  CKAN2D1BWP30P140LVT U2004 ( .A1(n11), .A2(i_data_bus[72]), .Z(N107) );
  CKAN2D1BWP30P140LVT U2005 ( .A1(n13), .A2(i_data_bus[71]), .Z(N106) );
  CKAN2D1BWP30P140LVT U2006 ( .A1(n14), .A2(i_data_bus[70]), .Z(N105) );
  CKAN2D1BWP30P140LVT U2007 ( .A1(n10), .A2(i_data_bus[69]), .Z(N104) );
  CKAN2D1BWP30P140LVT U2008 ( .A1(n10), .A2(i_data_bus[68]), .Z(N103) );
  CKAN2D1BWP30P140LVT U2009 ( .A1(n9), .A2(i_data_bus[799]), .Z(N834) );
  CKAN2D1BWP30P140LVT U2010 ( .A1(n10), .A2(i_data_bus[798]), .Z(N833) );
  CKAN2D1BWP30P140LVT U2011 ( .A1(n11), .A2(i_data_bus[954]), .Z(N989) );
  CKAN2D1BWP30P140LVT U2012 ( .A1(n11), .A2(i_data_bus[32]), .Z(N67) );
  CKAN2D1BWP30P140LVT U2013 ( .A1(n10), .A2(i_data_bus[961]), .Z(N996) );
  CKAN2D1BWP30P140LVT U2014 ( .A1(n11), .A2(i_data_bus[31]), .Z(N66) );
  CKAN2D1BWP30P140LVT U2015 ( .A1(n13), .A2(i_data_bus[30]), .Z(N65) );
  CKAN2D1BWP30P140LVT U2016 ( .A1(n9), .A2(i_data_bus[29]), .Z(N64) );
  CKAN2D1BWP30P140LVT U2017 ( .A1(n8), .A2(i_data_bus[28]), .Z(N63) );
  CKAN2D1BWP30P140LVT U2018 ( .A1(n12), .A2(i_data_bus[759]), .Z(N794) );
  CKAN2D1BWP30P140LVT U2019 ( .A1(n10), .A2(i_data_bus[27]), .Z(N62) );
  CKAN2D1BWP30P140LVT U2020 ( .A1(n13), .A2(i_data_bus[765]), .Z(N800) );
  CKAN2D1BWP30P140LVT U2021 ( .A1(n9), .A2(i_data_bus[24]), .Z(N59) );
  CKAN2D1BWP30P140LVT U2022 ( .A1(n8), .A2(i_data_bus[23]), .Z(N58) );
  CKAN2D1BWP30P140LVT U2023 ( .A1(n10), .A2(i_data_bus[22]), .Z(N57) );
  CKAN2D1BWP30P140LVT U2024 ( .A1(n12), .A2(i_data_bus[990]), .Z(N1025) );
  CKAN2D1BWP30P140LVT U2025 ( .A1(n7), .A2(i_data_bus[21]), .Z(N56) );
  CKAN2D1BWP30P140LVT U2026 ( .A1(n11), .A2(i_data_bus[20]), .Z(N55) );
  CKAN2D1BWP30P140LVT U2027 ( .A1(n9), .A2(i_data_bus[953]), .Z(N988) );
  CKAN2D1BWP30P140LVT U2028 ( .A1(n11), .A2(i_data_bus[970]), .Z(N1005) );
  CKAN2D1BWP30P140LVT U2029 ( .A1(n8), .A2(i_data_bus[955]), .Z(N990) );
  CKAN2D1BWP30P140LVT U2030 ( .A1(n9), .A2(i_data_bus[971]), .Z(N1006) );
  CKAN2D1BWP30P140LVT U2031 ( .A1(n10), .A2(i_data_bus[972]), .Z(N1007) );
  CKAN2D1BWP30P140LVT U2032 ( .A1(n11), .A2(i_data_bus[963]), .Z(N998) );
  CKAN2D1BWP30P140LVT U2033 ( .A1(n14), .A2(i_data_bus[1003]), .Z(N1038) );
  CKAN2D1BWP30P140LVT U2034 ( .A1(n13), .A2(i_data_bus[1012]), .Z(N1047) );
  CKAN2D1BWP30P140LVT U2035 ( .A1(n7), .A2(i_data_bus[1013]), .Z(N1048) );
  CKAN2D1BWP30P140LVT U2036 ( .A1(n11), .A2(i_data_bus[965]), .Z(N1000) );
  CKAN2D1BWP30P140LVT U2037 ( .A1(n8), .A2(i_data_bus[969]), .Z(N1004) );
  CKAN2D1BWP30P140LVT U2038 ( .A1(n9), .A2(i_data_bus[779]), .Z(N814) );
  CKAN2D1BWP30P140LVT U2039 ( .A1(n13), .A2(i_data_bus[778]), .Z(N813) );
  CKAN2D1BWP30P140LVT U2040 ( .A1(n8), .A2(i_data_bus[777]), .Z(N812) );
  CKAN2D1BWP30P140LVT U2041 ( .A1(n9), .A2(i_data_bus[992]), .Z(N1027) );
  CKAN2D1BWP30P140LVT U2042 ( .A1(n10), .A2(i_data_bus[993]), .Z(N1028) );
  CKAN2D1BWP30P140LVT U2043 ( .A1(n11), .A2(i_data_bus[776]), .Z(N811) );
  CKAN2D1BWP30P140LVT U2044 ( .A1(n8), .A2(i_data_bus[989]), .Z(N1024) );
  CKAN2D1BWP30P140LVT U2045 ( .A1(n9), .A2(i_data_bus[764]), .Z(N799) );
  CKAN2D1BWP30P140LVT U2046 ( .A1(n8), .A2(i_data_bus[991]), .Z(N1026) );
  CKAN2D1BWP30P140LVT U2047 ( .A1(n8), .A2(i_data_bus[766]), .Z(N801) );
  CKAN2D1BWP30P140LVT U2048 ( .A1(n12), .A2(i_data_bus[797]), .Z(N832) );
  CKAN2D1BWP30P140LVT U2049 ( .A1(n12), .A2(i_data_bus[775]), .Z(N810) );
  CKAN2D1BWP30P140LVT U2050 ( .A1(n12), .A2(i_data_bus[917]), .Z(N952) );
  CKAN2D1BWP30P140LVT U2051 ( .A1(n12), .A2(i_cmd[111]), .Z(N1170) );
  CKAN2D1BWP30P140LVT U2052 ( .A1(n12), .A2(i_data_bus[834]), .Z(N869) );
  CKAN2D1BWP30P140LVT U2053 ( .A1(n12), .A2(i_data_bus[951]), .Z(N986) );
  CKAN2D1BWP30P140LVT U2054 ( .A1(n12), .A2(i_cmd[13]), .Z(N1072) );
  CKAN2D1BWP30P140LVT U2055 ( .A1(n12), .A2(i_valid[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U2056 ( .A1(n12), .A2(i_data_bus[973]), .Z(N1008) );
  CKAN2D1BWP30P140LVT U2057 ( .A1(n12), .A2(i_cmd[252]), .Z(N1311) );
  CKAN2D1BWP30P140LVT U2058 ( .A1(n12), .A2(i_data_bus[980]), .Z(N1015) );
  CKAN2D1BWP30P140LVT U2059 ( .A1(n12), .A2(i_cmd[81]), .Z(N1140) );
  CKAN2D1BWP30P140LVT U2060 ( .A1(n12), .A2(i_cmd[39]), .Z(N1098) );
  CKAN2D1BWP30P140LVT U2061 ( .A1(n12), .A2(i_data_bus[931]), .Z(N966) );
  CKAN2D1BWP30P140LVT U2062 ( .A1(n12), .A2(i_valid[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U2063 ( .A1(n12), .A2(i_cmd[90]), .Z(N1149) );
  CKAN2D1BWP30P140LVT U2064 ( .A1(n12), .A2(i_cmd[1]), .Z(N1060) );
  CKAN2D1BWP30P140LVT U2065 ( .A1(n12), .A2(i_cmd[253]), .Z(N1312) );
  CKAN2D1BWP30P140LVT U2066 ( .A1(n12), .A2(i_data_bus[851]), .Z(N886) );
  CKAN2D1BWP30P140LVT U2067 ( .A1(n12), .A2(i_data_bus[994]), .Z(N1029) );
  CKAN2D1BWP30P140LVT U2068 ( .A1(n12), .A2(i_data_bus[871]), .Z(N906) );
  CKAN2D1BWP30P140LVT U2069 ( .A1(n12), .A2(i_cmd[254]), .Z(N1313) );
  CKAN2D1BWP30P140LVT U2070 ( .A1(n12), .A2(i_data_bus[809]), .Z(N844) );
  CKAN2D1BWP30P140LVT U2071 ( .A1(n12), .A2(i_cmd[47]), .Z(N1106) );
  CKAN2D1BWP30P140LVT U2072 ( .A1(n12), .A2(i_cmd[255]), .Z(N1314) );
  CKAN2D1BWP30P140LVT U2073 ( .A1(n12), .A2(i_data_bus[12]), .Z(N47) );
  CKAN2D1BWP30P140LVT U2074 ( .A1(n12), .A2(i_data_bus[11]), .Z(N46) );
  CKAN2D1BWP30P140LVT U2075 ( .A1(n12), .A2(i_data_bus[10]), .Z(N45) );
  CKAN2D1BWP30P140LVT U2076 ( .A1(n12), .A2(i_data_bus[9]), .Z(N44) );
  CKAN2D1BWP30P140LVT U2077 ( .A1(n12), .A2(i_data_bus[8]), .Z(N43) );
  CKAN2D1BWP30P140LVT U2078 ( .A1(n12), .A2(i_data_bus[3]), .Z(N38) );
  CKAN2D1BWP30P140LVT U2079 ( .A1(n12), .A2(i_data_bus[2]), .Z(N37) );
  CKAN2D1BWP30P140LVT U2080 ( .A1(n12), .A2(i_data_bus[1]), .Z(N36) );
  CKAN2D1BWP30P140LVT U2081 ( .A1(n12), .A2(i_data_bus[0]), .Z(N35) );
  CKAN2D1BWP30P140LVT U2082 ( .A1(n8), .A2(i_data_bus[909]), .Z(N944) );
  CKAN2D1BWP30P140LVT U2083 ( .A1(n11), .A2(i_data_bus[910]), .Z(N945) );
  CKAN2D1BWP30P140LVT U2084 ( .A1(n9), .A2(i_data_bus[760]), .Z(N795) );
  CKAN2D1BWP30P140LVT U2085 ( .A1(n8), .A2(i_data_bus[360]), .Z(N395) );
  CKAN2D1BWP30P140LVT U2086 ( .A1(n9), .A2(i_data_bus[359]), .Z(N394) );
  CKAN2D1BWP30P140LVT U2087 ( .A1(n13), .A2(i_data_bus[358]), .Z(N393) );
  CKAN2D1BWP30P140LVT U2088 ( .A1(n13), .A2(i_data_bus[902]), .Z(N937) );
  CKAN2D1BWP30P140LVT U2089 ( .A1(n7), .A2(i_data_bus[903]), .Z(N938) );
  CKAN2D1BWP30P140LVT U2090 ( .A1(n14), .A2(i_data_bus[904]), .Z(N939) );
  CKAN2D1BWP30P140LVT U2091 ( .A1(n11), .A2(i_data_bus[905]), .Z(N940) );
  CKAN2D1BWP30P140LVT U2092 ( .A1(n10), .A2(i_data_bus[906]), .Z(N941) );
  CKAN2D1BWP30P140LVT U2093 ( .A1(n14), .A2(i_data_bus[907]), .Z(N942) );
  CKAN2D1BWP30P140LVT U2094 ( .A1(n7), .A2(i_data_bus[357]), .Z(N392) );
  CKAN2D1BWP30P140LVT U2095 ( .A1(n10), .A2(i_data_bus[316]), .Z(N351) );
  CKAN2D1BWP30P140LVT U2096 ( .A1(n11), .A2(i_data_bus[923]), .Z(N958) );
  CKAN2D1BWP30P140LVT U2097 ( .A1(n8), .A2(i_data_bus[924]), .Z(N959) );
  CKAN2D1BWP30P140LVT U2098 ( .A1(n14), .A2(i_data_bus[925]), .Z(N960) );
  CKAN2D1BWP30P140LVT U2099 ( .A1(n10), .A2(i_data_bus[926]), .Z(N961) );
  CKAN2D1BWP30P140LVT U2100 ( .A1(n12), .A2(i_data_bus[927]), .Z(N962) );
  CKAN2D1BWP30P140LVT U2101 ( .A1(n14), .A2(i_data_bus[928]), .Z(N963) );
  CKAN2D1BWP30P140LVT U2102 ( .A1(n13), .A2(i_data_bus[929]), .Z(N964) );
  CKAN2D1BWP30P140LVT U2103 ( .A1(n10), .A2(i_data_bus[930]), .Z(N965) );
  CKAN2D1BWP30P140LVT U2104 ( .A1(n9), .A2(i_data_bus[315]), .Z(N350) );
  CKAN2D1BWP30P140LVT U2105 ( .A1(n13), .A2(i_data_bus[314]), .Z(N349) );
  CKAN2D1BWP30P140LVT U2106 ( .A1(n11), .A2(i_data_bus[313]), .Z(N348) );
  CKAN2D1BWP30P140LVT U2107 ( .A1(n14), .A2(i_data_bus[312]), .Z(N347) );
  CKAN2D1BWP30P140LVT U2108 ( .A1(n14), .A2(i_data_bus[311]), .Z(N346) );
  CKAN2D1BWP30P140LVT U2109 ( .A1(n8), .A2(i_data_bus[949]), .Z(N984) );
  CKAN2D1BWP30P140LVT U2110 ( .A1(n8), .A2(i_data_bus[950]), .Z(N985) );
  CKAN2D1BWP30P140LVT U2111 ( .A1(n14), .A2(i_data_bus[310]), .Z(N345) );
  CKAN2D1BWP30P140LVT U2112 ( .A1(n14), .A2(i_data_bus[309]), .Z(N344) );
  CKAN2D1BWP30P140LVT U2113 ( .A1(n14), .A2(i_data_bus[308]), .Z(N343) );
  CKAN2D1BWP30P140LVT U2114 ( .A1(n14), .A2(i_data_bus[911]), .Z(N946) );
  CKAN2D1BWP30P140LVT U2115 ( .A1(n8), .A2(i_data_bus[912]), .Z(N947) );
  CKAN2D1BWP30P140LVT U2116 ( .A1(n8), .A2(i_data_bus[913]), .Z(N948) );
  CKAN2D1BWP30P140LVT U2117 ( .A1(n14), .A2(i_data_bus[914]), .Z(N949) );
  CKAN2D1BWP30P140LVT U2118 ( .A1(n9), .A2(i_data_bus[915]), .Z(N950) );
  CKAN2D1BWP30P140LVT U2119 ( .A1(n9), .A2(i_data_bus[916]), .Z(N951) );
  CKAN2D1BWP30P140LVT U2120 ( .A1(n9), .A2(i_data_bus[356]), .Z(N391) );
  CKAN2D1BWP30P140LVT U2121 ( .A1(n14), .A2(i_data_bus[320]), .Z(N355) );
  CKAN2D1BWP30P140LVT U2122 ( .A1(n7), .A2(i_data_bus[319]), .Z(N354) );
  CKAN2D1BWP30P140LVT U2123 ( .A1(n10), .A2(i_data_bus[318]), .Z(N353) );
  CKAN2D1BWP30P140LVT U2124 ( .A1(n8), .A2(i_data_bus[317]), .Z(N352) );
  CKAN2D1BWP30P140LVT U2125 ( .A1(n13), .A2(i_data_bus[974]), .Z(N1009) );
  CKAN2D1BWP30P140LVT U2126 ( .A1(n13), .A2(i_data_bus[975]), .Z(N1010) );
  CKAN2D1BWP30P140LVT U2127 ( .A1(n14), .A2(i_data_bus[976]), .Z(N1011) );
  CKAN2D1BWP30P140LVT U2128 ( .A1(n9), .A2(i_data_bus[977]), .Z(N1012) );
  CKAN2D1BWP30P140LVT U2129 ( .A1(n13), .A2(i_data_bus[978]), .Z(N1013) );
  CKAN2D1BWP30P140LVT U2130 ( .A1(n14), .A2(i_data_bus[979]), .Z(N1014) );
  CKAN2D1BWP30P140LVT U2131 ( .A1(n11), .A2(i_data_bus[981]), .Z(N1016) );
  CKAN2D1BWP30P140LVT U2132 ( .A1(n11), .A2(i_data_bus[982]), .Z(N1017) );
  CKAN2D1BWP30P140LVT U2133 ( .A1(n14), .A2(i_data_bus[983]), .Z(N1018) );
  CKAN2D1BWP30P140LVT U2134 ( .A1(n13), .A2(i_data_bus[984]), .Z(N1019) );
  CKAN2D1BWP30P140LVT U2135 ( .A1(n11), .A2(i_data_bus[985]), .Z(N1020) );
  CKAN2D1BWP30P140LVT U2136 ( .A1(n14), .A2(i_data_bus[986]), .Z(N1021) );
  CKAN2D1BWP30P140LVT U2137 ( .A1(n9), .A2(i_data_bus[987]), .Z(N1022) );
  CKAN2D1BWP30P140LVT U2138 ( .A1(n7), .A2(i_data_bus[988]), .Z(N1023) );
  CKAN2D1BWP30P140LVT U2139 ( .A1(n7), .A2(i_data_bus[995]), .Z(N1030) );
  CKAN2D1BWP30P140LVT U2140 ( .A1(n7), .A2(i_data_bus[361]), .Z(N396) );
  CKAN2D1BWP30P140LVT U2141 ( .A1(n7), .A2(i_data_bus[996]), .Z(N1031) );
  CKAN2D1BWP30P140LVT U2142 ( .A1(n14), .A2(i_data_bus[997]), .Z(N1032) );
  CKAN2D1BWP30P140LVT U2143 ( .A1(n11), .A2(i_data_bus[998]), .Z(N1033) );
  CKAN2D1BWP30P140LVT U2144 ( .A1(n10), .A2(i_data_bus[999]), .Z(N1034) );
  CKAN2D1BWP30P140LVT U2145 ( .A1(n14), .A2(i_data_bus[1000]), .Z(N1035) );
  CKAN2D1BWP30P140LVT U2146 ( .A1(n13), .A2(i_data_bus[1001]), .Z(N1036) );
  CKAN2D1BWP30P140LVT U2147 ( .A1(n10), .A2(i_data_bus[1002]), .Z(N1037) );
  CKAN2D1BWP30P140LVT U2148 ( .A1(n14), .A2(i_cmd[128]), .Z(N1187) );
  CKAN2D1BWP30P140LVT U2149 ( .A1(n8), .A2(i_cmd[123]), .Z(N1182) );
  CKAN2D1BWP30P140LVT U2150 ( .A1(n11), .A2(i_cmd[122]), .Z(N1181) );
  CKAN2D1BWP30P140LVT U2151 ( .A1(n14), .A2(i_cmd[121]), .Z(N1180) );
  CKAN2D1BWP30P140LVT U2152 ( .A1(n8), .A2(i_cmd[120]), .Z(N1179) );
  CKAN2D1BWP30P140LVT U2153 ( .A1(n7), .A2(i_data_bus[1021]), .Z(N1056) );
  CKAN2D1BWP30P140LVT U2154 ( .A1(n9), .A2(i_data_bus[1022]), .Z(N1057) );
  CKAN2D1BWP30P140LVT U2155 ( .A1(n14), .A2(i_cmd[114]), .Z(N1173) );
  CKAN2D1BWP30P140LVT U2156 ( .A1(n7), .A2(i_cmd[95]), .Z(N1154) );
  CKAN2D1BWP30P140LVT U2157 ( .A1(n14), .A2(i_cmd[91]), .Z(N1150) );
  CKAN2D1BWP30P140LVT U2158 ( .A1(n13), .A2(i_cmd[85]), .Z(N1144) );
  CKAN2D1BWP30P140LVT U2159 ( .A1(n12), .A2(i_valid[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U2160 ( .A1(n12), .A2(i_valid[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U2161 ( .A1(n14), .A2(i_valid[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U2162 ( .A1(n12), .A2(i_valid[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U2163 ( .A1(n9), .A2(i_valid[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U2164 ( .A1(n14), .A2(i_valid[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U2165 ( .A1(n10), .A2(i_valid[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U2166 ( .A1(n11), .A2(i_valid[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U2167 ( .A1(n8), .A2(i_cmd[84]), .Z(N1143) );
  CKAN2D1BWP30P140LVT U2168 ( .A1(n14), .A2(i_cmd[83]), .Z(N1142) );
  CKAN2D1BWP30P140LVT U2169 ( .A1(n7), .A2(i_cmd[76]), .Z(N1135) );
  CKAN2D1BWP30P140LVT U2170 ( .A1(n9), .A2(i_cmd[75]), .Z(N1134) );
  CKAN2D1BWP30P140LVT U2171 ( .A1(n14), .A2(i_cmd[74]), .Z(N1133) );
  CKAN2D1BWP30P140LVT U2172 ( .A1(n13), .A2(i_cmd[73]), .Z(N1132) );
  CKAN2D1BWP30P140LVT U2173 ( .A1(n10), .A2(i_cmd[72]), .Z(N1131) );
  CKAN2D1BWP30P140LVT U2174 ( .A1(n14), .A2(i_cmd[31]), .Z(N1090) );
  CKAN2D1BWP30P140LVT U2175 ( .A1(n10), .A2(i_valid[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U2176 ( .A1(n13), .A2(i_valid[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U2177 ( .A1(n14), .A2(i_valid[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U2178 ( .A1(n11), .A2(i_valid[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U2179 ( .A1(n12), .A2(i_valid[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U2180 ( .A1(n14), .A2(i_valid[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U2181 ( .A1(n7), .A2(i_cmd[66]), .Z(N1125) );
  CKAN2D1BWP30P140LVT U2182 ( .A1(n11), .A2(i_valid[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U2183 ( .A1(n12), .A2(i_valid[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U2184 ( .A1(n14), .A2(i_cmd[65]), .Z(N1124) );
  CKAN2D1BWP30P140LVT U2185 ( .A1(n14), .A2(i_cmd[63]), .Z(N1122) );
  CKAN2D1BWP30P140LVT U2186 ( .A1(n14), .A2(i_cmd[57]), .Z(N1116) );
  CKAN2D1BWP30P140LVT U2187 ( .A1(n8), .A2(i_cmd[53]), .Z(N1112) );
  CKAN2D1BWP30P140LVT U2188 ( .A1(n8), .A2(i_cmd[6]), .Z(N1065) );
  CKAN2D1BWP30P140LVT U2189 ( .A1(n11), .A2(i_cmd[7]), .Z(N1066) );
  CKAN2D1BWP30P140LVT U2190 ( .A1(n14), .A2(i_cmd[8]), .Z(N1067) );
  CKAN2D1BWP30P140LVT U2191 ( .A1(n10), .A2(i_cmd[9]), .Z(N1068) );
  CKAN2D1BWP30P140LVT U2192 ( .A1(n9), .A2(i_cmd[10]), .Z(N1069) );
  CKAN2D1BWP30P140LVT U2193 ( .A1(n8), .A2(i_cmd[52]), .Z(N1111) );
  CKAN2D1BWP30P140LVT U2194 ( .A1(n14), .A2(i_cmd[51]), .Z(N1110) );
  CKAN2D1BWP30P140LVT U2195 ( .A1(n7), .A2(i_cmd[50]), .Z(N1109) );
  CKAN2D1BWP30P140LVT U2196 ( .A1(n9), .A2(i_cmd[49]), .Z(N1108) );
  CKAN2D1BWP30P140LVT U2197 ( .A1(n14), .A2(i_cmd[42]), .Z(N1101) );
  CKAN2D1BWP30P140LVT U2198 ( .A1(n13), .A2(i_cmd[18]), .Z(N1077) );
  CKAN2D1BWP30P140LVT U2199 ( .A1(n10), .A2(i_cmd[19]), .Z(N1078) );
  CKAN2D1BWP30P140LVT U2200 ( .A1(n14), .A2(i_cmd[20]), .Z(N1079) );
  CKAN2D1BWP30P140LVT U2201 ( .A1(n9), .A2(i_cmd[21]), .Z(N1080) );
  CKAN2D1BWP30P140LVT U2202 ( .A1(n13), .A2(i_cmd[22]), .Z(N1081) );
  CKAN2D1BWP30P140LVT U2203 ( .A1(n14), .A2(i_cmd[25]), .Z(N1084) );
  CKAN2D1BWP30P140LVT U2204 ( .A1(n11), .A2(i_cmd[33]), .Z(N1092) );
  CKAN2D1BWP30P140LVT U2205 ( .A1(n8), .A2(i_cmd[32]), .Z(N1091) );
  CKAN2D1BWP30P140LVT U2206 ( .A1(n11), .A2(i_cmd[29]), .Z(N1088) );
  CKAN2D1BWP30P140LVT U2207 ( .A1(n13), .A2(i_cmd[30]), .Z(N1089) );
  CKAN2D1BWP30P140LVT U2208 ( .A1(n11), .A2(i_data_bus[362]), .Z(N397) );
  CKAN2D1BWP30P140LVT U2209 ( .A1(n14), .A2(i_data_bus[762]), .Z(N797) );
  CKAN2D1BWP30P140LVT U2210 ( .A1(n7), .A2(i_data_bus[763]), .Z(N798) );
  CKAN2D1BWP30P140LVT U2211 ( .A1(n7), .A2(i_data_bus[588]), .Z(N623) );
  CKAN2D1BWP30P140LVT U2212 ( .A1(n12), .A2(i_data_bus[587]), .Z(N622) );
  CKAN2D1BWP30P140LVT U2213 ( .A1(n10), .A2(i_data_bus[586]), .Z(N621) );
  CKAN2D1BWP30P140LVT U2214 ( .A1(n7), .A2(i_data_bus[767]), .Z(N802) );
  CKAN2D1BWP30P140LVT U2215 ( .A1(n9), .A2(i_data_bus[768]), .Z(N803) );
  CKAN2D1BWP30P140LVT U2216 ( .A1(n14), .A2(i_data_bus[769]), .Z(N804) );
  CKAN2D1BWP30P140LVT U2217 ( .A1(n10), .A2(i_data_bus[770]), .Z(N805) );
  CKAN2D1BWP30P140LVT U2218 ( .A1(n12), .A2(i_data_bus[771]), .Z(N806) );
  CKAN2D1BWP30P140LVT U2219 ( .A1(n14), .A2(i_data_bus[772]), .Z(N807) );
  CKAN2D1BWP30P140LVT U2220 ( .A1(n7), .A2(i_data_bus[773]), .Z(N808) );
  CKAN2D1BWP30P140LVT U2221 ( .A1(n10), .A2(i_data_bus[774]), .Z(N809) );
  CKAN2D1BWP30P140LVT U2222 ( .A1(n8), .A2(i_data_bus[585]), .Z(N620) );
  CKAN2D1BWP30P140LVT U2223 ( .A1(n9), .A2(i_data_bus[584]), .Z(N619) );
  CKAN2D1BWP30P140LVT U2224 ( .A1(n13), .A2(i_data_bus[579]), .Z(N614) );
  CKAN2D1BWP30P140LVT U2225 ( .A1(n11), .A2(i_data_bus[578]), .Z(N613) );
  CKAN2D1BWP30P140LVT U2226 ( .A1(n7), .A2(i_data_bus[577]), .Z(N612) );
  CKAN2D1BWP30P140LVT U2227 ( .A1(n12), .A2(i_data_bus[576]), .Z(N611) );
  CKAN2D1BWP30P140LVT U2228 ( .A1(n10), .A2(i_data_bus[781]), .Z(N816) );
  CKAN2D1BWP30P140LVT U2229 ( .A1(n13), .A2(i_data_bus[782]), .Z(N817) );
  CKAN2D1BWP30P140LVT U2230 ( .A1(n14), .A2(i_data_bus[783]), .Z(N818) );
  CKAN2D1BWP30P140LVT U2231 ( .A1(n8), .A2(i_data_bus[784]), .Z(N819) );
  CKAN2D1BWP30P140LVT U2232 ( .A1(n10), .A2(i_data_bus[785]), .Z(N820) );
  CKAN2D1BWP30P140LVT U2233 ( .A1(n14), .A2(i_data_bus[786]), .Z(N821) );
  CKAN2D1BWP30P140LVT U2234 ( .A1(n12), .A2(i_data_bus[787]), .Z(N822) );
  CKAN2D1BWP30P140LVT U2235 ( .A1(n12), .A2(i_data_bus[575]), .Z(N610) );
  CKAN2D1BWP30P140LVT U2236 ( .A1(n8), .A2(i_data_bus[574]), .Z(N609) );
  CKAN2D1BWP30P140LVT U2237 ( .A1(n9), .A2(i_data_bus[573]), .Z(N608) );
  CKAN2D1BWP30P140LVT U2238 ( .A1(n13), .A2(i_data_bus[572]), .Z(N607) );
  CKAN2D1BWP30P140LVT U2239 ( .A1(n8), .A2(i_data_bus[559]), .Z(N594) );
  CKAN2D1BWP30P140LVT U2240 ( .A1(n10), .A2(i_data_bus[558]), .Z(N593) );
  CKAN2D1BWP30P140LVT U2241 ( .A1(n9), .A2(i_data_bus[557]), .Z(N592) );
  CKAN2D1BWP30P140LVT U2242 ( .A1(n10), .A2(i_data_bus[556]), .Z(N591) );
  CKAN2D1BWP30P140LVT U2243 ( .A1(n13), .A2(i_data_bus[796]), .Z(N831) );
  CKAN2D1BWP30P140LVT U2244 ( .A1(n11), .A2(i_data_bus[555]), .Z(N590) );
  CKAN2D1BWP30P140LVT U2245 ( .A1(n8), .A2(i_data_bus[554]), .Z(N589) );
  CKAN2D1BWP30P140LVT U2246 ( .A1(n7), .A2(i_data_bus[553]), .Z(N588) );
  CKAN2D1BWP30P140LVT U2247 ( .A1(n9), .A2(i_data_bus[552]), .Z(N587) );
  CKAN2D1BWP30P140LVT U2248 ( .A1(n12), .A2(i_data_bus[551]), .Z(N586) );
  CKAN2D1BWP30P140LVT U2249 ( .A1(n13), .A2(i_data_bus[550]), .Z(N585) );
  CKAN2D1BWP30P140LVT U2250 ( .A1(n12), .A2(i_data_bus[549]), .Z(N584) );
  CKAN2D1BWP30P140LVT U2251 ( .A1(n11), .A2(i_data_bus[548]), .Z(N583) );
  CKAN2D1BWP30P140LVT U2252 ( .A1(n11), .A2(i_data_bus[805]), .Z(N840) );
  CKAN2D1BWP30P140LVT U2253 ( .A1(n14), .A2(i_data_bus[806]), .Z(N841) );
  CKAN2D1BWP30P140LVT U2254 ( .A1(n7), .A2(i_data_bus[807]), .Z(N842) );
  CKAN2D1BWP30P140LVT U2255 ( .A1(n10), .A2(i_data_bus[808]), .Z(N843) );
  CKAN2D1BWP30P140LVT U2256 ( .A1(n8), .A2(i_data_bus[542]), .Z(N577) );
  CKAN2D1BWP30P140LVT U2257 ( .A1(n12), .A2(i_data_bus[541]), .Z(N576) );
  CKAN2D1BWP30P140LVT U2258 ( .A1(n9), .A2(i_data_bus[540]), .Z(N575) );
  CKAN2D1BWP30P140LVT U2259 ( .A1(n8), .A2(i_data_bus[539]), .Z(N574) );
  CKAN2D1BWP30P140LVT U2260 ( .A1(n13), .A2(i_data_bus[538]), .Z(N573) );
  CKAN2D1BWP30P140LVT U2261 ( .A1(n9), .A2(i_data_bus[537]), .Z(N572) );
  CKAN2D1BWP30P140LVT U2262 ( .A1(n14), .A2(i_data_bus[536]), .Z(N571) );
  CKAN2D1BWP30P140LVT U2263 ( .A1(n12), .A2(i_data_bus[535]), .Z(N570) );
  CKAN2D1BWP30P140LVT U2264 ( .A1(n10), .A2(i_data_bus[534]), .Z(N569) );
  CKAN2D1BWP30P140LVT U2265 ( .A1(n13), .A2(i_data_bus[533]), .Z(N568) );
  CKAN2D1BWP30P140LVT U2266 ( .A1(n13), .A2(i_data_bus[532]), .Z(N567) );
  CKAN2D1BWP30P140LVT U2267 ( .A1(n11), .A2(i_data_bus[531]), .Z(N566) );
  CKAN2D1BWP30P140LVT U2268 ( .A1(n7), .A2(i_data_bus[530]), .Z(N565) );
  CKAN2D1BWP30P140LVT U2269 ( .A1(n11), .A2(i_data_bus[529]), .Z(N564) );
  CKAN2D1BWP30P140LVT U2270 ( .A1(n14), .A2(i_data_bus[528]), .Z(N563) );
  CKAN2D1BWP30P140LVT U2271 ( .A1(n14), .A2(i_data_bus[527]), .Z(N562) );
  CKAN2D1BWP30P140LVT U2272 ( .A1(n14), .A2(i_data_bus[526]), .Z(N561) );
  CKAN2D1BWP30P140LVT U2273 ( .A1(n14), .A2(i_data_bus[525]), .Z(N560) );
  CKAN2D1BWP30P140LVT U2274 ( .A1(n14), .A2(i_data_bus[524]), .Z(N559) );
  CKAN2D1BWP30P140LVT U2275 ( .A1(n11), .A2(i_data_bus[516]), .Z(N551) );
  CKAN2D1BWP30P140LVT U2276 ( .A1(n7), .A2(i_data_bus[515]), .Z(N550) );
  CKAN2D1BWP30P140LVT U2277 ( .A1(n12), .A2(i_data_bus[514]), .Z(N549) );
  CKAN2D1BWP30P140LVT U2278 ( .A1(n12), .A2(i_data_bus[513]), .Z(N548) );
  CKAN2D1BWP30P140LVT U2279 ( .A1(n10), .A2(i_data_bus[512]), .Z(N547) );
  CKAN2D1BWP30P140LVT U2280 ( .A1(n8), .A2(i_data_bus[507]), .Z(N542) );
  CKAN2D1BWP30P140LVT U2281 ( .A1(n9), .A2(i_data_bus[506]), .Z(N541) );
  CKAN2D1BWP30P140LVT U2282 ( .A1(n14), .A2(i_data_bus[835]), .Z(N870) );
  CKAN2D1BWP30P140LVT U2283 ( .A1(n13), .A2(i_data_bus[505]), .Z(N540) );
  CKAN2D1BWP30P140LVT U2284 ( .A1(n11), .A2(i_data_bus[504]), .Z(N539) );
  CKAN2D1BWP30P140LVT U2285 ( .A1(n7), .A2(i_data_bus[503]), .Z(N538) );
  CKAN2D1BWP30P140LVT U2286 ( .A1(n12), .A2(i_data_bus[502]), .Z(N537) );
  CKAN2D1BWP30P140LVT U2287 ( .A1(n12), .A2(i_data_bus[501]), .Z(N536) );
  CKAN2D1BWP30P140LVT U2288 ( .A1(n11), .A2(i_data_bus[761]), .Z(N796) );
  CKAN2D1BWP30P140LVT U2289 ( .A1(n9), .A2(i_data_bus[363]), .Z(N398) );
  CKAN2D1BWP30P140LVT U2290 ( .A1(n13), .A2(i_data_bus[368]), .Z(N403) );
  CKAN2D1BWP30P140LVT U2291 ( .A1(n11), .A2(i_data_bus[369]), .Z(N404) );
  CKAN2D1BWP30P140LVT U2292 ( .A1(n7), .A2(i_data_bus[370]), .Z(N405) );
  CKAN2D1BWP30P140LVT U2293 ( .A1(n10), .A2(i_data_bus[371]), .Z(N406) );
  CKAN2D1BWP30P140LVT U2294 ( .A1(n8), .A2(i_data_bus[372]), .Z(N407) );
  CKAN2D1BWP30P140LVT U2295 ( .A1(n7), .A2(i_data_bus[380]), .Z(N415) );
  CKAN2D1BWP30P140LVT U2296 ( .A1(n10), .A2(i_data_bus[381]), .Z(N416) );
  CKAN2D1BWP30P140LVT U2297 ( .A1(n8), .A2(i_data_bus[382]), .Z(N417) );
  CKAN2D1BWP30P140LVT U2298 ( .A1(n9), .A2(i_data_bus[383]), .Z(N418) );
  CKAN2D1BWP30P140LVT U2299 ( .A1(n13), .A2(i_data_bus[384]), .Z(N419) );
  CKAN2D1BWP30P140LVT U2300 ( .A1(n14), .A2(i_data_bus[385]), .Z(N420) );
  CKAN2D1BWP30P140LVT U2301 ( .A1(n14), .A2(i_data_bus[386]), .Z(N421) );
  CKAN2D1BWP30P140LVT U2302 ( .A1(n14), .A2(i_data_bus[387]), .Z(N422) );
  CKAN2D1BWP30P140LVT U2303 ( .A1(n14), .A2(i_data_bus[388]), .Z(N423) );
  CKAN2D1BWP30P140LVT U2304 ( .A1(n8), .A2(i_data_bus[881]), .Z(N916) );
  CKAN2D1BWP30P140LVT U2305 ( .A1(n11), .A2(i_data_bus[880]), .Z(N915) );
  CKAN2D1BWP30P140LVT U2306 ( .A1(n14), .A2(i_data_bus[879]), .Z(N914) );
  CKAN2D1BWP30P140LVT U2307 ( .A1(n9), .A2(i_data_bus[878]), .Z(N913) );
  CKAN2D1BWP30P140LVT U2308 ( .A1(n7), .A2(i_data_bus[877]), .Z(N912) );
  CKAN2D1BWP30P140LVT U2309 ( .A1(n14), .A2(i_data_bus[389]), .Z(N424) );
  CKAN2D1BWP30P140LVT U2310 ( .A1(n14), .A2(i_data_bus[390]), .Z(N425) );
  CKAN2D1BWP30P140LVT U2311 ( .A1(n14), .A2(i_data_bus[391]), .Z(N426) );
  CKAN2D1BWP30P140LVT U2312 ( .A1(n7), .A2(i_data_bus[392]), .Z(N427) );
  CKAN2D1BWP30P140LVT U2313 ( .A1(n9), .A2(i_data_bus[428]), .Z(N463) );
  CKAN2D1BWP30P140LVT U2314 ( .A1(n13), .A2(i_data_bus[429]), .Z(N464) );
  CKAN2D1BWP30P140LVT U2315 ( .A1(n11), .A2(i_data_bus[430]), .Z(N465) );
  CKAN2D1BWP30P140LVT U2316 ( .A1(n7), .A2(i_data_bus[431]), .Z(N466) );
  CKAN2D1BWP30P140LVT U2317 ( .A1(n10), .A2(i_data_bus[432]), .Z(N467) );
  CKAN2D1BWP30P140LVT U2318 ( .A1(n8), .A2(i_data_bus[433]), .Z(N468) );
  CKAN2D1BWP30P140LVT U2319 ( .A1(n9), .A2(i_data_bus[434]), .Z(N469) );
  CKAN2D1BWP30P140LVT U2320 ( .A1(n13), .A2(i_data_bus[435]), .Z(N470) );
  CKAN2D1BWP30P140LVT U2321 ( .A1(n11), .A2(i_data_bus[440]), .Z(N475) );
  CKAN2D1BWP30P140LVT U2322 ( .A1(n7), .A2(i_data_bus[441]), .Z(N476) );
  CKAN2D1BWP30P140LVT U2323 ( .A1(n10), .A2(i_data_bus[442]), .Z(N477) );
  CKAN2D1BWP30P140LVT U2324 ( .A1(n8), .A2(i_data_bus[443]), .Z(N478) );
  CKAN2D1BWP30P140LVT U2325 ( .A1(n9), .A2(i_data_bus[444]), .Z(N479) );
  CKAN2D1BWP30P140LVT U2326 ( .A1(n7), .A2(i_data_bus[452]), .Z(N487) );
  CKAN2D1BWP30P140LVT U2327 ( .A1(n10), .A2(i_data_bus[453]), .Z(N488) );
  CKAN2D1BWP30P140LVT U2328 ( .A1(n13), .A2(i_data_bus[857]), .Z(N892) );
  CKAN2D1BWP30P140LVT U2329 ( .A1(n10), .A2(i_data_bus[856]), .Z(N891) );
  CKAN2D1BWP30P140LVT U2330 ( .A1(n14), .A2(i_data_bus[855]), .Z(N890) );
  CKAN2D1BWP30P140LVT U2331 ( .A1(n13), .A2(i_data_bus[854]), .Z(N889) );
  CKAN2D1BWP30P140LVT U2332 ( .A1(n12), .A2(i_cmd[67]), .Z(N1126) );
  CKAN2D1BWP30P140LVT U2333 ( .A1(n14), .A2(i_data_bus[852]), .Z(N887) );
  CKAN2D1BWP30P140LVT U2334 ( .A1(n8), .A2(i_data_bus[454]), .Z(N489) );
  CKAN2D1BWP30P140LVT U2335 ( .A1(n14), .A2(i_data_bus[463]), .Z(N498) );
  CKAN2D1BWP30P140LVT U2336 ( .A1(n9), .A2(i_data_bus[455]), .Z(N490) );
  CKAN2D1BWP30P140LVT U2337 ( .A1(n13), .A2(i_data_bus[456]), .Z(N491) );
  CKAN2D1BWP30P140LVT U2338 ( .A1(n14), .A2(i_data_bus[458]), .Z(N493) );
  CKAN2D1BWP30P140LVT U2339 ( .A1(n11), .A2(i_data_bus[464]), .Z(N499) );
  CKAN2D1BWP30P140LVT U2340 ( .A1(n12), .A2(i_data_bus[853]), .Z(N888) );
  CKAN2D1BWP30P140LVT U2341 ( .A1(n14), .A2(i_data_bus[459]), .Z(N494) );
  CKAN2D1BWP30P140LVT U2342 ( .A1(n14), .A2(i_data_bus[460]), .Z(N495) );
  CKAN2D1BWP30P140LVT U2343 ( .A1(n14), .A2(i_data_bus[461]), .Z(N496) );
  CKAN2D1BWP30P140LVT U2344 ( .A1(n14), .A2(i_data_bus[462]), .Z(N497) );
  CKAN2D1BWP30P140LVT U2345 ( .A1(n10), .A2(i_data_bus[500]), .Z(N535) );
  CKAN2D1BWP30P140LVT U2346 ( .A1(n14), .A2(i_data_bus[212]), .Z(N247) );
  CKAN2D1BWP30P140LVT U2347 ( .A1(n14), .A2(i_data_bus[213]), .Z(N248) );
  CKAN2D1BWP30P140LVT U2348 ( .A1(n14), .A2(i_data_bus[214]), .Z(N249) );
  CKAN2D1BWP30P140LVT U2349 ( .A1(n12), .A2(i_data_bus[215]), .Z(N250) );
  CKAN2D1BWP30P140LVT U2350 ( .A1(n14), .A2(i_data_bus[216]), .Z(N251) );
  CKAN2D1BWP30P140LVT U2351 ( .A1(n14), .A2(i_data_bus[217]), .Z(N252) );
  CKAN2D1BWP30P140LVT U2352 ( .A1(n7), .A2(i_data_bus[218]), .Z(N253) );
  CKAN2D1BWP30P140LVT U2353 ( .A1(n7), .A2(i_data_bus[219]), .Z(N254) );
  CKAN2D1BWP30P140LVT U2354 ( .A1(n8), .A2(i_data_bus[224]), .Z(N259) );
  CKAN2D1BWP30P140LVT U2355 ( .A1(n11), .A2(i_data_bus[225]), .Z(N260) );
  CKAN2D1BWP30P140LVT U2356 ( .A1(n13), .A2(i_data_bus[226]), .Z(N261) );
  CKAN2D1BWP30P140LVT U2357 ( .A1(n10), .A2(i_data_bus[227]), .Z(N262) );
  CKAN2D1BWP30P140LVT U2358 ( .A1(n14), .A2(i_data_bus[228]), .Z(N263) );
  CKAN2D1BWP30P140LVT U2359 ( .A1(n13), .A2(i_data_bus[284]), .Z(N319) );
  CKAN2D1BWP30P140LVT U2360 ( .A1(n13), .A2(i_data_bus[285]), .Z(N320) );
  CKAN2D1BWP30P140LVT U2361 ( .A1(n13), .A2(i_data_bus[286]), .Z(N321) );
  CKAN2D1BWP30P140LVT U2362 ( .A1(n13), .A2(i_data_bus[287]), .Z(N322) );
  CKAN2D1BWP30P140LVT U2363 ( .A1(n13), .A2(i_data_bus[288]), .Z(N323) );
  CKAN2D1BWP30P140LVT U2364 ( .A1(n13), .A2(i_data_bus[289]), .Z(N324) );
  CKAN2D1BWP30P140LVT U2365 ( .A1(n13), .A2(i_data_bus[290]), .Z(N325) );
  CKAN2D1BWP30P140LVT U2366 ( .A1(n13), .A2(i_data_bus[291]), .Z(N326) );
  CKAN2D1BWP30P140LVT U2367 ( .A1(n13), .A2(i_data_bus[296]), .Z(N331) );
  CKAN2D1BWP30P140LVT U2368 ( .A1(n13), .A2(i_data_bus[297]), .Z(N332) );
  CKAN2D1BWP30P140LVT U2369 ( .A1(n13), .A2(i_data_bus[298]), .Z(N333) );
  CKAN2D1BWP30P140LVT U2370 ( .A1(n13), .A2(i_data_bus[299]), .Z(N334) );
  CKAN2D1BWP30P140LVT U2371 ( .A1(n13), .A2(i_data_bus[300]), .Z(N335) );
  CKAN2D1BWP30P140LVT U2372 ( .A1(n13), .A2(i_data_bus[602]), .Z(N637) );
  CKAN2D1BWP30P140LVT U2373 ( .A1(n13), .A2(i_data_bus[603]), .Z(N638) );
  CKAN2D1BWP30P140LVT U2374 ( .A1(n14), .A2(i_data_bus[604]), .Z(N639) );
  CKAN2D1BWP30P140LVT U2375 ( .A1(n13), .A2(i_data_bus[605]), .Z(N640) );
  CKAN2D1BWP30P140LVT U2376 ( .A1(n10), .A2(i_data_bus[606]), .Z(N641) );
  CKAN2D1BWP30P140LVT U2377 ( .A1(n13), .A2(i_data_bus[607]), .Z(N642) );
  CKAN2D1BWP30P140LVT U2378 ( .A1(n7), .A2(i_data_bus[644]), .Z(N679) );
  CKAN2D1BWP30P140LVT U2379 ( .A1(n8), .A2(i_data_bus[645]), .Z(N680) );
  CKAN2D1BWP30P140LVT U2380 ( .A1(n9), .A2(i_data_bus[646]), .Z(N681) );
  CKAN2D1BWP30P140LVT U2381 ( .A1(n12), .A2(i_data_bus[647]), .Z(N682) );
  CKAN2D1BWP30P140LVT U2382 ( .A1(n12), .A2(i_data_bus[648]), .Z(N683) );
  CKAN2D1BWP30P140LVT U2383 ( .A1(n8), .A2(i_data_bus[649]), .Z(N684) );
  CKAN2D1BWP30P140LVT U2384 ( .A1(n9), .A2(i_data_bus[650]), .Z(N685) );
  CKAN2D1BWP30P140LVT U2385 ( .A1(n12), .A2(i_data_bus[651]), .Z(N686) );
  CKAN2D1BWP30P140LVT U2386 ( .A1(n13), .A2(i_data_bus[656]), .Z(N691) );
  CKAN2D1BWP30P140LVT U2387 ( .A1(n14), .A2(i_data_bus[657]), .Z(N692) );
  CKAN2D1BWP30P140LVT U2388 ( .A1(n11), .A2(i_data_bus[658]), .Z(N693) );
  CKAN2D1BWP30P140LVT U2389 ( .A1(n8), .A2(i_data_bus[659]), .Z(N694) );
  CKAN2D1BWP30P140LVT U2390 ( .A1(n9), .A2(i_data_bus[660]), .Z(N695) );
  CKAN2D1BWP30P140LVT U2391 ( .A1(n8), .A2(i_data_bus[668]), .Z(N703) );
  CKAN2D1BWP30P140LVT U2392 ( .A1(n9), .A2(i_data_bus[669]), .Z(N704) );
  CKAN2D1BWP30P140LVT U2393 ( .A1(n13), .A2(i_data_bus[670]), .Z(N705) );
  CKAN2D1BWP30P140LVT U2394 ( .A1(n7), .A2(i_data_bus[671]), .Z(N706) );
  CKAN2D1BWP30P140LVT U2395 ( .A1(n7), .A2(i_data_bus[672]), .Z(N707) );
  CKAN2D1BWP30P140LVT U2396 ( .A1(n9), .A2(i_data_bus[680]), .Z(N715) );
  CKAN2D1BWP30P140LVT U2397 ( .A1(n10), .A2(i_data_bus[716]), .Z(N751) );
  CKAN2D1BWP30P140LVT U2398 ( .A1(n10), .A2(i_data_bus[717]), .Z(N752) );
  CKAN2D1BWP30P140LVT U2399 ( .A1(n8), .A2(i_data_bus[718]), .Z(N753) );
  CKAN2D1BWP30P140LVT U2400 ( .A1(n9), .A2(i_data_bus[719]), .Z(N754) );
  CKAN2D1BWP30P140LVT U2401 ( .A1(n12), .A2(i_data_bus[720]), .Z(N755) );
  CKAN2D1BWP30P140LVT U2402 ( .A1(n10), .A2(i_data_bus[721]), .Z(N756) );
  CKAN2D1BWP30P140LVT U2403 ( .A1(n11), .A2(i_data_bus[722]), .Z(N757) );
  CKAN2D1BWP30P140LVT U2404 ( .A1(n8), .A2(i_data_bus[723]), .Z(N758) );
  CKAN2D1BWP30P140LVT U2405 ( .A1(n9), .A2(i_data_bus[728]), .Z(N763) );
  CKAN2D1BWP30P140LVT U2406 ( .A1(n12), .A2(i_data_bus[729]), .Z(N764) );
  CKAN2D1BWP30P140LVT U2407 ( .A1(n13), .A2(i_data_bus[730]), .Z(N765) );
  CKAN2D1BWP30P140LVT U2408 ( .A1(n12), .A2(i_data_bus[731]), .Z(N766) );
  CKAN2D1BWP30P140LVT U2409 ( .A1(n10), .A2(i_data_bus[732]), .Z(N767) );
  CKAN2D1BWP30P140LVT U2410 ( .A1(n14), .A2(i_data_bus[884]), .Z(N919) );
  CKAN2D1BWP30P140LVT U2411 ( .A1(n14), .A2(i_data_bus[885]), .Z(N920) );
  CKAN2D1BWP30P140LVT U2412 ( .A1(n14), .A2(i_data_bus[886]), .Z(N921) );
  CKAN2D1BWP30P140LVT U2413 ( .A1(n14), .A2(i_data_bus[887]), .Z(N922) );
  CKAN2D1BWP30P140LVT U2414 ( .A1(n14), .A2(i_data_bus[888]), .Z(N923) );
  CKAN2D1BWP30P140LVT U2415 ( .A1(n14), .A2(i_data_bus[896]), .Z(N931) );
  CKAN2D1BWP30P140LVT U2416 ( .A1(n10), .A2(i_data_bus[932]), .Z(N967) );
  CKAN2D1BWP30P140LVT U2417 ( .A1(n13), .A2(i_data_bus[933]), .Z(N968) );
  CKAN2D1BWP30P140LVT U2418 ( .A1(n9), .A2(i_data_bus[934]), .Z(N969) );
  CKAN2D1BWP30P140LVT U2419 ( .A1(n13), .A2(i_data_bus[935]), .Z(N970) );
  CKAN2D1BWP30P140LVT U2420 ( .A1(n11), .A2(i_data_bus[936]), .Z(N971) );
  CKAN2D1BWP30P140LVT U2421 ( .A1(n13), .A2(i_data_bus[937]), .Z(N972) );
  CKAN2D1BWP30P140LVT U2422 ( .A1(n13), .A2(i_data_bus[938]), .Z(N973) );
  CKAN2D1BWP30P140LVT U2423 ( .A1(n13), .A2(i_data_bus[939]), .Z(N974) );
  CKAN2D1BWP30P140LVT U2424 ( .A1(n14), .A2(i_data_bus[944]), .Z(N979) );
  CKAN2D1BWP30P140LVT U2425 ( .A1(n13), .A2(i_data_bus[945]), .Z(N980) );
  CKAN2D1BWP30P140LVT U2426 ( .A1(n14), .A2(i_data_bus[946]), .Z(N981) );
  CKAN2D1BWP30P140LVT U2427 ( .A1(n13), .A2(i_data_bus[947]), .Z(N982) );
  CKAN2D1BWP30P140LVT U2428 ( .A1(n12), .A2(i_data_bus[948]), .Z(N983) );
  CKAN2D1BWP30P140LVT U2429 ( .A1(n14), .A2(i_data_bus[966]), .Z(N1001) );
  CKAN2D1BWP30P140LVT U2430 ( .A1(n14), .A2(i_data_bus[967]), .Z(N1002) );
  CKAN2D1BWP30P140LVT U2431 ( .A1(n12), .A2(i_data_bus[1004]), .Z(N1039) );
  CKAN2D1BWP30P140LVT U2432 ( .A1(n13), .A2(i_data_bus[1005]), .Z(N1040) );
  CKAN2D1BWP30P140LVT U2433 ( .A1(n14), .A2(i_data_bus[1006]), .Z(N1041) );
  CKAN2D1BWP30P140LVT U2434 ( .A1(n7), .A2(i_data_bus[1007]), .Z(N1042) );
  CKAN2D1BWP30P140LVT U2435 ( .A1(n12), .A2(i_data_bus[1008]), .Z(N1043) );
  CKAN2D1BWP30P140LVT U2436 ( .A1(n7), .A2(i_data_bus[1009]), .Z(N1044) );
  CKAN2D1BWP30P140LVT U2437 ( .A1(n12), .A2(i_data_bus[1010]), .Z(N1045) );
  CKAN2D1BWP30P140LVT U2438 ( .A1(n7), .A2(i_data_bus[1011]), .Z(N1046) );
  CKAN2D1BWP30P140LVT U2439 ( .A1(n13), .A2(i_data_bus[1016]), .Z(N1051) );
  CKAN2D1BWP30P140LVT U2440 ( .A1(n7), .A2(i_data_bus[1017]), .Z(N1052) );
  CKAN2D1BWP30P140LVT U2441 ( .A1(n14), .A2(i_data_bus[1018]), .Z(N1053) );
  CKAN2D1BWP30P140LVT U2442 ( .A1(n11), .A2(i_data_bus[1019]), .Z(N1054) );
  CKAN2D1BWP30P140LVT U2443 ( .A1(n11), .A2(i_data_bus[1020]), .Z(N1055) );
endmodule

