`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module local_controller_prefetch_full(CLK, reset, init,  from_glob_controller_delay,  input_boundary_flag, prev_dest_address, from_glob_dest_addr, packet_out, boundary_next, dest_address, from_glob_controller_valid, ext_CEB, WEB, WEBM, D, BWEB, DM, BWEBM, ext_sample_address, ext_sample_address_M, write_flag, from_glob_prefetch_valid, from_glob_prefetch_start, from_glob_prefetch_stop, from_glob_prefetch_dest, prefetch_packet_out);

    // parameter
    	parameter N_sample = 256;
	parameter datawidth = 16;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 4; // 16 local controllers in subscaled system
	parameter sample_address_width = 8; /// assuming 1024 rows and 64 columns: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	

//=== IO Ports ===//

     // Normal Mode Input
        input WEB;
        input [31:0] D;
        input [31:0] BWEB;

     // BIST Mode Input
        input WEBM;
        input [31:0] DM;
        input [31:0] BWEBM;

    // input
    	input CLK; // system clock, generated by VCO
	input reset;
	input init;	
	input from_glob_controller_valid;
	input input_boundary_flag;
	input [address_vector_width - 1:0] prev_dest_address;
	input [address_vector_width - 1:0] from_glob_dest_addr;
	input [address_vector_width - 1:0] from_glob_prefetch_dest;
	input [sample_address_width - 1:0] from_glob_controller_delay;
        input [sample_address_width-1:0] ext_sample_address;	
        input [sample_address_width-1:0] ext_sample_address_M;
	input write_flag;
	input ext_CEB;
	input from_glob_prefetch_valid;
	input [sample_address_width - 1:0] from_glob_prefetch_start;
	input [sample_address_width - 1:0] from_glob_prefetch_stop;

    // output
        output reg [packet_width-1:0] packet_out;  
        output reg [packet_width-1:0] prefetch_packet_out;  
        output reg boundary_next;
        output reg [address_vector_width - 1:0] dest_address;

//////////// internal status regs/signals //////////////////////////////////
    //reg [packet_width-1:0] packet_out_internal;
    reg coeff_num;
    reg [sample_address_width - 1:0] delay;
    wire [2*datawidth - 1:0] data_from_sram;
    reg [2*datawidth - 1:0] packet_out_data;
    reg [sample_address_width-1:0] sample_address;	
    reg [sample_address_width-1:0] sample_address_M;
    reg [sample_address_width-1:0] prefetch_sample_address;
    reg prefetch_reqd;
    reg [address_vector_width - 1:0] prefetch_dest_addr;
    reg [sample_address_width - 1:0] prefetch_stop_address;



    reg BIST;
    reg AWT;
    reg SLP;
    reg SD;
    reg CEB;
    reg prefetch_CEB;
    reg CEBM;
    wire [sample_address_width-1:0] A;	
    wire [sample_address_width-1:0] AM;
    wire sram_CEB;
    wire CLK_n;


///////////////////////////////////////////////////////////////////////////////    

////////// logic part ///////////////////////////////////////////////////////  


    //assign packet_out = packet_out_internal;
    //assign CLK_n = ~CLK;
    assign A = write_flag ? ext_sample_address : (coeff_num ? sample_address: prefetch_sample_address);
    assign AM = write_flag ? ext_sample_address_M : sample_address_M;
    assign sram_CEB = write_flag ? ext_CEB : (CEB & prefetch_CEB);


////////////sequential logic
    always @ (posedge CLK_n) begin
        if (reset) begin

			sample_address <= 8'b0;
			sample_address_M <= 0;
			packet_out <= 40'bz;
			dest_address <= 0;
			coeff_num <= 0;
			delay <= 0;
			boundary_next <= 0;
			BIST <= 0;
			AWT <= 0;
			SLP <= 0;
			SD <= 0;
			CEB <= 1;
			CEBM <= 1;
			
        end
        else if (from_glob_controller_valid == 1) begin
			packet_out <= 40'bz;
			boundary_next <=0;
			sample_address <= from_glob_controller_delay;
			dest_address <= from_glob_dest_addr;
			coeff_num <= 1;
			delay <= from_glob_controller_delay;
			
			sample_address_M <= 0;

                        BIST <= 0;
			AWT <= 0;
			SLP <= 0;
			SD <= 0;
			CEB <= 1;
			CEBM <= 1;

	end
			

	else begin
			if (coeff_num == 1 && input_boundary_flag == 0 && boundary_next == 0) begin		// && write_flag == 0) begin
				packet_out <= {packet_out_data, dest_address};
				sample_address <= sample_address + 1;
				CEB <= 0;
				CEBM <= 1;
				dest_address <= dest_address;
				coeff_num <= coeff_num;
				if (sample_address == N_sample - 2) begin
					boundary_next <= 1;

				end
				else begin
					boundary_next <= 0;

				end

			end
			else if (coeff_num == 1 && input_boundary_flag == 0 && boundary_next == 1) begin		// && write_flag == 0) begin
				packet_out <= {packet_out_data, dest_address};
				sample_address <= sample_address + 1;   /// should automatically go to 0th address
				CEB <= 1;
				CEBM <= 1;
				dest_address <= dest_address;
				coeff_num <= 0;
				boundary_next <= 0;

			end

			else if (coeff_num == 0 && input_boundary_flag == 1 && boundary_next == 0) begin		// && write_flag == 0) begin
				packet_out <= 40'bz;
				sample_address <= 8'b0;   /// should automatically go to 0th address
				CEB <= 0;
				CEBM <= 1;
				dest_address <= prev_dest_address;
				coeff_num <= 1;
				boundary_next <= boundary_next;

			end

			else if (coeff_num == 0 && input_boundary_flag == 1 && boundary_next == 1) begin		// && write_flag == 0) begin
				packet_out <= 40'bz;
				sample_address <= 8'b0;   /// should automatically go to 0th address
				CEB <= 0;
				CEBM <= 1;
				dest_address <= prev_dest_address;
				coeff_num <= 1;
				boundary_next <= 0;

			end


			else begin
				packet_out <= 40'bz;
				sample_address <= sample_address;
				dest_address <= dest_address;
				coeff_num <= coeff_num;
				boundary_next <= boundary_next;
				CEB <= 1;
				CEBM <= 1;

			end

			delay <= delay;
			sample_address_M <= 0;
                        BIST <= 0;
			AWT <= 0;
			SLP <= 0;
			SD <= 0;

	end  
     end

     always @(posedge CLK_n) begin   //// merge with prev always block: prefetch sample address is assigned in both
        if (reset) begin
			prefetch_sample_address <= 8'b0;
			prefetch_packet_out <= 40'bz;
			prefetch_reqd <= 0;
			prefetch_dest_addr <= 0;
			prefetch_stop_address <= 0;
			prefetch_CEB <= 1;		
        end
        else if (init) begin

			prefetch_sample_address <= 8'b0;
			prefetch_packet_out <= 40'bz;
			prefetch_reqd <= 0;
			prefetch_dest_addr <= 0;
			prefetch_stop_address <= 0;
			prefetch_CEB <= 1;
        end
	else if (from_glob_prefetch_valid == 1) begin
		prefetch_dest_addr <= from_glob_prefetch_dest;
		prefetch_reqd <= 1;
		prefetch_sample_address <= from_glob_prefetch_start;
		prefetch_packet_out <= 40'bz;
		prefetch_stop_address <= from_glob_prefetch_stop;
		prefetch_CEB <= 1;
	end
	else if (coeff_num == 0 && input_boundary_flag == 0 && prefetch_reqd == 1)  begin
		prefetch_dest_addr <= prefetch_dest_addr;
		prefetch_stop_address <= prefetch_stop_address;
		prefetch_packet_out <= {packet_out_data,prefetch_dest_addr};
		prefetch_sample_address <= prefetch_sample_address + 1;
		if (prefetch_sample_address == prefetch_stop_address) begin
			prefetch_reqd <= 0;
			prefetch_CEB <= 1;
		end	
		else begin
			prefetch_reqd <= prefetch_reqd;
			prefetch_CEB <= 0;
		end		

	end
	else begin
		prefetch_dest_addr <= prefetch_dest_addr;
		prefetch_reqd <= prefetch_reqd;
		prefetch_stop_address <= prefetch_stop_address;
		prefetch_sample_address <= prefetch_sample_address;
		prefetch_packet_out <= 40'bz;
		prefetch_CEB <= prefetch_CEB;
	end


     end


     always @(posedge CLK) begin
	packet_out_data <= data_from_sram;

     end


    INVD6BWP30P140 UI_342 ( .I(CLK), .ZN(CLK_n) );

    TS1N28HPCPLVTB256X32M4SWBASO UI_dut_mem (.SLP(SLP), .SD(SD), .CLK(CLK), .CEB(sram_CEB), .WEB(WEB), .CEBM(CEBM), .WEBM(WEBM), .AWT(AWT), .A(A), .D(D), .BWEB(BWEB), .AM(AM), .DM(DM), .BWEBM(BWEBM), .BIST(BIST), .Q(data_from_sram));

	 
	 


   
endmodule
    
