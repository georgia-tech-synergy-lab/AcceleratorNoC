
module linear_network_unicast_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [31:0] i_data_bus;
  output [15:0] o_valid;
  output [511:0] o_data_bus;
  input [3:0] i_cmd;
  input clk, rst, i_valid, i_en;
  wire   N183, N184, N185, N186, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N320, N321, N322, N390, N391, N392, N393, N394,
         N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
         N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416,
         N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427,
         N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N457, N458, N526, N527, N528,
         N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539,
         N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550,
         N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561,
         N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572,
         N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583,
         N584, N585, N586, N587, N588, N589, N590, N591, N593, N594, N662,
         N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673,
         N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684,
         N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695,
         N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706,
         N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717,
         N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728,
         N730, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807,
         N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818,
         N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829,
         N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840,
         N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851,
         N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862,
         N864, N865, N866, N934, N935, N936, N937, N938, N939, N940, N941,
         N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952,
         N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963,
         N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974,
         N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985,
         N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996,
         N997, N998, N999, N1001, N1002, N1070, N1071, N1072, N1073, N1074,
         N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084,
         N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094,
         N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104,
         N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114,
         N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124,
         N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134,
         N1135, N1136, N1138, N1206, N1207, N1208, N1209, N1210, N1211, N1212,
         N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222,
         N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232,
         N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242,
         N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252,
         N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262,
         N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272,
         N1273, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350,
         N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360,
         N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370,
         N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380,
         N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390,
         N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400,
         N1401, N1402, N1403, N1404, N1405, N1406, N1408, N1409, N1410, N1478,
         N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488,
         N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498,
         N1499, N1500, N1501, N1502, N1503, N1504, N1505, N1506, N1507, N1508,
         N1509, N1510, N1511, N1512, N1513, N1514, N1515, N1516, N1517, N1518,
         N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528,
         N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538,
         N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1614, N1615, N1616,
         N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626,
         N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636,
         N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646,
         N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656,
         N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664, N1665, N1666,
         N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674, N1675, N1676,
         N1677, N1678, N1679, N1681, N1682, N1750, N1751, N1752, N1753, N1754,
         N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764,
         N1765, N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774,
         N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784,
         N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794,
         N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804,
         N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814,
         N1815, N1816, N1817, N1886, N1887, N1888, N1889, N1890, N1891, N1892,
         N1893, N1894, N1895, N1896, N1897, N1898, N1899, N1900, N1901, N1902,
         N1903, N1904, N1905, N1906, N1907, N1908, N1909, N1910, N1911, N1912,
         N1913, N1914, N1915, N1916, N1917, N1918, N1919, N1920, N1921, N1922,
         N1923, N1924, N1925, N1926, N1927, N1928, N1929, N1930, N1931, N1932,
         N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942,
         N1943, N1944, N1945, N1946, N1947, N1948, N1949, N1950, N1951, N1952,
         N1953, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030,
         N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2039, N2040,
         N2041, N2042, N2043, N2044, N2045, N2046, N2047, N2048, N2049, N2050,
         N2051, N2052, N2053, N2054, N2055, N2056, N2057, N2058, N2059, N2060,
         N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069, N2070,
         N2071, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079, N2080,
         N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2090, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304;
  wire   [479:0] o_data_forward_reg;
  wire   [0:14] o_valid_forward_reg;
  wire   [59:0] o_cmd_forward_reg;

  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__3_ ( .D(N186), .CP(clk), .Q(
        o_cmd_forward_reg[59]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__2_ ( .D(N185), .CP(clk), .Q(
        o_cmd_forward_reg[58]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__1_ ( .D(N184), .CP(clk), .Q(
        o_cmd_forward_reg[57]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__0_ ( .D(N183), .CP(clk), .Q(
        o_cmd_forward_reg[56]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__31_ ( .D(n209), .CP(clk), .Q(
        o_data_forward_reg[479]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__30_ ( .D(n208), .CP(clk), .Q(
        o_data_forward_reg[478]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__29_ ( .D(n207), .CP(clk), .Q(
        o_data_forward_reg[477]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__28_ ( .D(n206), .CP(clk), .Q(
        o_data_forward_reg[476]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__27_ ( .D(n205), .CP(clk), .Q(
        o_data_forward_reg[475]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__26_ ( .D(n204), .CP(clk), .Q(
        o_data_forward_reg[474]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__25_ ( .D(n203), .CP(clk), .Q(
        o_data_forward_reg[473]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__24_ ( .D(n202), .CP(clk), .Q(
        o_data_forward_reg[472]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__23_ ( .D(n201), .CP(clk), .Q(
        o_data_forward_reg[471]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__22_ ( .D(n200), .CP(clk), .Q(
        o_data_forward_reg[470]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__21_ ( .D(n199), .CP(clk), .Q(
        o_data_forward_reg[469]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__20_ ( .D(n198), .CP(clk), .Q(
        o_data_forward_reg[468]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__19_ ( .D(n197), .CP(clk), .Q(
        o_data_forward_reg[467]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__18_ ( .D(n196), .CP(clk), .Q(
        o_data_forward_reg[466]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__17_ ( .D(n195), .CP(clk), .Q(
        o_data_forward_reg[465]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__16_ ( .D(n194), .CP(clk), .Q(
        o_data_forward_reg[464]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__15_ ( .D(n193), .CP(clk), .Q(
        o_data_forward_reg[463]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__14_ ( .D(n192), .CP(clk), .Q(
        o_data_forward_reg[462]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__13_ ( .D(n191), .CP(clk), .Q(
        o_data_forward_reg[461]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__12_ ( .D(n190), .CP(clk), .Q(
        o_data_forward_reg[460]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__11_ ( .D(n189), .CP(clk), .Q(
        o_data_forward_reg[459]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__10_ ( .D(n188), .CP(clk), .Q(
        o_data_forward_reg[458]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__9_ ( .D(n187), .CP(clk), .Q(
        o_data_forward_reg[457]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__8_ ( .D(n186), .CP(clk), .Q(
        o_data_forward_reg[456]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__7_ ( .D(n185), .CP(clk), .Q(
        o_data_forward_reg[455]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__6_ ( .D(n184), .CP(clk), .Q(
        o_data_forward_reg[454]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__5_ ( .D(n183), .CP(clk), .Q(
        o_data_forward_reg[453]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__4_ ( .D(n182), .CP(clk), .Q(
        o_data_forward_reg[452]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__3_ ( .D(n181), .CP(clk), .Q(
        o_data_forward_reg[451]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__2_ ( .D(n180), .CP(clk), .Q(
        o_data_forward_reg[450]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__1_ ( .D(n179), .CP(clk), .Q(
        o_data_forward_reg[449]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__0_ ( .D(n178), .CP(clk), .Q(
        o_data_forward_reg[448]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_0_ ( .D(n295), .CP(clk), .Q(
        o_valid_forward_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__3_ ( .D(N322), .CP(clk), .Q(
        o_cmd_forward_reg[55]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__2_ ( .D(N321), .CP(clk), .Q(
        o_cmd_forward_reg[54]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__1_ ( .D(N320), .CP(clk), .Q(
        o_cmd_forward_reg[53]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__0_ ( .D(n296), .CP(clk), .Q(
        o_cmd_forward_reg[52]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__31_ ( .D(N317), .CP(clk), .Q(
        o_data_forward_reg[447]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__30_ ( .D(N316), .CP(clk), .Q(
        o_data_forward_reg[446]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__29_ ( .D(N315), .CP(clk), .Q(
        o_data_forward_reg[445]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__28_ ( .D(N314), .CP(clk), .Q(
        o_data_forward_reg[444]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__27_ ( .D(N313), .CP(clk), .Q(
        o_data_forward_reg[443]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__26_ ( .D(N312), .CP(clk), .Q(
        o_data_forward_reg[442]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__25_ ( .D(N311), .CP(clk), .Q(
        o_data_forward_reg[441]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__24_ ( .D(N310), .CP(clk), .Q(
        o_data_forward_reg[440]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__23_ ( .D(N309), .CP(clk), .Q(
        o_data_forward_reg[439]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__22_ ( .D(N308), .CP(clk), .Q(
        o_data_forward_reg[438]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__21_ ( .D(N307), .CP(clk), .Q(
        o_data_forward_reg[437]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__20_ ( .D(N306), .CP(clk), .Q(
        o_data_forward_reg[436]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__19_ ( .D(N305), .CP(clk), .Q(
        o_data_forward_reg[435]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__18_ ( .D(N304), .CP(clk), .Q(
        o_data_forward_reg[434]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__17_ ( .D(N303), .CP(clk), .Q(
        o_data_forward_reg[433]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__16_ ( .D(N302), .CP(clk), .Q(
        o_data_forward_reg[432]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__15_ ( .D(N301), .CP(clk), .Q(
        o_data_forward_reg[431]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__14_ ( .D(N300), .CP(clk), .Q(
        o_data_forward_reg[430]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__13_ ( .D(N299), .CP(clk), .Q(
        o_data_forward_reg[429]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__12_ ( .D(N298), .CP(clk), .Q(
        o_data_forward_reg[428]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__11_ ( .D(N297), .CP(clk), .Q(
        o_data_forward_reg[427]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__10_ ( .D(N296), .CP(clk), .Q(
        o_data_forward_reg[426]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__9_ ( .D(N295), .CP(clk), .Q(
        o_data_forward_reg[425]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__8_ ( .D(N294), .CP(clk), .Q(
        o_data_forward_reg[424]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__7_ ( .D(N293), .CP(clk), .Q(
        o_data_forward_reg[423]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__6_ ( .D(N292), .CP(clk), .Q(
        o_data_forward_reg[422]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__5_ ( .D(N291), .CP(clk), .Q(
        o_data_forward_reg[421]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__4_ ( .D(N290), .CP(clk), .Q(
        o_data_forward_reg[420]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__3_ ( .D(N289), .CP(clk), .Q(
        o_data_forward_reg[419]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__2_ ( .D(N288), .CP(clk), .Q(
        o_data_forward_reg[418]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__1_ ( .D(N287), .CP(clk), .Q(
        o_data_forward_reg[417]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__0_ ( .D(N286), .CP(clk), .Q(
        o_data_forward_reg[416]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_1_ ( .D(N318), .CP(clk), .Q(
        o_valid_forward_reg[1]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__3_ ( .D(N458), .CP(clk), .Q(
        o_cmd_forward_reg[51]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__2_ ( .D(N457), .CP(clk), .Q(
        o_cmd_forward_reg[50]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__1_ ( .D(n293), .CP(clk), .Q(
        o_cmd_forward_reg[49]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__0_ ( .D(N455), .CP(clk), .Q(
        o_cmd_forward_reg[48]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__31_ ( .D(N453), .CP(clk), .Q(
        o_data_forward_reg[415]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__30_ ( .D(N452), .CP(clk), .Q(
        o_data_forward_reg[414]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__29_ ( .D(N451), .CP(clk), .Q(
        o_data_forward_reg[413]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__28_ ( .D(N450), .CP(clk), .Q(
        o_data_forward_reg[412]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__27_ ( .D(N449), .CP(clk), .Q(
        o_data_forward_reg[411]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__26_ ( .D(N448), .CP(clk), .Q(
        o_data_forward_reg[410]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__25_ ( .D(N447), .CP(clk), .Q(
        o_data_forward_reg[409]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__24_ ( .D(N446), .CP(clk), .Q(
        o_data_forward_reg[408]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__23_ ( .D(N445), .CP(clk), .Q(
        o_data_forward_reg[407]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__22_ ( .D(N444), .CP(clk), .Q(
        o_data_forward_reg[406]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__21_ ( .D(N443), .CP(clk), .Q(
        o_data_forward_reg[405]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__20_ ( .D(N442), .CP(clk), .Q(
        o_data_forward_reg[404]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__19_ ( .D(N441), .CP(clk), .Q(
        o_data_forward_reg[403]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__18_ ( .D(N440), .CP(clk), .Q(
        o_data_forward_reg[402]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__17_ ( .D(N439), .CP(clk), .Q(
        o_data_forward_reg[401]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__16_ ( .D(N438), .CP(clk), .Q(
        o_data_forward_reg[400]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__15_ ( .D(N437), .CP(clk), .Q(
        o_data_forward_reg[399]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__14_ ( .D(N436), .CP(clk), .Q(
        o_data_forward_reg[398]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__13_ ( .D(N435), .CP(clk), .Q(
        o_data_forward_reg[397]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__12_ ( .D(N434), .CP(clk), .Q(
        o_data_forward_reg[396]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__11_ ( .D(N433), .CP(clk), .Q(
        o_data_forward_reg[395]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__10_ ( .D(N432), .CP(clk), .Q(
        o_data_forward_reg[394]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__9_ ( .D(N431), .CP(clk), .Q(
        o_data_forward_reg[393]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__8_ ( .D(N430), .CP(clk), .Q(
        o_data_forward_reg[392]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__7_ ( .D(N429), .CP(clk), .Q(
        o_data_forward_reg[391]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__6_ ( .D(N428), .CP(clk), .Q(
        o_data_forward_reg[390]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__5_ ( .D(N427), .CP(clk), .Q(
        o_data_forward_reg[389]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__4_ ( .D(N426), .CP(clk), .Q(
        o_data_forward_reg[388]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__3_ ( .D(N425), .CP(clk), .Q(
        o_data_forward_reg[387]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__2_ ( .D(N424), .CP(clk), .Q(
        o_data_forward_reg[386]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__1_ ( .D(N423), .CP(clk), .Q(
        o_data_forward_reg[385]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__0_ ( .D(N422), .CP(clk), .Q(
        o_data_forward_reg[384]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_2_ ( .D(N454), .CP(clk), .Q(
        o_valid_forward_reg[2]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_3__3_ ( .D(N594), .CP(clk), .Q(
        o_cmd_forward_reg[47]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_3__2_ ( .D(N593), .CP(clk), .Q(
        o_cmd_forward_reg[46]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_3__1_ ( .D(n297), .CP(clk), .Q(
        o_cmd_forward_reg[45]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_3__0_ ( .D(N591), .CP(clk), .Q(
        o_cmd_forward_reg[44]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__31_ ( .D(N589), .CP(clk), .Q(
        o_data_forward_reg[383]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__30_ ( .D(N588), .CP(clk), .Q(
        o_data_forward_reg[382]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__29_ ( .D(N587), .CP(clk), .Q(
        o_data_forward_reg[381]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__28_ ( .D(N586), .CP(clk), .Q(
        o_data_forward_reg[380]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__27_ ( .D(N585), .CP(clk), .Q(
        o_data_forward_reg[379]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__26_ ( .D(N584), .CP(clk), .Q(
        o_data_forward_reg[378]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__25_ ( .D(N583), .CP(clk), .Q(
        o_data_forward_reg[377]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__24_ ( .D(N582), .CP(clk), .Q(
        o_data_forward_reg[376]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__23_ ( .D(N581), .CP(clk), .Q(
        o_data_forward_reg[375]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__22_ ( .D(N580), .CP(clk), .Q(
        o_data_forward_reg[374]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__21_ ( .D(N579), .CP(clk), .Q(
        o_data_forward_reg[373]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__20_ ( .D(N578), .CP(clk), .Q(
        o_data_forward_reg[372]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__19_ ( .D(N577), .CP(clk), .Q(
        o_data_forward_reg[371]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__18_ ( .D(N576), .CP(clk), .Q(
        o_data_forward_reg[370]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__17_ ( .D(N575), .CP(clk), .Q(
        o_data_forward_reg[369]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__16_ ( .D(N574), .CP(clk), .Q(
        o_data_forward_reg[368]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__15_ ( .D(N573), .CP(clk), .Q(
        o_data_forward_reg[367]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__14_ ( .D(N572), .CP(clk), .Q(
        o_data_forward_reg[366]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__13_ ( .D(N571), .CP(clk), .Q(
        o_data_forward_reg[365]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__12_ ( .D(N570), .CP(clk), .Q(
        o_data_forward_reg[364]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__11_ ( .D(N569), .CP(clk), .Q(
        o_data_forward_reg[363]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__10_ ( .D(N568), .CP(clk), .Q(
        o_data_forward_reg[362]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__9_ ( .D(N567), .CP(clk), .Q(
        o_data_forward_reg[361]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__8_ ( .D(N566), .CP(clk), .Q(
        o_data_forward_reg[360]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__7_ ( .D(N565), .CP(clk), .Q(
        o_data_forward_reg[359]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__6_ ( .D(N564), .CP(clk), .Q(
        o_data_forward_reg[358]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__5_ ( .D(N563), .CP(clk), .Q(
        o_data_forward_reg[357]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__4_ ( .D(N562), .CP(clk), .Q(
        o_data_forward_reg[356]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__3_ ( .D(N561), .CP(clk), .Q(
        o_data_forward_reg[355]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__2_ ( .D(N560), .CP(clk), .Q(
        o_data_forward_reg[354]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__1_ ( .D(N559), .CP(clk), .Q(
        o_data_forward_reg[353]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__0_ ( .D(N558), .CP(clk), .Q(
        o_data_forward_reg[352]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_3_ ( .D(N590), .CP(clk), .Q(
        o_valid_forward_reg[3]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_4__3_ ( .D(N730), .CP(clk), .Q(
        o_cmd_forward_reg[43]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_4__2_ ( .D(n290), .CP(clk), .Q(
        o_cmd_forward_reg[42]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_4__1_ ( .D(N728), .CP(clk), .Q(
        o_cmd_forward_reg[41]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_4__0_ ( .D(N727), .CP(clk), .Q(
        o_cmd_forward_reg[40]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__31_ ( .D(N725), .CP(clk), .Q(
        o_data_forward_reg[351]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__30_ ( .D(N724), .CP(clk), .Q(
        o_data_forward_reg[350]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__29_ ( .D(N723), .CP(clk), .Q(
        o_data_forward_reg[349]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__28_ ( .D(N722), .CP(clk), .Q(
        o_data_forward_reg[348]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__27_ ( .D(N721), .CP(clk), .Q(
        o_data_forward_reg[347]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__26_ ( .D(N720), .CP(clk), .Q(
        o_data_forward_reg[346]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__25_ ( .D(N719), .CP(clk), .Q(
        o_data_forward_reg[345]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__24_ ( .D(N718), .CP(clk), .Q(
        o_data_forward_reg[344]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__23_ ( .D(N717), .CP(clk), .Q(
        o_data_forward_reg[343]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__22_ ( .D(N716), .CP(clk), .Q(
        o_data_forward_reg[342]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__21_ ( .D(N715), .CP(clk), .Q(
        o_data_forward_reg[341]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__20_ ( .D(N714), .CP(clk), .Q(
        o_data_forward_reg[340]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__19_ ( .D(N713), .CP(clk), .Q(
        o_data_forward_reg[339]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__18_ ( .D(N712), .CP(clk), .Q(
        o_data_forward_reg[338]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__17_ ( .D(N711), .CP(clk), .Q(
        o_data_forward_reg[337]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__16_ ( .D(N710), .CP(clk), .Q(
        o_data_forward_reg[336]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__15_ ( .D(N709), .CP(clk), .Q(
        o_data_forward_reg[335]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__14_ ( .D(N708), .CP(clk), .Q(
        o_data_forward_reg[334]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__13_ ( .D(N707), .CP(clk), .Q(
        o_data_forward_reg[333]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__12_ ( .D(N706), .CP(clk), .Q(
        o_data_forward_reg[332]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__11_ ( .D(N705), .CP(clk), .Q(
        o_data_forward_reg[331]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__10_ ( .D(N704), .CP(clk), .Q(
        o_data_forward_reg[330]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__9_ ( .D(N703), .CP(clk), .Q(
        o_data_forward_reg[329]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__8_ ( .D(N702), .CP(clk), .Q(
        o_data_forward_reg[328]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__7_ ( .D(N701), .CP(clk), .Q(
        o_data_forward_reg[327]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__6_ ( .D(N700), .CP(clk), .Q(
        o_data_forward_reg[326]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__5_ ( .D(N699), .CP(clk), .Q(
        o_data_forward_reg[325]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__4_ ( .D(N698), .CP(clk), .Q(
        o_data_forward_reg[324]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__3_ ( .D(N697), .CP(clk), .Q(
        o_data_forward_reg[323]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__2_ ( .D(N696), .CP(clk), .Q(
        o_data_forward_reg[322]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__1_ ( .D(N695), .CP(clk), .Q(
        o_data_forward_reg[321]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__0_ ( .D(N694), .CP(clk), .Q(
        o_data_forward_reg[320]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_4_ ( .D(N726), .CP(clk), .Q(
        o_valid_forward_reg[4]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_5__3_ ( .D(N866), .CP(clk), .Q(
        o_cmd_forward_reg[39]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_5__2_ ( .D(N865), .CP(clk), .Q(
        o_cmd_forward_reg[38]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_5__1_ ( .D(N864), .CP(clk), .Q(
        o_cmd_forward_reg[37]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_5__0_ ( .D(n298), .CP(clk), .Q(
        o_cmd_forward_reg[36]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__31_ ( .D(N861), .CP(clk), .Q(
        o_data_forward_reg[319]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__30_ ( .D(N860), .CP(clk), .Q(
        o_data_forward_reg[318]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__29_ ( .D(N859), .CP(clk), .Q(
        o_data_forward_reg[317]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__28_ ( .D(N858), .CP(clk), .Q(
        o_data_forward_reg[316]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__27_ ( .D(N857), .CP(clk), .Q(
        o_data_forward_reg[315]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__26_ ( .D(N856), .CP(clk), .Q(
        o_data_forward_reg[314]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__25_ ( .D(N855), .CP(clk), .Q(
        o_data_forward_reg[313]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__24_ ( .D(N854), .CP(clk), .Q(
        o_data_forward_reg[312]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__23_ ( .D(N853), .CP(clk), .Q(
        o_data_forward_reg[311]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__22_ ( .D(N852), .CP(clk), .Q(
        o_data_forward_reg[310]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__21_ ( .D(N851), .CP(clk), .Q(
        o_data_forward_reg[309]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__20_ ( .D(N850), .CP(clk), .Q(
        o_data_forward_reg[308]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__19_ ( .D(N849), .CP(clk), .Q(
        o_data_forward_reg[307]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__18_ ( .D(N848), .CP(clk), .Q(
        o_data_forward_reg[306]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__17_ ( .D(N847), .CP(clk), .Q(
        o_data_forward_reg[305]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__16_ ( .D(N846), .CP(clk), .Q(
        o_data_forward_reg[304]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__15_ ( .D(N845), .CP(clk), .Q(
        o_data_forward_reg[303]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__14_ ( .D(N844), .CP(clk), .Q(
        o_data_forward_reg[302]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__13_ ( .D(N843), .CP(clk), .Q(
        o_data_forward_reg[301]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__12_ ( .D(N842), .CP(clk), .Q(
        o_data_forward_reg[300]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__11_ ( .D(N841), .CP(clk), .Q(
        o_data_forward_reg[299]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__10_ ( .D(N840), .CP(clk), .Q(
        o_data_forward_reg[298]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__9_ ( .D(N839), .CP(clk), .Q(
        o_data_forward_reg[297]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__8_ ( .D(N838), .CP(clk), .Q(
        o_data_forward_reg[296]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__7_ ( .D(N837), .CP(clk), .Q(
        o_data_forward_reg[295]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__6_ ( .D(N836), .CP(clk), .Q(
        o_data_forward_reg[294]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__5_ ( .D(N835), .CP(clk), .Q(
        o_data_forward_reg[293]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__4_ ( .D(N834), .CP(clk), .Q(
        o_data_forward_reg[292]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__3_ ( .D(N833), .CP(clk), .Q(
        o_data_forward_reg[291]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__2_ ( .D(N832), .CP(clk), .Q(
        o_data_forward_reg[290]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__1_ ( .D(N831), .CP(clk), .Q(
        o_data_forward_reg[289]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__0_ ( .D(N830), .CP(clk), .Q(
        o_data_forward_reg[288]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_5_ ( .D(N862), .CP(clk), .Q(
        o_valid_forward_reg[5]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_6__3_ ( .D(N1002), .CP(clk), .Q(
        o_cmd_forward_reg[35]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_6__2_ ( .D(N1001), .CP(clk), .Q(
        o_cmd_forward_reg[34]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_6__1_ ( .D(n287), .CP(clk), .Q(
        o_cmd_forward_reg[33]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_6__0_ ( .D(N999), .CP(clk), .Q(
        o_cmd_forward_reg[32]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__31_ ( .D(N997), .CP(clk), .Q(
        o_data_forward_reg[287]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__30_ ( .D(N996), .CP(clk), .Q(
        o_data_forward_reg[286]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__29_ ( .D(N995), .CP(clk), .Q(
        o_data_forward_reg[285]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__28_ ( .D(N994), .CP(clk), .Q(
        o_data_forward_reg[284]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__27_ ( .D(N993), .CP(clk), .Q(
        o_data_forward_reg[283]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__26_ ( .D(N992), .CP(clk), .Q(
        o_data_forward_reg[282]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__25_ ( .D(N991), .CP(clk), .Q(
        o_data_forward_reg[281]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__24_ ( .D(N990), .CP(clk), .Q(
        o_data_forward_reg[280]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__23_ ( .D(N989), .CP(clk), .Q(
        o_data_forward_reg[279]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__22_ ( .D(N988), .CP(clk), .Q(
        o_data_forward_reg[278]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__21_ ( .D(N987), .CP(clk), .Q(
        o_data_forward_reg[277]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__20_ ( .D(N986), .CP(clk), .Q(
        o_data_forward_reg[276]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__19_ ( .D(N985), .CP(clk), .Q(
        o_data_forward_reg[275]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__18_ ( .D(N984), .CP(clk), .Q(
        o_data_forward_reg[274]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__17_ ( .D(N983), .CP(clk), .Q(
        o_data_forward_reg[273]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__16_ ( .D(N982), .CP(clk), .Q(
        o_data_forward_reg[272]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__15_ ( .D(N981), .CP(clk), .Q(
        o_data_forward_reg[271]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__14_ ( .D(N980), .CP(clk), .Q(
        o_data_forward_reg[270]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__13_ ( .D(N979), .CP(clk), .Q(
        o_data_forward_reg[269]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__12_ ( .D(N978), .CP(clk), .Q(
        o_data_forward_reg[268]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__11_ ( .D(N977), .CP(clk), .Q(
        o_data_forward_reg[267]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__10_ ( .D(N976), .CP(clk), .Q(
        o_data_forward_reg[266]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__9_ ( .D(N975), .CP(clk), .Q(
        o_data_forward_reg[265]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__8_ ( .D(N974), .CP(clk), .Q(
        o_data_forward_reg[264]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__7_ ( .D(N973), .CP(clk), .Q(
        o_data_forward_reg[263]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__6_ ( .D(N972), .CP(clk), .Q(
        o_data_forward_reg[262]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__5_ ( .D(N971), .CP(clk), .Q(
        o_data_forward_reg[261]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__4_ ( .D(N970), .CP(clk), .Q(
        o_data_forward_reg[260]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__3_ ( .D(N969), .CP(clk), .Q(
        o_data_forward_reg[259]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__2_ ( .D(N968), .CP(clk), .Q(
        o_data_forward_reg[258]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__1_ ( .D(N967), .CP(clk), .Q(
        o_data_forward_reg[257]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__0_ ( .D(N966), .CP(clk), .Q(
        o_data_forward_reg[256]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_6_ ( .D(N998), .CP(clk), .Q(
        o_valid_forward_reg[6]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_7__3_ ( .D(N1138), .CP(clk), .Q(
        o_cmd_forward_reg[31]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_7__2_ ( .D(n301), .CP(clk), .Q(
        o_cmd_forward_reg[30]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_7__1_ ( .D(N1136), .CP(clk), .Q(
        o_cmd_forward_reg[29]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_7__0_ ( .D(N1135), .CP(clk), .Q(
        o_cmd_forward_reg[28]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__31_ ( .D(N1133), .CP(clk), .Q(
        o_data_forward_reg[255]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__30_ ( .D(N1132), .CP(clk), .Q(
        o_data_forward_reg[254]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__29_ ( .D(N1131), .CP(clk), .Q(
        o_data_forward_reg[253]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__28_ ( .D(N1130), .CP(clk), .Q(
        o_data_forward_reg[252]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__27_ ( .D(N1129), .CP(clk), .Q(
        o_data_forward_reg[251]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__26_ ( .D(N1128), .CP(clk), .Q(
        o_data_forward_reg[250]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__25_ ( .D(N1127), .CP(clk), .Q(
        o_data_forward_reg[249]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__24_ ( .D(N1126), .CP(clk), .Q(
        o_data_forward_reg[248]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__23_ ( .D(N1125), .CP(clk), .Q(
        o_data_forward_reg[247]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__22_ ( .D(N1124), .CP(clk), .Q(
        o_data_forward_reg[246]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__21_ ( .D(N1123), .CP(clk), .Q(
        o_data_forward_reg[245]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__20_ ( .D(N1122), .CP(clk), .Q(
        o_data_forward_reg[244]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__19_ ( .D(N1121), .CP(clk), .Q(
        o_data_forward_reg[243]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__18_ ( .D(N1120), .CP(clk), .Q(
        o_data_forward_reg[242]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__17_ ( .D(N1119), .CP(clk), .Q(
        o_data_forward_reg[241]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__16_ ( .D(N1118), .CP(clk), .Q(
        o_data_forward_reg[240]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__15_ ( .D(N1117), .CP(clk), .Q(
        o_data_forward_reg[239]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__14_ ( .D(N1116), .CP(clk), .Q(
        o_data_forward_reg[238]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__13_ ( .D(N1115), .CP(clk), .Q(
        o_data_forward_reg[237]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__12_ ( .D(N1114), .CP(clk), .Q(
        o_data_forward_reg[236]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__11_ ( .D(N1113), .CP(clk), .Q(
        o_data_forward_reg[235]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__10_ ( .D(N1112), .CP(clk), .Q(
        o_data_forward_reg[234]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__9_ ( .D(N1111), .CP(clk), .Q(
        o_data_forward_reg[233]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__8_ ( .D(N1110), .CP(clk), .Q(
        o_data_forward_reg[232]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__7_ ( .D(N1109), .CP(clk), .Q(
        o_data_forward_reg[231]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__6_ ( .D(N1108), .CP(clk), .Q(
        o_data_forward_reg[230]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__5_ ( .D(N1107), .CP(clk), .Q(
        o_data_forward_reg[229]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__4_ ( .D(N1106), .CP(clk), .Q(
        o_data_forward_reg[228]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__3_ ( .D(N1105), .CP(clk), .Q(
        o_data_forward_reg[227]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__2_ ( .D(N1104), .CP(clk), .Q(
        o_data_forward_reg[226]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__1_ ( .D(N1103), .CP(clk), .Q(
        o_data_forward_reg[225]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__0_ ( .D(N1102), .CP(clk), .Q(
        o_data_forward_reg[224]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_7_ ( .D(N1134), .CP(clk), .Q(
        o_valid_forward_reg[7]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_8__3_ ( .D(n284), .CP(clk), .Q(
        o_cmd_forward_reg[27]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_8__2_ ( .D(N1273), .CP(clk), .Q(
        o_cmd_forward_reg[26]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_8__1_ ( .D(N1272), .CP(clk), .Q(
        o_cmd_forward_reg[25]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_8__0_ ( .D(N1271), .CP(clk), .Q(
        o_cmd_forward_reg[24]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__31_ ( .D(N1269), .CP(clk), .Q(
        o_data_forward_reg[223]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__30_ ( .D(N1268), .CP(clk), .Q(
        o_data_forward_reg[222]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__29_ ( .D(N1267), .CP(clk), .Q(
        o_data_forward_reg[221]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__28_ ( .D(N1266), .CP(clk), .Q(
        o_data_forward_reg[220]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__27_ ( .D(N1265), .CP(clk), .Q(
        o_data_forward_reg[219]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__26_ ( .D(N1264), .CP(clk), .Q(
        o_data_forward_reg[218]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__25_ ( .D(N1263), .CP(clk), .Q(
        o_data_forward_reg[217]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__24_ ( .D(N1262), .CP(clk), .Q(
        o_data_forward_reg[216]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__23_ ( .D(N1261), .CP(clk), .Q(
        o_data_forward_reg[215]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__22_ ( .D(N1260), .CP(clk), .Q(
        o_data_forward_reg[214]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__21_ ( .D(N1259), .CP(clk), .Q(
        o_data_forward_reg[213]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__20_ ( .D(N1258), .CP(clk), .Q(
        o_data_forward_reg[212]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__19_ ( .D(N1257), .CP(clk), .Q(
        o_data_forward_reg[211]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__18_ ( .D(N1256), .CP(clk), .Q(
        o_data_forward_reg[210]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__17_ ( .D(N1255), .CP(clk), .Q(
        o_data_forward_reg[209]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__16_ ( .D(N1254), .CP(clk), .Q(
        o_data_forward_reg[208]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__15_ ( .D(N1253), .CP(clk), .Q(
        o_data_forward_reg[207]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__14_ ( .D(N1252), .CP(clk), .Q(
        o_data_forward_reg[206]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__13_ ( .D(N1251), .CP(clk), .Q(
        o_data_forward_reg[205]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__12_ ( .D(N1250), .CP(clk), .Q(
        o_data_forward_reg[204]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__11_ ( .D(N1249), .CP(clk), .Q(
        o_data_forward_reg[203]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__10_ ( .D(N1248), .CP(clk), .Q(
        o_data_forward_reg[202]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__9_ ( .D(N1247), .CP(clk), .Q(
        o_data_forward_reg[201]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__8_ ( .D(N1246), .CP(clk), .Q(
        o_data_forward_reg[200]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__7_ ( .D(N1245), .CP(clk), .Q(
        o_data_forward_reg[199]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__6_ ( .D(N1244), .CP(clk), .Q(
        o_data_forward_reg[198]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__5_ ( .D(N1243), .CP(clk), .Q(
        o_data_forward_reg[197]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__4_ ( .D(N1242), .CP(clk), .Q(
        o_data_forward_reg[196]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__3_ ( .D(N1241), .CP(clk), .Q(
        o_data_forward_reg[195]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__2_ ( .D(N1240), .CP(clk), .Q(
        o_data_forward_reg[194]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__1_ ( .D(N1239), .CP(clk), .Q(
        o_data_forward_reg[193]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__0_ ( .D(N1238), .CP(clk), .Q(
        o_data_forward_reg[192]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_8_ ( .D(N1270), .CP(clk), .Q(
        o_valid_forward_reg[8]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_9__3_ ( .D(N1410), .CP(clk), .Q(
        o_cmd_forward_reg[23]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_9__2_ ( .D(N1409), .CP(clk), .Q(
        o_cmd_forward_reg[22]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_9__1_ ( .D(N1408), .CP(clk), .Q(
        o_cmd_forward_reg[21]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_9__0_ ( .D(n299), .CP(clk), .Q(
        o_cmd_forward_reg[20]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__31_ ( .D(N1405), .CP(clk), .Q(
        o_data_forward_reg[191]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__30_ ( .D(N1404), .CP(clk), .Q(
        o_data_forward_reg[190]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__29_ ( .D(N1403), .CP(clk), .Q(
        o_data_forward_reg[189]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__28_ ( .D(N1402), .CP(clk), .Q(
        o_data_forward_reg[188]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__27_ ( .D(N1401), .CP(clk), .Q(
        o_data_forward_reg[187]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__26_ ( .D(N1400), .CP(clk), .Q(
        o_data_forward_reg[186]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__25_ ( .D(N1399), .CP(clk), .Q(
        o_data_forward_reg[185]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__24_ ( .D(N1398), .CP(clk), .Q(
        o_data_forward_reg[184]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__23_ ( .D(N1397), .CP(clk), .Q(
        o_data_forward_reg[183]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__22_ ( .D(N1396), .CP(clk), .Q(
        o_data_forward_reg[182]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__21_ ( .D(N1395), .CP(clk), .Q(
        o_data_forward_reg[181]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__20_ ( .D(N1394), .CP(clk), .Q(
        o_data_forward_reg[180]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__19_ ( .D(N1393), .CP(clk), .Q(
        o_data_forward_reg[179]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__18_ ( .D(N1392), .CP(clk), .Q(
        o_data_forward_reg[178]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__17_ ( .D(N1391), .CP(clk), .Q(
        o_data_forward_reg[177]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__16_ ( .D(N1390), .CP(clk), .Q(
        o_data_forward_reg[176]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__15_ ( .D(N1389), .CP(clk), .Q(
        o_data_forward_reg[175]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__14_ ( .D(N1388), .CP(clk), .Q(
        o_data_forward_reg[174]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__13_ ( .D(N1387), .CP(clk), .Q(
        o_data_forward_reg[173]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__12_ ( .D(N1386), .CP(clk), .Q(
        o_data_forward_reg[172]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__11_ ( .D(N1385), .CP(clk), .Q(
        o_data_forward_reg[171]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__10_ ( .D(N1384), .CP(clk), .Q(
        o_data_forward_reg[170]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__9_ ( .D(N1383), .CP(clk), .Q(
        o_data_forward_reg[169]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__8_ ( .D(N1382), .CP(clk), .Q(
        o_data_forward_reg[168]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__7_ ( .D(N1381), .CP(clk), .Q(
        o_data_forward_reg[167]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__6_ ( .D(N1380), .CP(clk), .Q(
        o_data_forward_reg[166]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__5_ ( .D(N1379), .CP(clk), .Q(
        o_data_forward_reg[165]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__4_ ( .D(N1378), .CP(clk), .Q(
        o_data_forward_reg[164]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__3_ ( .D(N1377), .CP(clk), .Q(
        o_data_forward_reg[163]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__2_ ( .D(N1376), .CP(clk), .Q(
        o_data_forward_reg[162]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__1_ ( .D(N1375), .CP(clk), .Q(
        o_data_forward_reg[161]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__0_ ( .D(N1374), .CP(clk), .Q(
        o_data_forward_reg[160]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_9_ ( .D(N1406), .CP(clk), .Q(
        o_valid_forward_reg[9]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_10__3_ ( .D(n300), .CP(clk), .Q(
        o_cmd_forward_reg[19]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_10__2_ ( .D(N1545), .CP(clk), .Q(
        o_cmd_forward_reg[18]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_10__1_ ( .D(N1544), .CP(clk), .Q(
        o_cmd_forward_reg[17]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_10__0_ ( .D(N1543), .CP(clk), .Q(
        o_cmd_forward_reg[16]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__31_ ( .D(N1541), .CP(clk), .Q(
        o_data_forward_reg[159]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__30_ ( .D(N1540), .CP(clk), .Q(
        o_data_forward_reg[158]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__29_ ( .D(N1539), .CP(clk), .Q(
        o_data_forward_reg[157]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__28_ ( .D(N1538), .CP(clk), .Q(
        o_data_forward_reg[156]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__27_ ( .D(N1537), .CP(clk), .Q(
        o_data_forward_reg[155]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__26_ ( .D(N1536), .CP(clk), .Q(
        o_data_forward_reg[154]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__25_ ( .D(N1535), .CP(clk), .Q(
        o_data_forward_reg[153]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__24_ ( .D(N1534), .CP(clk), .Q(
        o_data_forward_reg[152]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__23_ ( .D(N1533), .CP(clk), .Q(
        o_data_forward_reg[151]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__22_ ( .D(N1532), .CP(clk), .Q(
        o_data_forward_reg[150]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__21_ ( .D(N1531), .CP(clk), .Q(
        o_data_forward_reg[149]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__20_ ( .D(N1530), .CP(clk), .Q(
        o_data_forward_reg[148]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__19_ ( .D(N1529), .CP(clk), .Q(
        o_data_forward_reg[147]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__18_ ( .D(N1528), .CP(clk), .Q(
        o_data_forward_reg[146]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__17_ ( .D(N1527), .CP(clk), .Q(
        o_data_forward_reg[145]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__16_ ( .D(N1526), .CP(clk), .Q(
        o_data_forward_reg[144]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__15_ ( .D(N1525), .CP(clk), .Q(
        o_data_forward_reg[143]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__14_ ( .D(N1524), .CP(clk), .Q(
        o_data_forward_reg[142]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__13_ ( .D(N1523), .CP(clk), .Q(
        o_data_forward_reg[141]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__12_ ( .D(N1522), .CP(clk), .Q(
        o_data_forward_reg[140]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__11_ ( .D(N1521), .CP(clk), .Q(
        o_data_forward_reg[139]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__10_ ( .D(N1520), .CP(clk), .Q(
        o_data_forward_reg[138]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__9_ ( .D(N1519), .CP(clk), .Q(
        o_data_forward_reg[137]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__8_ ( .D(N1518), .CP(clk), .Q(
        o_data_forward_reg[136]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__7_ ( .D(N1517), .CP(clk), .Q(
        o_data_forward_reg[135]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__6_ ( .D(N1516), .CP(clk), .Q(
        o_data_forward_reg[134]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__5_ ( .D(N1515), .CP(clk), .Q(
        o_data_forward_reg[133]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__4_ ( .D(N1514), .CP(clk), .Q(
        o_data_forward_reg[132]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__3_ ( .D(N1513), .CP(clk), .Q(
        o_data_forward_reg[131]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__2_ ( .D(N1512), .CP(clk), .Q(
        o_data_forward_reg[130]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__1_ ( .D(N1511), .CP(clk), .Q(
        o_data_forward_reg[129]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__0_ ( .D(N1510), .CP(clk), .Q(
        o_data_forward_reg[128]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_10_ ( .D(N1542), .CP(clk), .Q(
        o_valid_forward_reg[10]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_11__3_ ( .D(N1682), .CP(clk), .Q(
        o_cmd_forward_reg[15]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_11__2_ ( .D(N1681), .CP(clk), .Q(
        o_cmd_forward_reg[14]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_11__1_ ( .D(n302), .CP(clk), .Q(
        o_cmd_forward_reg[13]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_11__0_ ( .D(N1679), .CP(clk), .Q(
        o_cmd_forward_reg[12]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__31_ ( .D(N1677), .CP(clk), .Q(
        o_data_forward_reg[127]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__30_ ( .D(N1676), .CP(clk), .Q(
        o_data_forward_reg[126]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__29_ ( .D(N1675), .CP(clk), .Q(
        o_data_forward_reg[125]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__28_ ( .D(N1674), .CP(clk), .Q(
        o_data_forward_reg[124]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__27_ ( .D(N1673), .CP(clk), .Q(
        o_data_forward_reg[123]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__26_ ( .D(N1672), .CP(clk), .Q(
        o_data_forward_reg[122]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__25_ ( .D(N1671), .CP(clk), .Q(
        o_data_forward_reg[121]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__24_ ( .D(N1670), .CP(clk), .Q(
        o_data_forward_reg[120]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__23_ ( .D(N1669), .CP(clk), .Q(
        o_data_forward_reg[119]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__22_ ( .D(N1668), .CP(clk), .Q(
        o_data_forward_reg[118]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__21_ ( .D(N1667), .CP(clk), .Q(
        o_data_forward_reg[117]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__20_ ( .D(N1666), .CP(clk), .Q(
        o_data_forward_reg[116]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__19_ ( .D(N1665), .CP(clk), .Q(
        o_data_forward_reg[115]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__18_ ( .D(N1664), .CP(clk), .Q(
        o_data_forward_reg[114]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__17_ ( .D(N1663), .CP(clk), .Q(
        o_data_forward_reg[113]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__16_ ( .D(N1662), .CP(clk), .Q(
        o_data_forward_reg[112]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__15_ ( .D(N1661), .CP(clk), .Q(
        o_data_forward_reg[111]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__14_ ( .D(N1660), .CP(clk), .Q(
        o_data_forward_reg[110]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__13_ ( .D(N1659), .CP(clk), .Q(
        o_data_forward_reg[109]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__12_ ( .D(N1658), .CP(clk), .Q(
        o_data_forward_reg[108]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__11_ ( .D(N1657), .CP(clk), .Q(
        o_data_forward_reg[107]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__10_ ( .D(N1656), .CP(clk), .Q(
        o_data_forward_reg[106]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__9_ ( .D(N1655), .CP(clk), .Q(
        o_data_forward_reg[105]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__8_ ( .D(N1654), .CP(clk), .Q(
        o_data_forward_reg[104]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__7_ ( .D(N1653), .CP(clk), .Q(
        o_data_forward_reg[103]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__6_ ( .D(N1652), .CP(clk), .Q(
        o_data_forward_reg[102]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__5_ ( .D(N1651), .CP(clk), .Q(
        o_data_forward_reg[101]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__4_ ( .D(N1650), .CP(clk), .Q(
        o_data_forward_reg[100]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__3_ ( .D(N1649), .CP(clk), .Q(
        o_data_forward_reg[99]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__2_ ( .D(N1648), .CP(clk), .Q(
        o_data_forward_reg[98]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__1_ ( .D(N1647), .CP(clk), .Q(
        o_data_forward_reg[97]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__0_ ( .D(N1646), .CP(clk), .Q(
        o_data_forward_reg[96]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_11_ ( .D(N1678), .CP(clk), .Q(
        o_valid_forward_reg[11]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_12__3_ ( .D(n304), .CP(clk), .Q(
        o_cmd_forward_reg[11]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_12__2_ ( .D(N1817), .CP(clk), .Q(
        o_cmd_forward_reg[10]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_12__1_ ( .D(N1816), .CP(clk), .Q(
        o_cmd_forward_reg[9]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_12__0_ ( .D(N1815), .CP(clk), .Q(
        o_cmd_forward_reg[8]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__31_ ( .D(N1813), .CP(clk), .Q(
        o_data_forward_reg[95]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__30_ ( .D(N1812), .CP(clk), .Q(
        o_data_forward_reg[94]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__29_ ( .D(N1811), .CP(clk), .Q(
        o_data_forward_reg[93]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__28_ ( .D(N1810), .CP(clk), .Q(
        o_data_forward_reg[92]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__27_ ( .D(N1809), .CP(clk), .Q(
        o_data_forward_reg[91]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__26_ ( .D(N1808), .CP(clk), .Q(
        o_data_forward_reg[90]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__25_ ( .D(N1807), .CP(clk), .Q(
        o_data_forward_reg[89]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__24_ ( .D(N1806), .CP(clk), .Q(
        o_data_forward_reg[88]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__23_ ( .D(N1805), .CP(clk), .Q(
        o_data_forward_reg[87]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__22_ ( .D(N1804), .CP(clk), .Q(
        o_data_forward_reg[86]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__21_ ( .D(N1803), .CP(clk), .Q(
        o_data_forward_reg[85]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__20_ ( .D(N1802), .CP(clk), .Q(
        o_data_forward_reg[84]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__19_ ( .D(N1801), .CP(clk), .Q(
        o_data_forward_reg[83]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__18_ ( .D(N1800), .CP(clk), .Q(
        o_data_forward_reg[82]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__17_ ( .D(N1799), .CP(clk), .Q(
        o_data_forward_reg[81]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__16_ ( .D(N1798), .CP(clk), .Q(
        o_data_forward_reg[80]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__15_ ( .D(N1797), .CP(clk), .Q(
        o_data_forward_reg[79]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__14_ ( .D(N1796), .CP(clk), .Q(
        o_data_forward_reg[78]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__13_ ( .D(N1795), .CP(clk), .Q(
        o_data_forward_reg[77]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__12_ ( .D(N1794), .CP(clk), .Q(
        o_data_forward_reg[76]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__11_ ( .D(N1793), .CP(clk), .Q(
        o_data_forward_reg[75]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__10_ ( .D(N1792), .CP(clk), .Q(
        o_data_forward_reg[74]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__9_ ( .D(N1791), .CP(clk), .Q(
        o_data_forward_reg[73]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__8_ ( .D(N1790), .CP(clk), .Q(
        o_data_forward_reg[72]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__7_ ( .D(N1789), .CP(clk), .Q(
        o_data_forward_reg[71]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__6_ ( .D(N1788), .CP(clk), .Q(
        o_data_forward_reg[70]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__5_ ( .D(N1787), .CP(clk), .Q(
        o_data_forward_reg[69]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__4_ ( .D(N1786), .CP(clk), .Q(
        o_data_forward_reg[68]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__3_ ( .D(N1785), .CP(clk), .Q(
        o_data_forward_reg[67]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__2_ ( .D(N1784), .CP(clk), .Q(
        o_data_forward_reg[66]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__1_ ( .D(N1783), .CP(clk), .Q(
        o_data_forward_reg[65]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__0_ ( .D(N1782), .CP(clk), .Q(
        o_data_forward_reg[64]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_12_ ( .D(N1814), .CP(clk), .Q(
        o_valid_forward_reg[12]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_13__3_ ( .D(n303), .CP(clk), .Q(
        o_cmd_forward_reg[7]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_13__2_ ( .D(N1953), .CP(clk), .Q(
        o_cmd_forward_reg[6]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_13__1_ ( .D(N1952), .CP(clk), .Q(
        o_cmd_forward_reg[5]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_13__0_ ( .D(N1951), .CP(clk), .Q(
        o_cmd_forward_reg[4]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__31_ ( .D(N1949), .CP(clk), .Q(
        o_data_forward_reg[63]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__30_ ( .D(N1948), .CP(clk), .Q(
        o_data_forward_reg[62]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__29_ ( .D(N1947), .CP(clk), .Q(
        o_data_forward_reg[61]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__28_ ( .D(N1946), .CP(clk), .Q(
        o_data_forward_reg[60]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__27_ ( .D(N1945), .CP(clk), .Q(
        o_data_forward_reg[59]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__26_ ( .D(N1944), .CP(clk), .Q(
        o_data_forward_reg[58]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__25_ ( .D(N1943), .CP(clk), .Q(
        o_data_forward_reg[57]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__24_ ( .D(N1942), .CP(clk), .Q(
        o_data_forward_reg[56]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__23_ ( .D(N1941), .CP(clk), .Q(
        o_data_forward_reg[55]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__22_ ( .D(N1940), .CP(clk), .Q(
        o_data_forward_reg[54]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__21_ ( .D(N1939), .CP(clk), .Q(
        o_data_forward_reg[53]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__20_ ( .D(N1938), .CP(clk), .Q(
        o_data_forward_reg[52]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__19_ ( .D(N1937), .CP(clk), .Q(
        o_data_forward_reg[51]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__18_ ( .D(N1936), .CP(clk), .Q(
        o_data_forward_reg[50]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__17_ ( .D(N1935), .CP(clk), .Q(
        o_data_forward_reg[49]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__16_ ( .D(N1934), .CP(clk), .Q(
        o_data_forward_reg[48]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__15_ ( .D(N1933), .CP(clk), .Q(
        o_data_forward_reg[47]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__14_ ( .D(N1932), .CP(clk), .Q(
        o_data_forward_reg[46]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__13_ ( .D(N1931), .CP(clk), .Q(
        o_data_forward_reg[45]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__12_ ( .D(N1930), .CP(clk), .Q(
        o_data_forward_reg[44]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__11_ ( .D(N1929), .CP(clk), .Q(
        o_data_forward_reg[43]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__10_ ( .D(N1928), .CP(clk), .Q(
        o_data_forward_reg[42]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__9_ ( .D(N1927), .CP(clk), .Q(
        o_data_forward_reg[41]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__8_ ( .D(N1926), .CP(clk), .Q(
        o_data_forward_reg[40]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__7_ ( .D(N1925), .CP(clk), .Q(
        o_data_forward_reg[39]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__6_ ( .D(N1924), .CP(clk), .Q(
        o_data_forward_reg[38]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__5_ ( .D(N1923), .CP(clk), .Q(
        o_data_forward_reg[37]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__4_ ( .D(N1922), .CP(clk), .Q(
        o_data_forward_reg[36]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__3_ ( .D(N1921), .CP(clk), .Q(
        o_data_forward_reg[35]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__2_ ( .D(N1920), .CP(clk), .Q(
        o_data_forward_reg[34]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__1_ ( .D(N1919), .CP(clk), .Q(
        o_data_forward_reg[33]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__0_ ( .D(N1918), .CP(clk), .Q(
        o_data_forward_reg[32]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_13_ ( .D(N1950), .CP(clk), .Q(
        o_valid_forward_reg[13]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_14__3_ ( .D(N2090), .CP(clk), .Q(
        o_cmd_forward_reg[3]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_14__2_ ( .D(n277), .CP(clk), .Q(
        o_cmd_forward_reg[2]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_14__1_ ( .D(N2088), .CP(clk), .Q(
        o_cmd_forward_reg[1]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_14__0_ ( .D(N2087), .CP(clk), .Q(
        o_cmd_forward_reg[0]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__31_ ( .D(N2085), .CP(clk), .Q(
        o_data_forward_reg[31]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__30_ ( .D(N2084), .CP(clk), .Q(
        o_data_forward_reg[30]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__29_ ( .D(N2083), .CP(clk), .Q(
        o_data_forward_reg[29]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__28_ ( .D(N2082), .CP(clk), .Q(
        o_data_forward_reg[28]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__27_ ( .D(N2081), .CP(clk), .Q(
        o_data_forward_reg[27]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__26_ ( .D(N2080), .CP(clk), .Q(
        o_data_forward_reg[26]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__25_ ( .D(N2079), .CP(clk), .Q(
        o_data_forward_reg[25]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__24_ ( .D(N2078), .CP(clk), .Q(
        o_data_forward_reg[24]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__23_ ( .D(N2077), .CP(clk), .Q(
        o_data_forward_reg[23]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__22_ ( .D(N2076), .CP(clk), .Q(
        o_data_forward_reg[22]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__21_ ( .D(N2075), .CP(clk), .Q(
        o_data_forward_reg[21]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__20_ ( .D(N2074), .CP(clk), .Q(
        o_data_forward_reg[20]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__19_ ( .D(N2073), .CP(clk), .Q(
        o_data_forward_reg[19]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__18_ ( .D(N2072), .CP(clk), .Q(
        o_data_forward_reg[18]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__17_ ( .D(N2071), .CP(clk), .Q(
        o_data_forward_reg[17]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__16_ ( .D(N2070), .CP(clk), .Q(
        o_data_forward_reg[16]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__15_ ( .D(N2069), .CP(clk), .Q(
        o_data_forward_reg[15]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__14_ ( .D(N2068), .CP(clk), .Q(
        o_data_forward_reg[14]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__13_ ( .D(N2067), .CP(clk), .Q(
        o_data_forward_reg[13]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__12_ ( .D(N2066), .CP(clk), .Q(
        o_data_forward_reg[12]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__11_ ( .D(N2065), .CP(clk), .Q(
        o_data_forward_reg[11]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__10_ ( .D(N2064), .CP(clk), .Q(
        o_data_forward_reg[10]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__9_ ( .D(N2063), .CP(clk), .Q(
        o_data_forward_reg[9]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__8_ ( .D(N2062), .CP(clk), .Q(
        o_data_forward_reg[8]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__7_ ( .D(N2061), .CP(clk), .Q(
        o_data_forward_reg[7]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__6_ ( .D(N2060), .CP(clk), .Q(
        o_data_forward_reg[6]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__5_ ( .D(N2059), .CP(clk), .Q(
        o_data_forward_reg[5]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__4_ ( .D(N2058), .CP(clk), .Q(
        o_data_forward_reg[4]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__3_ ( .D(N2057), .CP(clk), .Q(
        o_data_forward_reg[3]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__2_ ( .D(N2056), .CP(clk), .Q(
        o_data_forward_reg[2]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__1_ ( .D(N2055), .CP(clk), .Q(
        o_data_forward_reg[1]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__0_ ( .D(N2054), .CP(clk), .Q(
        o_data_forward_reg[0]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_14_ ( .D(N2086), .CP(clk), .Q(
        o_valid_forward_reg[14]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_15_ ( .D(n275), .CP(clk), .Q(o_valid[15])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_14_ ( .D(n276), .CP(clk), .Q(o_valid[14])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_13_ ( .D(n278), .CP(clk), .Q(o_valid[13])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_12_ ( .D(n20), .CP(clk), .Q(o_valid[12])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_11_ ( .D(n280), .CP(clk), .Q(o_valid[11])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_10_ ( .D(n21), .CP(clk), .Q(o_valid[10])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_9_ ( .D(n282), .CP(clk), .Q(o_valid[9]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_8_ ( .D(n283), .CP(clk), .Q(o_valid[8]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_7_ ( .D(n19), .CP(clk), .Q(o_valid[7]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_6_ ( .D(n286), .CP(clk), .Q(o_valid[6]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_5_ ( .D(n288), .CP(clk), .Q(o_valid[5]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_4_ ( .D(n289), .CP(clk), .Q(o_valid[4]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_3_ ( .D(n291), .CP(clk), .Q(o_valid[3]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_2_ ( .D(n292), .CP(clk), .Q(o_valid[2]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_1_ ( .D(n294), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_0_ ( .D(n274), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_511_ ( .D(n267), .CP(clk), .Q(
        o_data_bus[511]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_510_ ( .D(n266), .CP(clk), .Q(
        o_data_bus[510]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_509_ ( .D(n265), .CP(clk), .Q(
        o_data_bus[509]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_508_ ( .D(n264), .CP(clk), .Q(
        o_data_bus[508]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_507_ ( .D(n263), .CP(clk), .Q(
        o_data_bus[507]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_506_ ( .D(n262), .CP(clk), .Q(
        o_data_bus[506]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_505_ ( .D(n235), .CP(clk), .Q(
        o_data_bus[505]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_504_ ( .D(n234), .CP(clk), .Q(
        o_data_bus[504]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_503_ ( .D(n233), .CP(clk), .Q(
        o_data_bus[503]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_502_ ( .D(n232), .CP(clk), .Q(
        o_data_bus[502]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_501_ ( .D(n231), .CP(clk), .Q(
        o_data_bus[501]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_500_ ( .D(n230), .CP(clk), .Q(
        o_data_bus[500]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_499_ ( .D(n229), .CP(clk), .Q(
        o_data_bus[499]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_498_ ( .D(n228), .CP(clk), .Q(
        o_data_bus[498]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_497_ ( .D(n227), .CP(clk), .Q(
        o_data_bus[497]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_496_ ( .D(n226), .CP(clk), .Q(
        o_data_bus[496]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_495_ ( .D(n225), .CP(clk), .Q(
        o_data_bus[495]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_494_ ( .D(n224), .CP(clk), .Q(
        o_data_bus[494]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_493_ ( .D(n223), .CP(clk), .Q(
        o_data_bus[493]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_492_ ( .D(n222), .CP(clk), .Q(
        o_data_bus[492]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_491_ ( .D(n221), .CP(clk), .Q(
        o_data_bus[491]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_490_ ( .D(n220), .CP(clk), .Q(
        o_data_bus[490]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_489_ ( .D(n219), .CP(clk), .Q(
        o_data_bus[489]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_488_ ( .D(n218), .CP(clk), .Q(
        o_data_bus[488]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_487_ ( .D(n217), .CP(clk), .Q(
        o_data_bus[487]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_486_ ( .D(n216), .CP(clk), .Q(
        o_data_bus[486]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_485_ ( .D(n215), .CP(clk), .Q(
        o_data_bus[485]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_484_ ( .D(n214), .CP(clk), .Q(
        o_data_bus[484]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_483_ ( .D(n213), .CP(clk), .Q(
        o_data_bus[483]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_482_ ( .D(n212), .CP(clk), .Q(
        o_data_bus[482]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_481_ ( .D(n211), .CP(clk), .Q(
        o_data_bus[481]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_480_ ( .D(n210), .CP(clk), .Q(
        o_data_bus[480]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_479_ ( .D(N2053), .CP(clk), .Q(
        o_data_bus[479]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_478_ ( .D(N2052), .CP(clk), .Q(
        o_data_bus[478]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_477_ ( .D(N2051), .CP(clk), .Q(
        o_data_bus[477]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_476_ ( .D(N2050), .CP(clk), .Q(
        o_data_bus[476]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_475_ ( .D(N2049), .CP(clk), .Q(
        o_data_bus[475]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_474_ ( .D(N2048), .CP(clk), .Q(
        o_data_bus[474]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_473_ ( .D(N2047), .CP(clk), .Q(
        o_data_bus[473]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_472_ ( .D(N2046), .CP(clk), .Q(
        o_data_bus[472]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_471_ ( .D(N2045), .CP(clk), .Q(
        o_data_bus[471]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_470_ ( .D(N2044), .CP(clk), .Q(
        o_data_bus[470]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_469_ ( .D(N2043), .CP(clk), .Q(
        o_data_bus[469]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_468_ ( .D(N2042), .CP(clk), .Q(
        o_data_bus[468]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_467_ ( .D(N2041), .CP(clk), .Q(
        o_data_bus[467]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_466_ ( .D(N2040), .CP(clk), .Q(
        o_data_bus[466]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_465_ ( .D(N2039), .CP(clk), .Q(
        o_data_bus[465]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_464_ ( .D(N2038), .CP(clk), .Q(
        o_data_bus[464]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_463_ ( .D(N2037), .CP(clk), .Q(
        o_data_bus[463]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_462_ ( .D(N2036), .CP(clk), .Q(
        o_data_bus[462]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_461_ ( .D(N2035), .CP(clk), .Q(
        o_data_bus[461]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_460_ ( .D(N2034), .CP(clk), .Q(
        o_data_bus[460]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_459_ ( .D(N2033), .CP(clk), .Q(
        o_data_bus[459]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_458_ ( .D(N2032), .CP(clk), .Q(
        o_data_bus[458]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_457_ ( .D(N2031), .CP(clk), .Q(
        o_data_bus[457]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_456_ ( .D(N2030), .CP(clk), .Q(
        o_data_bus[456]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_455_ ( .D(N2029), .CP(clk), .Q(
        o_data_bus[455]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_454_ ( .D(N2028), .CP(clk), .Q(
        o_data_bus[454]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_453_ ( .D(N2027), .CP(clk), .Q(
        o_data_bus[453]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_452_ ( .D(N2026), .CP(clk), .Q(
        o_data_bus[452]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_451_ ( .D(N2025), .CP(clk), .Q(
        o_data_bus[451]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_450_ ( .D(N2024), .CP(clk), .Q(
        o_data_bus[450]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_449_ ( .D(N2023), .CP(clk), .Q(
        o_data_bus[449]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_448_ ( .D(N2022), .CP(clk), .Q(
        o_data_bus[448]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_447_ ( .D(N1917), .CP(clk), .Q(
        o_data_bus[447]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_446_ ( .D(N1916), .CP(clk), .Q(
        o_data_bus[446]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_445_ ( .D(N1915), .CP(clk), .Q(
        o_data_bus[445]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_444_ ( .D(N1914), .CP(clk), .Q(
        o_data_bus[444]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_443_ ( .D(N1913), .CP(clk), .Q(
        o_data_bus[443]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_442_ ( .D(N1912), .CP(clk), .Q(
        o_data_bus[442]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_441_ ( .D(N1911), .CP(clk), .Q(
        o_data_bus[441]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_440_ ( .D(N1910), .CP(clk), .Q(
        o_data_bus[440]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_439_ ( .D(N1909), .CP(clk), .Q(
        o_data_bus[439]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_438_ ( .D(N1908), .CP(clk), .Q(
        o_data_bus[438]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_437_ ( .D(N1907), .CP(clk), .Q(
        o_data_bus[437]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_436_ ( .D(N1906), .CP(clk), .Q(
        o_data_bus[436]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_435_ ( .D(N1905), .CP(clk), .Q(
        o_data_bus[435]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_434_ ( .D(N1904), .CP(clk), .Q(
        o_data_bus[434]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_433_ ( .D(N1903), .CP(clk), .Q(
        o_data_bus[433]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_432_ ( .D(N1902), .CP(clk), .Q(
        o_data_bus[432]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_431_ ( .D(N1901), .CP(clk), .Q(
        o_data_bus[431]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_430_ ( .D(N1900), .CP(clk), .Q(
        o_data_bus[430]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_429_ ( .D(N1899), .CP(clk), .Q(
        o_data_bus[429]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_428_ ( .D(N1898), .CP(clk), .Q(
        o_data_bus[428]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_427_ ( .D(N1897), .CP(clk), .Q(
        o_data_bus[427]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_426_ ( .D(N1896), .CP(clk), .Q(
        o_data_bus[426]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_425_ ( .D(N1895), .CP(clk), .Q(
        o_data_bus[425]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_424_ ( .D(N1894), .CP(clk), .Q(
        o_data_bus[424]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_423_ ( .D(N1893), .CP(clk), .Q(
        o_data_bus[423]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_422_ ( .D(N1892), .CP(clk), .Q(
        o_data_bus[422]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_421_ ( .D(N1891), .CP(clk), .Q(
        o_data_bus[421]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_420_ ( .D(N1890), .CP(clk), .Q(
        o_data_bus[420]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_419_ ( .D(N1889), .CP(clk), .Q(
        o_data_bus[419]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_418_ ( .D(N1888), .CP(clk), .Q(
        o_data_bus[418]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_417_ ( .D(N1887), .CP(clk), .Q(
        o_data_bus[417]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_416_ ( .D(N1886), .CP(clk), .Q(
        o_data_bus[416]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_415_ ( .D(N1781), .CP(clk), .Q(
        o_data_bus[415]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_414_ ( .D(N1780), .CP(clk), .Q(
        o_data_bus[414]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_413_ ( .D(N1779), .CP(clk), .Q(
        o_data_bus[413]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_412_ ( .D(N1778), .CP(clk), .Q(
        o_data_bus[412]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_411_ ( .D(N1777), .CP(clk), .Q(
        o_data_bus[411]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_410_ ( .D(N1776), .CP(clk), .Q(
        o_data_bus[410]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_409_ ( .D(N1775), .CP(clk), .Q(
        o_data_bus[409]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_408_ ( .D(N1774), .CP(clk), .Q(
        o_data_bus[408]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_407_ ( .D(N1773), .CP(clk), .Q(
        o_data_bus[407]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_406_ ( .D(N1772), .CP(clk), .Q(
        o_data_bus[406]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_405_ ( .D(N1771), .CP(clk), .Q(
        o_data_bus[405]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_404_ ( .D(N1770), .CP(clk), .Q(
        o_data_bus[404]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_403_ ( .D(N1769), .CP(clk), .Q(
        o_data_bus[403]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_402_ ( .D(N1768), .CP(clk), .Q(
        o_data_bus[402]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_401_ ( .D(N1767), .CP(clk), .Q(
        o_data_bus[401]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_400_ ( .D(N1766), .CP(clk), .Q(
        o_data_bus[400]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_399_ ( .D(N1765), .CP(clk), .Q(
        o_data_bus[399]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_398_ ( .D(N1764), .CP(clk), .Q(
        o_data_bus[398]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_397_ ( .D(N1763), .CP(clk), .Q(
        o_data_bus[397]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_396_ ( .D(N1762), .CP(clk), .Q(
        o_data_bus[396]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_395_ ( .D(N1761), .CP(clk), .Q(
        o_data_bus[395]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_394_ ( .D(N1760), .CP(clk), .Q(
        o_data_bus[394]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_393_ ( .D(N1759), .CP(clk), .Q(
        o_data_bus[393]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_392_ ( .D(N1758), .CP(clk), .Q(
        o_data_bus[392]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_391_ ( .D(N1757), .CP(clk), .Q(
        o_data_bus[391]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_390_ ( .D(N1756), .CP(clk), .Q(
        o_data_bus[390]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_389_ ( .D(N1755), .CP(clk), .Q(
        o_data_bus[389]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_388_ ( .D(N1754), .CP(clk), .Q(
        o_data_bus[388]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_387_ ( .D(N1753), .CP(clk), .Q(
        o_data_bus[387]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_386_ ( .D(N1752), .CP(clk), .Q(
        o_data_bus[386]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_385_ ( .D(N1751), .CP(clk), .Q(
        o_data_bus[385]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_384_ ( .D(N1750), .CP(clk), .Q(
        o_data_bus[384]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_383_ ( .D(N1645), .CP(clk), .Q(
        o_data_bus[383]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_382_ ( .D(N1644), .CP(clk), .Q(
        o_data_bus[382]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_381_ ( .D(N1643), .CP(clk), .Q(
        o_data_bus[381]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_380_ ( .D(N1642), .CP(clk), .Q(
        o_data_bus[380]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_379_ ( .D(N1641), .CP(clk), .Q(
        o_data_bus[379]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_378_ ( .D(N1640), .CP(clk), .Q(
        o_data_bus[378]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_377_ ( .D(N1639), .CP(clk), .Q(
        o_data_bus[377]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_376_ ( .D(N1638), .CP(clk), .Q(
        o_data_bus[376]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_375_ ( .D(N1637), .CP(clk), .Q(
        o_data_bus[375]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_374_ ( .D(N1636), .CP(clk), .Q(
        o_data_bus[374]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_373_ ( .D(N1635), .CP(clk), .Q(
        o_data_bus[373]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_372_ ( .D(N1634), .CP(clk), .Q(
        o_data_bus[372]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_371_ ( .D(N1633), .CP(clk), .Q(
        o_data_bus[371]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_370_ ( .D(N1632), .CP(clk), .Q(
        o_data_bus[370]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_369_ ( .D(N1631), .CP(clk), .Q(
        o_data_bus[369]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_368_ ( .D(N1630), .CP(clk), .Q(
        o_data_bus[368]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_367_ ( .D(N1629), .CP(clk), .Q(
        o_data_bus[367]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_366_ ( .D(N1628), .CP(clk), .Q(
        o_data_bus[366]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_365_ ( .D(N1627), .CP(clk), .Q(
        o_data_bus[365]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_364_ ( .D(N1626), .CP(clk), .Q(
        o_data_bus[364]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_363_ ( .D(N1625), .CP(clk), .Q(
        o_data_bus[363]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_362_ ( .D(N1624), .CP(clk), .Q(
        o_data_bus[362]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_361_ ( .D(N1623), .CP(clk), .Q(
        o_data_bus[361]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_360_ ( .D(N1622), .CP(clk), .Q(
        o_data_bus[360]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_359_ ( .D(N1621), .CP(clk), .Q(
        o_data_bus[359]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_358_ ( .D(N1620), .CP(clk), .Q(
        o_data_bus[358]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_357_ ( .D(N1619), .CP(clk), .Q(
        o_data_bus[357]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_356_ ( .D(N1618), .CP(clk), .Q(
        o_data_bus[356]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_355_ ( .D(N1617), .CP(clk), .Q(
        o_data_bus[355]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_354_ ( .D(N1616), .CP(clk), .Q(
        o_data_bus[354]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_353_ ( .D(N1615), .CP(clk), .Q(
        o_data_bus[353]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_352_ ( .D(N1614), .CP(clk), .Q(
        o_data_bus[352]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_351_ ( .D(N1509), .CP(clk), .Q(
        o_data_bus[351]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_350_ ( .D(N1508), .CP(clk), .Q(
        o_data_bus[350]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_349_ ( .D(N1507), .CP(clk), .Q(
        o_data_bus[349]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_348_ ( .D(N1506), .CP(clk), .Q(
        o_data_bus[348]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_347_ ( .D(N1505), .CP(clk), .Q(
        o_data_bus[347]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_346_ ( .D(N1504), .CP(clk), .Q(
        o_data_bus[346]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_345_ ( .D(N1503), .CP(clk), .Q(
        o_data_bus[345]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_344_ ( .D(N1502), .CP(clk), .Q(
        o_data_bus[344]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_343_ ( .D(N1501), .CP(clk), .Q(
        o_data_bus[343]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_342_ ( .D(N1500), .CP(clk), .Q(
        o_data_bus[342]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_341_ ( .D(N1499), .CP(clk), .Q(
        o_data_bus[341]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_340_ ( .D(N1498), .CP(clk), .Q(
        o_data_bus[340]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_339_ ( .D(N1497), .CP(clk), .Q(
        o_data_bus[339]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_338_ ( .D(N1496), .CP(clk), .Q(
        o_data_bus[338]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_337_ ( .D(N1495), .CP(clk), .Q(
        o_data_bus[337]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_336_ ( .D(N1494), .CP(clk), .Q(
        o_data_bus[336]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_335_ ( .D(N1493), .CP(clk), .Q(
        o_data_bus[335]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_334_ ( .D(N1492), .CP(clk), .Q(
        o_data_bus[334]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_333_ ( .D(N1491), .CP(clk), .Q(
        o_data_bus[333]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_332_ ( .D(N1490), .CP(clk), .Q(
        o_data_bus[332]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_331_ ( .D(N1489), .CP(clk), .Q(
        o_data_bus[331]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_330_ ( .D(N1488), .CP(clk), .Q(
        o_data_bus[330]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_329_ ( .D(N1487), .CP(clk), .Q(
        o_data_bus[329]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_328_ ( .D(N1486), .CP(clk), .Q(
        o_data_bus[328]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_327_ ( .D(N1485), .CP(clk), .Q(
        o_data_bus[327]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_326_ ( .D(N1484), .CP(clk), .Q(
        o_data_bus[326]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_325_ ( .D(N1483), .CP(clk), .Q(
        o_data_bus[325]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_324_ ( .D(N1482), .CP(clk), .Q(
        o_data_bus[324]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_323_ ( .D(N1481), .CP(clk), .Q(
        o_data_bus[323]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_322_ ( .D(N1480), .CP(clk), .Q(
        o_data_bus[322]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_321_ ( .D(N1479), .CP(clk), .Q(
        o_data_bus[321]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_320_ ( .D(N1478), .CP(clk), .Q(
        o_data_bus[320]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_319_ ( .D(N1373), .CP(clk), .Q(
        o_data_bus[319]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_318_ ( .D(N1372), .CP(clk), .Q(
        o_data_bus[318]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_317_ ( .D(N1371), .CP(clk), .Q(
        o_data_bus[317]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_316_ ( .D(N1370), .CP(clk), .Q(
        o_data_bus[316]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_315_ ( .D(N1369), .CP(clk), .Q(
        o_data_bus[315]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_314_ ( .D(N1368), .CP(clk), .Q(
        o_data_bus[314]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_313_ ( .D(N1367), .CP(clk), .Q(
        o_data_bus[313]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_312_ ( .D(N1366), .CP(clk), .Q(
        o_data_bus[312]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_311_ ( .D(N1365), .CP(clk), .Q(
        o_data_bus[311]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_310_ ( .D(N1364), .CP(clk), .Q(
        o_data_bus[310]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_309_ ( .D(N1363), .CP(clk), .Q(
        o_data_bus[309]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_308_ ( .D(N1362), .CP(clk), .Q(
        o_data_bus[308]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_307_ ( .D(N1361), .CP(clk), .Q(
        o_data_bus[307]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_306_ ( .D(N1360), .CP(clk), .Q(
        o_data_bus[306]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_305_ ( .D(N1359), .CP(clk), .Q(
        o_data_bus[305]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_304_ ( .D(N1358), .CP(clk), .Q(
        o_data_bus[304]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_303_ ( .D(N1357), .CP(clk), .Q(
        o_data_bus[303]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_302_ ( .D(N1356), .CP(clk), .Q(
        o_data_bus[302]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_301_ ( .D(N1355), .CP(clk), .Q(
        o_data_bus[301]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_300_ ( .D(N1354), .CP(clk), .Q(
        o_data_bus[300]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_299_ ( .D(N1353), .CP(clk), .Q(
        o_data_bus[299]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_298_ ( .D(N1352), .CP(clk), .Q(
        o_data_bus[298]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_297_ ( .D(N1351), .CP(clk), .Q(
        o_data_bus[297]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_296_ ( .D(N1350), .CP(clk), .Q(
        o_data_bus[296]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_295_ ( .D(N1349), .CP(clk), .Q(
        o_data_bus[295]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_294_ ( .D(N1348), .CP(clk), .Q(
        o_data_bus[294]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_293_ ( .D(N1347), .CP(clk), .Q(
        o_data_bus[293]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_292_ ( .D(N1346), .CP(clk), .Q(
        o_data_bus[292]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_291_ ( .D(N1345), .CP(clk), .Q(
        o_data_bus[291]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_290_ ( .D(N1344), .CP(clk), .Q(
        o_data_bus[290]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_289_ ( .D(N1343), .CP(clk), .Q(
        o_data_bus[289]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_288_ ( .D(N1342), .CP(clk), .Q(
        o_data_bus[288]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N1101), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N1100), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N1099), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N1098), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N1097), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N1096), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N1095), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N1094), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N1093), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N1092), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N1091), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N1090), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N1089), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N1088), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N1087), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N1086), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N1085), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N1084), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N1083), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N1082), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N1081), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N1080), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N1079), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N1078), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N1077), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N1076), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N1075), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N1074), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N1073), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N1072), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N1071), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N1070), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N965), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N964), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N963), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N962), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N961), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N960), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N959), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N958), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N957), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N956), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N955), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N954), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N953), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N952), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N951), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N950), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N949), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N948), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N947), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N946), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N945), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N944), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N943), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N942), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N941), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N940), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N939), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N938), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N937), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N936), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N935), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N934), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N829), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N828), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N827), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N826), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N825), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N824), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N823), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N822), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N821), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N820), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N819), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N818), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N817), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N816), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N815), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N814), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N813), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N812), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N811), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N810), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N809), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N808), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N807), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N806), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N805), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N804), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N803), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N802), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N801), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N800), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N799), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N798), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N557), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N556), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N555), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N554), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N553), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N552), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N551), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N550), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N549), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N548), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N547), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N546), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N545), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N544), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N543), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N542), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N541), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N540), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N539), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N538), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N537), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N536), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N535), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N534), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N533), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N532), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N531), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N530), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N529), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N528), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N527), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N526), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(n273), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(n272), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(n271), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(n270), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(n269), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(n268), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(n261), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(n260), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(n259), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(n258), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(n257), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(n256), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(n255), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(n254), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(n253), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(n252), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(n251), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(n250), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(n249), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(n248), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(n247), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(n246), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(n245), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(n244), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(n243), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(n242), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(n241), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(n240), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(n239), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(n238), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(n237), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(n236), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_287_ ( .D(N1237), .CP(clk), .Q(
        o_data_bus[287]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_286_ ( .D(N1236), .CP(clk), .Q(
        o_data_bus[286]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_285_ ( .D(N1235), .CP(clk), .Q(
        o_data_bus[285]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_284_ ( .D(N1234), .CP(clk), .Q(
        o_data_bus[284]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_283_ ( .D(N1233), .CP(clk), .Q(
        o_data_bus[283]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_282_ ( .D(N1232), .CP(clk), .Q(
        o_data_bus[282]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_281_ ( .D(N1231), .CP(clk), .Q(
        o_data_bus[281]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_280_ ( .D(N1230), .CP(clk), .Q(
        o_data_bus[280]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_279_ ( .D(N1229), .CP(clk), .Q(
        o_data_bus[279]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_278_ ( .D(N1228), .CP(clk), .Q(
        o_data_bus[278]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_277_ ( .D(N1227), .CP(clk), .Q(
        o_data_bus[277]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_276_ ( .D(N1226), .CP(clk), .Q(
        o_data_bus[276]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_275_ ( .D(N1225), .CP(clk), .Q(
        o_data_bus[275]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_274_ ( .D(N1224), .CP(clk), .Q(
        o_data_bus[274]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_273_ ( .D(N1223), .CP(clk), .Q(
        o_data_bus[273]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_272_ ( .D(N1222), .CP(clk), .Q(
        o_data_bus[272]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_271_ ( .D(N1221), .CP(clk), .Q(
        o_data_bus[271]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_270_ ( .D(N1220), .CP(clk), .Q(
        o_data_bus[270]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_269_ ( .D(N1219), .CP(clk), .Q(
        o_data_bus[269]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_268_ ( .D(N1218), .CP(clk), .Q(
        o_data_bus[268]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_267_ ( .D(N1217), .CP(clk), .Q(
        o_data_bus[267]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_266_ ( .D(N1216), .CP(clk), .Q(
        o_data_bus[266]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_265_ ( .D(N1215), .CP(clk), .Q(
        o_data_bus[265]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_264_ ( .D(N1214), .CP(clk), .Q(
        o_data_bus[264]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_263_ ( .D(N1213), .CP(clk), .Q(
        o_data_bus[263]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_262_ ( .D(N1212), .CP(clk), .Q(
        o_data_bus[262]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_261_ ( .D(N1211), .CP(clk), .Q(
        o_data_bus[261]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_260_ ( .D(N1210), .CP(clk), .Q(
        o_data_bus[260]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_259_ ( .D(N1209), .CP(clk), .Q(
        o_data_bus[259]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_258_ ( .D(N1208), .CP(clk), .Q(
        o_data_bus[258]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_257_ ( .D(N1207), .CP(clk), .Q(
        o_data_bus[257]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_256_ ( .D(N1206), .CP(clk), .Q(
        o_data_bus[256]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N693), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N692), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N691), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N690), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N689), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N688), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N687), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N686), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N685), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N684), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N683), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N682), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N681), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N680), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N679), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N678), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N677), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N676), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N675), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N674), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N673), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N672), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N671), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N670), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N669), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N668), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N667), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N666), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N665), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N664), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N663), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N662), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N265), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N264), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N263), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N262), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N261), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N260), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N259), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N258), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N257), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N256), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N255), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N254), .CP(clk), .Q(
        o_data_bus[32]) );
  ND2OPTIBD1BWP30P140LVT U1103 ( .A1(n22), .A2(n27), .ZN(n28) );
  INR2D1BWP30P140LVT U1104 ( .A1(o_cmd_forward_reg[15]), .B1(n18), .ZN(n304)
         );
  INR2D1BWP30P140LVT U1105 ( .A1(o_cmd_forward_reg[23]), .B1(n18), .ZN(n300)
         );
  INR2D1BWP30P140LVT U1106 ( .A1(o_cmd_forward_reg[34]), .B1(n18), .ZN(n301)
         );
  NR3D1P5BWP30P140LVT U1107 ( .A1(n26), .A2(n25), .A3(n24), .ZN(n275) );
  INVD2BWP30P140LVT U1108 ( .I(n48), .ZN(n18) );
  NR2D1BWP30P140LVT U1109 ( .A1(o_cmd_forward_reg[25]), .A2(
        o_cmd_forward_reg[26]), .ZN(n47) );
  NR2D1BWP30P140LVT U1110 ( .A1(o_cmd_forward_reg[41]), .A2(
        o_cmd_forward_reg[43]), .ZN(n46) );
  ND2D1BWP30P140LVT U1111 ( .A1(n23), .A2(i_en), .ZN(n49) );
  NR2D1BWP30P140LVT U1112 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n27) );
  NR2D1BWP30P140LVT U1113 ( .A1(i_cmd[0]), .A2(i_cmd[1]), .ZN(n29) );
  CKAN2D1BWP30P140LVT U1114 ( .A1(i_valid), .A2(n48), .Z(n22) );
  CKAN2D1BWP30P140LVT U1115 ( .A1(o_cmd_forward_reg[24]), .A2(n48), .Z(n299)
         );
  CKAN2D1BWP30P140LVT U1116 ( .A1(o_cmd_forward_reg[40]), .A2(n48), .Z(n298)
         );
  CKAN2D1BWP30P140LVT U1117 ( .A1(o_cmd_forward_reg[17]), .A2(n48), .Z(n302)
         );
  CKAN2D1BWP30P140LVT U1118 ( .A1(o_cmd_forward_reg[11]), .A2(n48), .Z(n303)
         );
  CKAN2D1BWP30P140LVT U1119 ( .A1(o_cmd_forward_reg[6]), .A2(n48), .Z(n277) );
  AN4D1BWP30P140LVT U1120 ( .A1(n298), .A2(n46), .A3(o_cmd_forward_reg[42]), 
        .A4(o_valid_forward_reg[4]), .Z(n288) );
  AN4D1BWP30P140LVT U1121 ( .A1(n299), .A2(n47), .A3(o_cmd_forward_reg[27]), 
        .A4(o_valid_forward_reg[8]), .Z(n282) );
  AN4D1BWP30P140LVT U1122 ( .A1(n44), .A2(n302), .A3(o_cmd_forward_reg[19]), 
        .A4(o_valid_forward_reg[10]), .Z(n280) );
  AN4D1BWP30P140LVT U1123 ( .A1(n45), .A2(n303), .A3(o_cmd_forward_reg[10]), 
        .A4(o_valid_forward_reg[12]), .Z(n278) );
  AN4D1BWP30P140LVT U1124 ( .A1(n43), .A2(n277), .A3(o_cmd_forward_reg[7]), 
        .A4(o_valid_forward_reg[13]), .Z(n276) );
  ND2D1BWP30P140LVT U1125 ( .A1(o_cmd_forward_reg[2]), .A2(
        o_cmd_forward_reg[1]), .ZN(n26) );
  ND2D1BWP30P140LVT U1126 ( .A1(o_valid_forward_reg[14]), .A2(
        o_cmd_forward_reg[3]), .ZN(n25) );
  ND2D1BWP30P140LVT U1127 ( .A1(o_cmd_forward_reg[0]), .A2(n48), .ZN(n24) );
  NR2D1BWP30P140LVT U1128 ( .A1(n41), .A2(n18), .ZN(n284) );
  INVD1BWP30P140LVT U1129 ( .I(o_cmd_forward_reg[31]), .ZN(n41) );
  NR2D1BWP30P140LVT U1130 ( .A1(n35), .A2(n18), .ZN(n290) );
  INVD1BWP30P140LVT U1131 ( .I(o_cmd_forward_reg[46]), .ZN(n35) );
  NR2D1BWP30P140LVT U1132 ( .A1(n39), .A2(n49), .ZN(n293) );
  INVD1BWP30P140LVT U1133 ( .I(o_cmd_forward_reg[53]), .ZN(n39) );
  NR2D1BWP30P140LVT U1134 ( .A1(n37), .A2(n49), .ZN(n296) );
  INVD1BWP30P140LVT U1135 ( .I(o_cmd_forward_reg[56]), .ZN(n37) );
  INR2D1BWP30P140LVT U1136 ( .A1(i_valid), .B1(n49), .ZN(n295) );
  BUFFD2BWP30P140LVT U1137 ( .I(n285), .Z(n19) );
  INR3D0BWP30P140LVT U1138 ( .A1(o_valid_forward_reg[6]), .B1(
        o_cmd_forward_reg[35]), .B2(n30), .ZN(n285) );
  BUFFD2BWP30P140LVT U1139 ( .I(n279), .Z(n20) );
  INR3D0BWP30P140LVT U1140 ( .A1(o_valid_forward_reg[11]), .B1(
        o_cmd_forward_reg[12]), .B2(n33), .ZN(n279) );
  BUFFD2BWP30P140LVT U1141 ( .I(n281), .Z(n21) );
  INR3D0BWP30P140LVT U1142 ( .A1(o_valid_forward_reg[9]), .B1(
        o_cmd_forward_reg[20]), .B2(n34), .ZN(n281) );
  CKAN2D1BWP30P140LVT U1143 ( .A1(o_cmd_forward_reg[37]), .A2(n48), .Z(n287)
         );
  CKAN2D1BWP30P140LVT U1144 ( .A1(o_cmd_forward_reg[49]), .A2(n48), .Z(n297)
         );
  INVD1BWP30P140LVT U1145 ( .I(n49), .ZN(n48) );
  INVD1BWP30P140LVT U1146 ( .I(rst), .ZN(n23) );
  CKAN2D1BWP30P140LVT U1147 ( .A1(i_data_bus[27]), .A2(n48), .Z(n205) );
  CKAN2D1BWP30P140LVT U1148 ( .A1(i_data_bus[31]), .A2(n48), .Z(n209) );
  CKAN2D1BWP30P140LVT U1149 ( .A1(i_data_bus[25]), .A2(n48), .Z(n203) );
  CKAN2D1BWP30P140LVT U1150 ( .A1(i_data_bus[20]), .A2(n48), .Z(n198) );
  CKAN2D1BWP30P140LVT U1151 ( .A1(i_data_bus[12]), .A2(n48), .Z(n190) );
  CKAN2D1BWP30P140LVT U1152 ( .A1(i_data_bus[15]), .A2(n48), .Z(n193) );
  CKAN2D1BWP30P140LVT U1153 ( .A1(i_data_bus[14]), .A2(n48), .Z(n192) );
  CKAN2D1BWP30P140LVT U1154 ( .A1(i_data_bus[17]), .A2(n48), .Z(n195) );
  CKAN2D1BWP30P140LVT U1155 ( .A1(i_data_bus[11]), .A2(n48), .Z(n189) );
  CKAN2D1BWP30P140LVT U1156 ( .A1(i_data_bus[19]), .A2(n48), .Z(n197) );
  CKAN2D1BWP30P140LVT U1157 ( .A1(i_data_bus[16]), .A2(n48), .Z(n194) );
  CKAN2D1BWP30P140LVT U1158 ( .A1(i_data_bus[21]), .A2(n48), .Z(n199) );
  CKAN2D1BWP30P140LVT U1159 ( .A1(i_data_bus[22]), .A2(n48), .Z(n200) );
  CKAN2D1BWP30P140LVT U1160 ( .A1(i_data_bus[24]), .A2(n48), .Z(n202) );
  CKAN2D1BWP30P140LVT U1161 ( .A1(i_data_bus[13]), .A2(n48), .Z(n191) );
  CKAN2D1BWP30P140LVT U1162 ( .A1(i_data_bus[23]), .A2(n48), .Z(n201) );
  CKAN2D1BWP30P140LVT U1163 ( .A1(i_data_bus[18]), .A2(n48), .Z(n196) );
  CKAN2D1BWP30P140LVT U1164 ( .A1(i_data_bus[0]), .A2(n48), .Z(n178) );
  CKAN2D1BWP30P140LVT U1165 ( .A1(i_data_bus[8]), .A2(n48), .Z(n186) );
  CKAN2D1BWP30P140LVT U1166 ( .A1(i_data_bus[1]), .A2(n48), .Z(n179) );
  CKAN2D1BWP30P140LVT U1167 ( .A1(i_data_bus[4]), .A2(n48), .Z(n182) );
  CKAN2D1BWP30P140LVT U1168 ( .A1(i_data_bus[9]), .A2(n48), .Z(n187) );
  CKAN2D1BWP30P140LVT U1169 ( .A1(i_data_bus[6]), .A2(n48), .Z(n184) );
  CKAN2D1BWP30P140LVT U1170 ( .A1(i_data_bus[7]), .A2(n48), .Z(n185) );
  CKAN2D1BWP30P140LVT U1171 ( .A1(i_data_bus[3]), .A2(n48), .Z(n181) );
  CKAN2D1BWP30P140LVT U1172 ( .A1(i_data_bus[5]), .A2(n48), .Z(n183) );
  CKAN2D1BWP30P140LVT U1173 ( .A1(i_data_bus[10]), .A2(n48), .Z(n188) );
  CKAN2D1BWP30P140LVT U1174 ( .A1(i_data_bus[2]), .A2(n48), .Z(n180) );
  INR2D2BWP30P140LVT U1175 ( .A1(n29), .B1(n28), .ZN(n274) );
  ND3D1BWP30P140LVT U1176 ( .A1(n301), .A2(o_cmd_forward_reg[33]), .A3(
        o_cmd_forward_reg[32]), .ZN(n30) );
  IND3D1BWP30P140LVT U1177 ( .A1(o_cmd_forward_reg[51]), .B1(
        o_cmd_forward_reg[48]), .B2(n297), .ZN(n31) );
  INR3D2BWP30P140LVT U1178 ( .A1(o_valid_forward_reg[2]), .B1(
        o_cmd_forward_reg[50]), .B2(n31), .ZN(n291) );
  IND3D1BWP30P140LVT U1179 ( .A1(o_cmd_forward_reg[39]), .B1(
        o_valid_forward_reg[5]), .B2(n287), .ZN(n32) );
  INR3D2BWP30P140LVT U1180 ( .A1(o_cmd_forward_reg[38]), .B1(
        o_cmd_forward_reg[36]), .B2(n32), .ZN(n286) );
  IND3D1BWP30P140LVT U1181 ( .A1(o_cmd_forward_reg[13]), .B1(
        o_cmd_forward_reg[14]), .B2(n304), .ZN(n33) );
  IND3D1BWP30P140LVT U1182 ( .A1(o_cmd_forward_reg[22]), .B1(
        o_cmd_forward_reg[21]), .B2(n300), .ZN(n34) );
  IND2D1BWP30P140LVT U1183 ( .A1(o_cmd_forward_reg[44]), .B1(
        o_valid_forward_reg[3]), .ZN(n36) );
  INR4D2BWP30P140LVT U1184 ( .A1(n290), .B1(o_cmd_forward_reg[45]), .B2(
        o_cmd_forward_reg[47]), .B3(n36), .ZN(n289) );
  IND2D1BWP30P140LVT U1185 ( .A1(o_cmd_forward_reg[57]), .B1(
        o_valid_forward_reg[0]), .ZN(n38) );
  INR4D2BWP30P140LVT U1186 ( .A1(n296), .B1(o_cmd_forward_reg[58]), .B2(
        o_cmd_forward_reg[59]), .B3(n38), .ZN(n294) );
  IND2D1BWP30P140LVT U1187 ( .A1(o_cmd_forward_reg[52]), .B1(
        o_valid_forward_reg[1]), .ZN(n40) );
  INR4D2BWP30P140LVT U1188 ( .A1(n293), .B1(o_cmd_forward_reg[54]), .B2(
        o_cmd_forward_reg[55]), .B3(n40), .ZN(n292) );
  IND2D1BWP30P140LVT U1189 ( .A1(o_cmd_forward_reg[28]), .B1(
        o_valid_forward_reg[7]), .ZN(n42) );
  INR4D2BWP30P140LVT U1190 ( .A1(n284), .B1(o_cmd_forward_reg[29]), .B2(
        o_cmd_forward_reg[30]), .B3(n42), .ZN(n283) );
  INR2D1BWP30P140LVT U1191 ( .A1(o_cmd_forward_reg[5]), .B1(
        o_cmd_forward_reg[4]), .ZN(n43) );
  CKAN2D1BWP30P140LVT U1192 ( .A1(n276), .A2(o_data_forward_reg[45]), .Z(N2035) );
  CKAN2D1BWP30P140LVT U1193 ( .A1(n276), .A2(o_data_forward_reg[50]), .Z(N2040) );
  CKAN2D1BWP30P140LVT U1194 ( .A1(n276), .A2(o_data_forward_reg[48]), .Z(N2038) );
  CKAN2D1BWP30P140LVT U1195 ( .A1(n276), .A2(o_data_forward_reg[47]), .Z(N2037) );
  CKAN2D1BWP30P140LVT U1196 ( .A1(n276), .A2(o_data_forward_reg[42]), .Z(N2032) );
  CKAN2D1BWP30P140LVT U1197 ( .A1(n276), .A2(o_data_forward_reg[49]), .Z(N2039) );
  CKAN2D1BWP30P140LVT U1198 ( .A1(n276), .A2(o_data_forward_reg[44]), .Z(N2034) );
  CKAN2D1BWP30P140LVT U1199 ( .A1(n276), .A2(o_data_forward_reg[32]), .Z(N2022) );
  CKAN2D1BWP30P140LVT U1200 ( .A1(n276), .A2(o_data_forward_reg[59]), .Z(N2049) );
  CKAN2D1BWP30P140LVT U1201 ( .A1(n276), .A2(o_data_forward_reg[60]), .Z(N2050) );
  CKAN2D1BWP30P140LVT U1202 ( .A1(n276), .A2(o_data_forward_reg[46]), .Z(N2036) );
  CKAN2D1BWP30P140LVT U1203 ( .A1(n276), .A2(o_data_forward_reg[62]), .Z(N2052) );
  CKAN2D1BWP30P140LVT U1204 ( .A1(n276), .A2(o_data_forward_reg[33]), .Z(N2023) );
  CKAN2D1BWP30P140LVT U1205 ( .A1(n276), .A2(o_data_forward_reg[51]), .Z(N2041) );
  CKAN2D1BWP30P140LVT U1206 ( .A1(n276), .A2(o_data_forward_reg[52]), .Z(N2042) );
  CKAN2D1BWP30P140LVT U1207 ( .A1(n276), .A2(o_data_forward_reg[61]), .Z(N2051) );
  CKAN2D1BWP30P140LVT U1208 ( .A1(n276), .A2(o_data_forward_reg[54]), .Z(N2044) );
  CKAN2D1BWP30P140LVT U1209 ( .A1(n276), .A2(o_data_forward_reg[55]), .Z(N2045) );
  CKAN2D1BWP30P140LVT U1210 ( .A1(n276), .A2(o_data_forward_reg[39]), .Z(N2029) );
  CKAN2D1BWP30P140LVT U1211 ( .A1(n276), .A2(o_data_forward_reg[40]), .Z(N2030) );
  CKAN2D1BWP30P140LVT U1212 ( .A1(n276), .A2(o_data_forward_reg[41]), .Z(N2031) );
  CKAN2D1BWP30P140LVT U1213 ( .A1(n276), .A2(o_data_forward_reg[38]), .Z(N2028) );
  CKAN2D1BWP30P140LVT U1214 ( .A1(n276), .A2(o_data_forward_reg[43]), .Z(N2033) );
  CKAN2D1BWP30P140LVT U1215 ( .A1(n276), .A2(o_data_forward_reg[57]), .Z(N2047) );
  CKAN2D1BWP30P140LVT U1216 ( .A1(n276), .A2(o_data_forward_reg[58]), .Z(N2048) );
  CKAN2D1BWP30P140LVT U1217 ( .A1(n276), .A2(o_data_forward_reg[34]), .Z(N2024) );
  CKAN2D1BWP30P140LVT U1218 ( .A1(n276), .A2(o_data_forward_reg[35]), .Z(N2025) );
  CKAN2D1BWP30P140LVT U1219 ( .A1(n276), .A2(o_data_forward_reg[53]), .Z(N2043) );
  CKAN2D1BWP30P140LVT U1220 ( .A1(n276), .A2(o_data_forward_reg[37]), .Z(N2027) );
  CKAN2D1BWP30P140LVT U1221 ( .A1(n276), .A2(o_data_forward_reg[63]), .Z(N2053) );
  CKAN2D1BWP30P140LVT U1222 ( .A1(n276), .A2(o_data_forward_reg[56]), .Z(N2046) );
  CKAN2D1BWP30P140LVT U1223 ( .A1(n276), .A2(o_data_forward_reg[36]), .Z(N2026) );
  INR2D1BWP30P140LVT U1224 ( .A1(o_cmd_forward_reg[16]), .B1(
        o_cmd_forward_reg[18]), .ZN(n44) );
  CKAN2D1BWP30P140LVT U1225 ( .A1(n280), .A2(o_data_forward_reg[133]), .Z(
        N1619) );
  CKAN2D1BWP30P140LVT U1226 ( .A1(n280), .A2(o_data_forward_reg[132]), .Z(
        N1618) );
  CKAN2D1BWP30P140LVT U1227 ( .A1(n280), .A2(o_data_forward_reg[128]), .Z(
        N1614) );
  CKAN2D1BWP30P140LVT U1228 ( .A1(n280), .A2(o_data_forward_reg[134]), .Z(
        N1620) );
  CKAN2D1BWP30P140LVT U1229 ( .A1(n280), .A2(o_data_forward_reg[129]), .Z(
        N1615) );
  CKAN2D1BWP30P140LVT U1230 ( .A1(n280), .A2(o_data_forward_reg[130]), .Z(
        N1616) );
  CKAN2D1BWP30P140LVT U1231 ( .A1(n280), .A2(o_data_forward_reg[141]), .Z(
        N1627) );
  CKAN2D1BWP30P140LVT U1232 ( .A1(n280), .A2(o_data_forward_reg[142]), .Z(
        N1628) );
  CKAN2D1BWP30P140LVT U1233 ( .A1(n280), .A2(o_data_forward_reg[131]), .Z(
        N1617) );
  CKAN2D1BWP30P140LVT U1234 ( .A1(n280), .A2(o_data_forward_reg[144]), .Z(
        N1630) );
  CKAN2D1BWP30P140LVT U1235 ( .A1(n280), .A2(o_data_forward_reg[135]), .Z(
        N1621) );
  CKAN2D1BWP30P140LVT U1236 ( .A1(n280), .A2(o_data_forward_reg[136]), .Z(
        N1622) );
  CKAN2D1BWP30P140LVT U1237 ( .A1(n280), .A2(o_data_forward_reg[137]), .Z(
        N1623) );
  CKAN2D1BWP30P140LVT U1238 ( .A1(n280), .A2(o_data_forward_reg[143]), .Z(
        N1629) );
  CKAN2D1BWP30P140LVT U1239 ( .A1(n280), .A2(o_data_forward_reg[139]), .Z(
        N1625) );
  CKAN2D1BWP30P140LVT U1240 ( .A1(n280), .A2(o_data_forward_reg[140]), .Z(
        N1626) );
  CKAN2D1BWP30P140LVT U1241 ( .A1(n280), .A2(o_data_forward_reg[145]), .Z(
        N1631) );
  CKAN2D1BWP30P140LVT U1242 ( .A1(n280), .A2(o_data_forward_reg[146]), .Z(
        N1632) );
  CKAN2D1BWP30P140LVT U1243 ( .A1(n280), .A2(o_data_forward_reg[147]), .Z(
        N1633) );
  CKAN2D1BWP30P140LVT U1244 ( .A1(n280), .A2(o_data_forward_reg[148]), .Z(
        N1634) );
  CKAN2D1BWP30P140LVT U1245 ( .A1(n280), .A2(o_data_forward_reg[149]), .Z(
        N1635) );
  CKAN2D1BWP30P140LVT U1246 ( .A1(n280), .A2(o_data_forward_reg[150]), .Z(
        N1636) );
  CKAN2D1BWP30P140LVT U1247 ( .A1(n280), .A2(o_data_forward_reg[151]), .Z(
        N1637) );
  CKAN2D1BWP30P140LVT U1248 ( .A1(n280), .A2(o_data_forward_reg[152]), .Z(
        N1638) );
  CKAN2D1BWP30P140LVT U1249 ( .A1(n280), .A2(o_data_forward_reg[138]), .Z(
        N1624) );
  CKAN2D1BWP30P140LVT U1250 ( .A1(n280), .A2(o_data_forward_reg[153]), .Z(
        N1639) );
  CKAN2D1BWP30P140LVT U1251 ( .A1(n280), .A2(o_data_forward_reg[154]), .Z(
        N1640) );
  CKAN2D1BWP30P140LVT U1252 ( .A1(n280), .A2(o_data_forward_reg[155]), .Z(
        N1641) );
  CKAN2D1BWP30P140LVT U1253 ( .A1(n280), .A2(o_data_forward_reg[156]), .Z(
        N1642) );
  CKAN2D1BWP30P140LVT U1254 ( .A1(n280), .A2(o_data_forward_reg[157]), .Z(
        N1643) );
  CKAN2D1BWP30P140LVT U1255 ( .A1(n280), .A2(o_data_forward_reg[158]), .Z(
        N1644) );
  CKAN2D1BWP30P140LVT U1256 ( .A1(n280), .A2(o_data_forward_reg[159]), .Z(
        N1645) );
  INR2D1BWP30P140LVT U1257 ( .A1(o_cmd_forward_reg[8]), .B1(
        o_cmd_forward_reg[9]), .ZN(n45) );
  CKAN2D1BWP30P140LVT U1258 ( .A1(n278), .A2(o_data_forward_reg[64]), .Z(N1886) );
  CKAN2D1BWP30P140LVT U1259 ( .A1(n278), .A2(o_data_forward_reg[65]), .Z(N1887) );
  CKAN2D1BWP30P140LVT U1260 ( .A1(n278), .A2(o_data_forward_reg[66]), .Z(N1888) );
  CKAN2D1BWP30P140LVT U1261 ( .A1(n278), .A2(o_data_forward_reg[67]), .Z(N1889) );
  CKAN2D1BWP30P140LVT U1262 ( .A1(n278), .A2(o_data_forward_reg[68]), .Z(N1890) );
  CKAN2D1BWP30P140LVT U1263 ( .A1(n278), .A2(o_data_forward_reg[69]), .Z(N1891) );
  CKAN2D1BWP30P140LVT U1264 ( .A1(n278), .A2(o_data_forward_reg[70]), .Z(N1892) );
  CKAN2D1BWP30P140LVT U1265 ( .A1(n278), .A2(o_data_forward_reg[71]), .Z(N1893) );
  CKAN2D1BWP30P140LVT U1266 ( .A1(n278), .A2(o_data_forward_reg[72]), .Z(N1894) );
  CKAN2D1BWP30P140LVT U1267 ( .A1(n278), .A2(o_data_forward_reg[73]), .Z(N1895) );
  CKAN2D1BWP30P140LVT U1268 ( .A1(n278), .A2(o_data_forward_reg[74]), .Z(N1896) );
  CKAN2D1BWP30P140LVT U1269 ( .A1(n278), .A2(o_data_forward_reg[75]), .Z(N1897) );
  CKAN2D1BWP30P140LVT U1270 ( .A1(n278), .A2(o_data_forward_reg[76]), .Z(N1898) );
  CKAN2D1BWP30P140LVT U1271 ( .A1(n278), .A2(o_data_forward_reg[77]), .Z(N1899) );
  CKAN2D1BWP30P140LVT U1272 ( .A1(n278), .A2(o_data_forward_reg[78]), .Z(N1900) );
  CKAN2D1BWP30P140LVT U1273 ( .A1(n278), .A2(o_data_forward_reg[79]), .Z(N1901) );
  CKAN2D1BWP30P140LVT U1274 ( .A1(n278), .A2(o_data_forward_reg[80]), .Z(N1902) );
  CKAN2D1BWP30P140LVT U1275 ( .A1(n278), .A2(o_data_forward_reg[81]), .Z(N1903) );
  CKAN2D1BWP30P140LVT U1276 ( .A1(n278), .A2(o_data_forward_reg[82]), .Z(N1904) );
  CKAN2D1BWP30P140LVT U1277 ( .A1(n278), .A2(o_data_forward_reg[83]), .Z(N1905) );
  CKAN2D1BWP30P140LVT U1278 ( .A1(n278), .A2(o_data_forward_reg[84]), .Z(N1906) );
  CKAN2D1BWP30P140LVT U1279 ( .A1(n278), .A2(o_data_forward_reg[87]), .Z(N1909) );
  CKAN2D1BWP30P140LVT U1280 ( .A1(n278), .A2(o_data_forward_reg[88]), .Z(N1910) );
  CKAN2D1BWP30P140LVT U1281 ( .A1(n278), .A2(o_data_forward_reg[94]), .Z(N1916) );
  CKAN2D1BWP30P140LVT U1282 ( .A1(n278), .A2(o_data_forward_reg[89]), .Z(N1911) );
  CKAN2D1BWP30P140LVT U1283 ( .A1(n278), .A2(o_data_forward_reg[90]), .Z(N1912) );
  CKAN2D1BWP30P140LVT U1284 ( .A1(n278), .A2(o_data_forward_reg[91]), .Z(N1913) );
  CKAN2D1BWP30P140LVT U1285 ( .A1(n278), .A2(o_data_forward_reg[92]), .Z(N1914) );
  CKAN2D1BWP30P140LVT U1286 ( .A1(n278), .A2(o_data_forward_reg[93]), .Z(N1915) );
  CKAN2D1BWP30P140LVT U1287 ( .A1(n278), .A2(o_data_forward_reg[95]), .Z(N1917) );
  CKAN2D1BWP30P140LVT U1288 ( .A1(n278), .A2(o_data_forward_reg[86]), .Z(N1908) );
  CKAN2D1BWP30P140LVT U1289 ( .A1(n278), .A2(o_data_forward_reg[85]), .Z(N1907) );
  CKAN2D1BWP30P140LVT U1290 ( .A1(n288), .A2(o_data_forward_reg[322]), .Z(N800) );
  CKAN2D1BWP30P140LVT U1291 ( .A1(n288), .A2(o_data_forward_reg[332]), .Z(N810) );
  CKAN2D1BWP30P140LVT U1292 ( .A1(n288), .A2(o_data_forward_reg[334]), .Z(N812) );
  CKAN2D1BWP30P140LVT U1293 ( .A1(n288), .A2(o_data_forward_reg[335]), .Z(N813) );
  CKAN2D1BWP30P140LVT U1294 ( .A1(n288), .A2(o_data_forward_reg[336]), .Z(N814) );
  CKAN2D1BWP30P140LVT U1295 ( .A1(n288), .A2(o_data_forward_reg[331]), .Z(N809) );
  CKAN2D1BWP30P140LVT U1296 ( .A1(n288), .A2(o_data_forward_reg[338]), .Z(N816) );
  CKAN2D1BWP30P140LVT U1297 ( .A1(n288), .A2(o_data_forward_reg[333]), .Z(N811) );
  CKAN2D1BWP30P140LVT U1298 ( .A1(n288), .A2(o_data_forward_reg[339]), .Z(N817) );
  CKAN2D1BWP30P140LVT U1299 ( .A1(n288), .A2(o_data_forward_reg[340]), .Z(N818) );
  CKAN2D1BWP30P140LVT U1300 ( .A1(n288), .A2(o_data_forward_reg[341]), .Z(N819) );
  CKAN2D1BWP30P140LVT U1301 ( .A1(n288), .A2(o_data_forward_reg[343]), .Z(N821) );
  CKAN2D1BWP30P140LVT U1302 ( .A1(n288), .A2(o_data_forward_reg[344]), .Z(N822) );
  CKAN2D1BWP30P140LVT U1303 ( .A1(n288), .A2(o_data_forward_reg[345]), .Z(N823) );
  CKAN2D1BWP30P140LVT U1304 ( .A1(n288), .A2(o_data_forward_reg[346]), .Z(N824) );
  CKAN2D1BWP30P140LVT U1305 ( .A1(n288), .A2(o_data_forward_reg[347]), .Z(N825) );
  CKAN2D1BWP30P140LVT U1306 ( .A1(n288), .A2(o_data_forward_reg[348]), .Z(N826) );
  CKAN2D1BWP30P140LVT U1307 ( .A1(n288), .A2(o_data_forward_reg[349]), .Z(N827) );
  CKAN2D1BWP30P140LVT U1308 ( .A1(n288), .A2(o_data_forward_reg[350]), .Z(N828) );
  CKAN2D1BWP30P140LVT U1309 ( .A1(n288), .A2(o_data_forward_reg[337]), .Z(N815) );
  CKAN2D1BWP30P140LVT U1310 ( .A1(n288), .A2(o_data_forward_reg[320]), .Z(N798) );
  CKAN2D1BWP30P140LVT U1311 ( .A1(n288), .A2(o_data_forward_reg[321]), .Z(N799) );
  CKAN2D1BWP30P140LVT U1312 ( .A1(n288), .A2(o_data_forward_reg[351]), .Z(N829) );
  CKAN2D1BWP30P140LVT U1313 ( .A1(n288), .A2(o_data_forward_reg[323]), .Z(N801) );
  CKAN2D1BWP30P140LVT U1314 ( .A1(n288), .A2(o_data_forward_reg[324]), .Z(N802) );
  CKAN2D1BWP30P140LVT U1315 ( .A1(n288), .A2(o_data_forward_reg[325]), .Z(N803) );
  CKAN2D1BWP30P140LVT U1316 ( .A1(n288), .A2(o_data_forward_reg[326]), .Z(N804) );
  CKAN2D1BWP30P140LVT U1317 ( .A1(n288), .A2(o_data_forward_reg[327]), .Z(N805) );
  CKAN2D1BWP30P140LVT U1318 ( .A1(n288), .A2(o_data_forward_reg[328]), .Z(N806) );
  CKAN2D1BWP30P140LVT U1319 ( .A1(n288), .A2(o_data_forward_reg[329]), .Z(N807) );
  CKAN2D1BWP30P140LVT U1320 ( .A1(n288), .A2(o_data_forward_reg[330]), .Z(N808) );
  CKAN2D1BWP30P140LVT U1321 ( .A1(n288), .A2(o_data_forward_reg[342]), .Z(N820) );
  CKAN2D1BWP30P140LVT U1322 ( .A1(n282), .A2(o_data_forward_reg[214]), .Z(
        N1364) );
  CKAN2D1BWP30P140LVT U1323 ( .A1(n282), .A2(o_data_forward_reg[213]), .Z(
        N1363) );
  CKAN2D1BWP30P140LVT U1324 ( .A1(n282), .A2(o_data_forward_reg[212]), .Z(
        N1362) );
  CKAN2D1BWP30P140LVT U1325 ( .A1(n282), .A2(o_data_forward_reg[211]), .Z(
        N1361) );
  CKAN2D1BWP30P140LVT U1326 ( .A1(n282), .A2(o_data_forward_reg[210]), .Z(
        N1360) );
  CKAN2D1BWP30P140LVT U1327 ( .A1(n282), .A2(o_data_forward_reg[209]), .Z(
        N1359) );
  CKAN2D1BWP30P140LVT U1328 ( .A1(n282), .A2(o_data_forward_reg[208]), .Z(
        N1358) );
  CKAN2D1BWP30P140LVT U1329 ( .A1(n282), .A2(o_data_forward_reg[207]), .Z(
        N1357) );
  CKAN2D1BWP30P140LVT U1330 ( .A1(n282), .A2(o_data_forward_reg[206]), .Z(
        N1356) );
  CKAN2D1BWP30P140LVT U1331 ( .A1(n282), .A2(o_data_forward_reg[205]), .Z(
        N1355) );
  CKAN2D1BWP30P140LVT U1332 ( .A1(n282), .A2(o_data_forward_reg[204]), .Z(
        N1354) );
  CKAN2D1BWP30P140LVT U1333 ( .A1(n282), .A2(o_data_forward_reg[203]), .Z(
        N1353) );
  CKAN2D1BWP30P140LVT U1334 ( .A1(n282), .A2(o_data_forward_reg[202]), .Z(
        N1352) );
  CKAN2D1BWP30P140LVT U1335 ( .A1(n282), .A2(o_data_forward_reg[201]), .Z(
        N1351) );
  CKAN2D1BWP30P140LVT U1336 ( .A1(n282), .A2(o_data_forward_reg[200]), .Z(
        N1350) );
  CKAN2D1BWP30P140LVT U1337 ( .A1(n282), .A2(o_data_forward_reg[199]), .Z(
        N1349) );
  CKAN2D1BWP30P140LVT U1338 ( .A1(n282), .A2(o_data_forward_reg[198]), .Z(
        N1348) );
  CKAN2D1BWP30P140LVT U1339 ( .A1(n282), .A2(o_data_forward_reg[197]), .Z(
        N1347) );
  CKAN2D1BWP30P140LVT U1340 ( .A1(n282), .A2(o_data_forward_reg[196]), .Z(
        N1346) );
  CKAN2D1BWP30P140LVT U1341 ( .A1(n282), .A2(o_data_forward_reg[195]), .Z(
        N1345) );
  CKAN2D1BWP30P140LVT U1342 ( .A1(n282), .A2(o_data_forward_reg[194]), .Z(
        N1344) );
  CKAN2D1BWP30P140LVT U1343 ( .A1(n282), .A2(o_data_forward_reg[193]), .Z(
        N1343) );
  CKAN2D1BWP30P140LVT U1344 ( .A1(n282), .A2(o_data_forward_reg[192]), .Z(
        N1342) );
  CKAN2D1BWP30P140LVT U1345 ( .A1(n282), .A2(o_data_forward_reg[222]), .Z(
        N1372) );
  CKAN2D1BWP30P140LVT U1346 ( .A1(n282), .A2(o_data_forward_reg[219]), .Z(
        N1369) );
  CKAN2D1BWP30P140LVT U1347 ( .A1(n282), .A2(o_data_forward_reg[215]), .Z(
        N1365) );
  CKAN2D1BWP30P140LVT U1348 ( .A1(n282), .A2(o_data_forward_reg[216]), .Z(
        N1366) );
  CKAN2D1BWP30P140LVT U1349 ( .A1(n282), .A2(o_data_forward_reg[217]), .Z(
        N1367) );
  CKAN2D1BWP30P140LVT U1350 ( .A1(n282), .A2(o_data_forward_reg[218]), .Z(
        N1368) );
  CKAN2D1BWP30P140LVT U1351 ( .A1(n282), .A2(o_data_forward_reg[220]), .Z(
        N1370) );
  CKAN2D1BWP30P140LVT U1352 ( .A1(n282), .A2(o_data_forward_reg[221]), .Z(
        N1371) );
  CKAN2D1BWP30P140LVT U1353 ( .A1(n282), .A2(o_data_forward_reg[223]), .Z(
        N1373) );
  INR2D1BWP30P140LVT U1354 ( .A1(o_data_forward_reg[390]), .B1(n18), .ZN(N564)
         );
  INR2D1BWP30P140LVT U1355 ( .A1(o_data_forward_reg[479]), .B1(n18), .ZN(N317)
         );
  INR2D1BWP30P140LVT U1356 ( .A1(o_data_forward_reg[389]), .B1(n18), .ZN(N563)
         );
  INR2D1BWP30P140LVT U1357 ( .A1(o_data_forward_reg[394]), .B1(n18), .ZN(N568)
         );
  INR2D1BWP30P140LVT U1358 ( .A1(o_data_forward_reg[395]), .B1(n18), .ZN(N569)
         );
  INR2D1BWP30P140LVT U1359 ( .A1(o_data_forward_reg[396]), .B1(n18), .ZN(N570)
         );
  INR2D1BWP30P140LVT U1360 ( .A1(o_data_forward_reg[397]), .B1(n49), .ZN(N571)
         );
  INR2D1BWP30P140LVT U1361 ( .A1(o_data_forward_reg[398]), .B1(n49), .ZN(N572)
         );
  INR2D1BWP30P140LVT U1362 ( .A1(o_data_forward_reg[399]), .B1(n49), .ZN(N573)
         );
  INR2D1BWP30P140LVT U1363 ( .A1(o_data_forward_reg[400]), .B1(n18), .ZN(N574)
         );
  INR2D1BWP30P140LVT U1364 ( .A1(o_data_forward_reg[393]), .B1(n18), .ZN(N567)
         );
  INR2D1BWP30P140LVT U1365 ( .A1(o_data_forward_reg[416]), .B1(n18), .ZN(N422)
         );
  INR2D1BWP30P140LVT U1366 ( .A1(o_data_forward_reg[417]), .B1(n49), .ZN(N423)
         );
  INR2D1BWP30P140LVT U1367 ( .A1(o_data_forward_reg[418]), .B1(n49), .ZN(N424)
         );
  INR2D1BWP30P140LVT U1368 ( .A1(o_data_forward_reg[419]), .B1(n18), .ZN(N425)
         );
  INR2D1BWP30P140LVT U1369 ( .A1(o_data_forward_reg[420]), .B1(n18), .ZN(N426)
         );
  INR2D1BWP30P140LVT U1370 ( .A1(o_data_forward_reg[391]), .B1(n18), .ZN(N565)
         );
  INR2D1BWP30P140LVT U1371 ( .A1(o_data_forward_reg[422]), .B1(n18), .ZN(N428)
         );
  INR2D1BWP30P140LVT U1372 ( .A1(o_data_forward_reg[423]), .B1(n18), .ZN(N429)
         );
  INR2D1BWP30P140LVT U1373 ( .A1(o_data_forward_reg[392]), .B1(n49), .ZN(N566)
         );
  INR2D1BWP30P140LVT U1374 ( .A1(o_data_forward_reg[425]), .B1(n18), .ZN(N431)
         );
  INR2D1BWP30P140LVT U1375 ( .A1(o_data_forward_reg[426]), .B1(n18), .ZN(N432)
         );
  INR2D1BWP30P140LVT U1376 ( .A1(o_data_forward_reg[427]), .B1(n49), .ZN(N433)
         );
  INR2D1BWP30P140LVT U1377 ( .A1(o_data_forward_reg[421]), .B1(n18), .ZN(N427)
         );
  INR2D1BWP30P140LVT U1378 ( .A1(o_data_forward_reg[401]), .B1(n18), .ZN(N575)
         );
  INR2D1BWP30P140LVT U1379 ( .A1(o_data_forward_reg[424]), .B1(n49), .ZN(N430)
         );
  INR2D1BWP30P140LVT U1380 ( .A1(o_data_forward_reg[429]), .B1(n18), .ZN(N435)
         );
  INR2D1BWP30P140LVT U1381 ( .A1(o_data_forward_reg[432]), .B1(n49), .ZN(N438)
         );
  INR2D1BWP30P140LVT U1382 ( .A1(o_data_forward_reg[430]), .B1(n18), .ZN(N436)
         );
  INR2D1BWP30P140LVT U1383 ( .A1(o_data_forward_reg[428]), .B1(n18), .ZN(N434)
         );
  INR2D1BWP30P140LVT U1384 ( .A1(o_data_forward_reg[435]), .B1(n18), .ZN(N441)
         );
  INR2D1BWP30P140LVT U1385 ( .A1(o_data_forward_reg[436]), .B1(n49), .ZN(N442)
         );
  INR2D1BWP30P140LVT U1386 ( .A1(o_data_forward_reg[437]), .B1(n18), .ZN(N443)
         );
  INR2D1BWP30P140LVT U1387 ( .A1(o_data_forward_reg[438]), .B1(n18), .ZN(N444)
         );
  INR2D1BWP30P140LVT U1388 ( .A1(o_data_forward_reg[431]), .B1(n18), .ZN(N437)
         );
  INR2D1BWP30P140LVT U1389 ( .A1(o_data_forward_reg[439]), .B1(n49), .ZN(N445)
         );
  INR2D1BWP30P140LVT U1390 ( .A1(o_data_forward_reg[440]), .B1(n18), .ZN(N446)
         );
  INR2D1BWP30P140LVT U1391 ( .A1(o_data_forward_reg[434]), .B1(n18), .ZN(N440)
         );
  INR2D1BWP30P140LVT U1392 ( .A1(o_data_forward_reg[433]), .B1(n18), .ZN(N439)
         );
  INR2D1BWP30P140LVT U1393 ( .A1(o_data_forward_reg[465]), .B1(n18), .ZN(N303)
         );
  INR2D1BWP30P140LVT U1394 ( .A1(o_data_forward_reg[453]), .B1(n18), .ZN(N291)
         );
  INR2D1BWP30P140LVT U1395 ( .A1(o_data_forward_reg[454]), .B1(n49), .ZN(N292)
         );
  INR2D1BWP30P140LVT U1396 ( .A1(o_data_forward_reg[455]), .B1(n18), .ZN(N293)
         );
  INR2D1BWP30P140LVT U1397 ( .A1(o_data_forward_reg[456]), .B1(n18), .ZN(N294)
         );
  INR2D1BWP30P140LVT U1398 ( .A1(o_data_forward_reg[457]), .B1(n18), .ZN(N295)
         );
  INR2D1BWP30P140LVT U1399 ( .A1(o_data_forward_reg[458]), .B1(n18), .ZN(N296)
         );
  INR2D1BWP30P140LVT U1400 ( .A1(o_data_forward_reg[459]), .B1(n49), .ZN(N297)
         );
  INR2D1BWP30P140LVT U1401 ( .A1(o_data_forward_reg[460]), .B1(n18), .ZN(N298)
         );
  INR2D1BWP30P140LVT U1402 ( .A1(o_data_forward_reg[461]), .B1(n49), .ZN(N299)
         );
  INR2D1BWP30P140LVT U1403 ( .A1(o_data_forward_reg[462]), .B1(n18), .ZN(N300)
         );
  INR2D1BWP30P140LVT U1404 ( .A1(o_data_forward_reg[463]), .B1(n18), .ZN(N301)
         );
  INR2D1BWP30P140LVT U1405 ( .A1(o_data_forward_reg[464]), .B1(n49), .ZN(N302)
         );
  INR2D1BWP30P140LVT U1406 ( .A1(o_data_forward_reg[332]), .B1(n18), .ZN(N842)
         );
  INR2D1BWP30P140LVT U1407 ( .A1(o_data_forward_reg[335]), .B1(n49), .ZN(N845)
         );
  INR2D1BWP30P140LVT U1408 ( .A1(o_data_forward_reg[336]), .B1(n18), .ZN(N846)
         );
  INR2D1BWP30P140LVT U1409 ( .A1(o_data_forward_reg[334]), .B1(n18), .ZN(N844)
         );
  INR2D1BWP30P140LVT U1410 ( .A1(o_data_forward_reg[337]), .B1(n18), .ZN(N847)
         );
  INR2D1BWP30P140LVT U1411 ( .A1(o_data_forward_reg[412]), .B1(n18), .ZN(N586)
         );
  INR2D1BWP30P140LVT U1412 ( .A1(o_data_forward_reg[411]), .B1(n49), .ZN(N585)
         );
  INR2D1BWP30P140LVT U1413 ( .A1(o_data_forward_reg[410]), .B1(n18), .ZN(N584)
         );
  INR2D1BWP30P140LVT U1414 ( .A1(o_data_forward_reg[409]), .B1(n49), .ZN(N583)
         );
  INR2D1BWP30P140LVT U1415 ( .A1(o_data_forward_reg[408]), .B1(n18), .ZN(N582)
         );
  INR2D1BWP30P140LVT U1416 ( .A1(o_data_forward_reg[407]), .B1(n18), .ZN(N581)
         );
  INR2D1BWP30P140LVT U1417 ( .A1(o_data_forward_reg[406]), .B1(n18), .ZN(N580)
         );
  INR2D1BWP30P140LVT U1418 ( .A1(o_data_forward_reg[405]), .B1(n18), .ZN(N579)
         );
  INR2D1BWP30P140LVT U1419 ( .A1(o_data_forward_reg[404]), .B1(n18), .ZN(N578)
         );
  INR2D1BWP30P140LVT U1420 ( .A1(o_data_forward_reg[328]), .B1(n49), .ZN(N838)
         );
  INR2D1BWP30P140LVT U1421 ( .A1(o_data_forward_reg[414]), .B1(n18), .ZN(N588)
         );
  INR2D1BWP30P140LVT U1422 ( .A1(o_data_forward_reg[333]), .B1(n18), .ZN(N843)
         );
  INR2D1BWP30P140LVT U1423 ( .A1(o_data_forward_reg[330]), .B1(n18), .ZN(N840)
         );
  INR2D1BWP30P140LVT U1424 ( .A1(o_data_forward_reg[329]), .B1(n18), .ZN(N839)
         );
  INR2D1BWP30P140LVT U1425 ( .A1(o_data_forward_reg[327]), .B1(n18), .ZN(N837)
         );
  INR2D1BWP30P140LVT U1426 ( .A1(o_data_forward_reg[326]), .B1(n18), .ZN(N836)
         );
  INR2D1BWP30P140LVT U1427 ( .A1(o_data_forward_reg[413]), .B1(n18), .ZN(N587)
         );
  INR2D1BWP30P140LVT U1428 ( .A1(o_data_forward_reg[325]), .B1(n18), .ZN(N835)
         );
  INR2D1BWP30P140LVT U1429 ( .A1(o_data_forward_reg[331]), .B1(n18), .ZN(N841)
         );
  INR2D1BWP30P140LVT U1430 ( .A1(o_data_forward_reg[403]), .B1(n49), .ZN(N577)
         );
  INR2D1BWP30P140LVT U1431 ( .A1(o_data_forward_reg[402]), .B1(n18), .ZN(N576)
         );
  INR2D1BWP30P140LVT U1432 ( .A1(o_data_forward_reg[363]), .B1(n18), .ZN(N705)
         );
  INR2D1BWP30P140LVT U1433 ( .A1(o_data_forward_reg[359]), .B1(n49), .ZN(N701)
         );
  INR2D1BWP30P140LVT U1434 ( .A1(o_data_forward_reg[355]), .B1(n18), .ZN(N697)
         );
  INR2D1BWP30P140LVT U1435 ( .A1(o_data_forward_reg[352]), .B1(n18), .ZN(N694)
         );
  INR2D1BWP30P140LVT U1436 ( .A1(o_data_forward_reg[356]), .B1(n18), .ZN(N698)
         );
  INR2D1BWP30P140LVT U1437 ( .A1(o_data_forward_reg[358]), .B1(n18), .ZN(N700)
         );
  INR2D1BWP30P140LVT U1438 ( .A1(o_data_forward_reg[354]), .B1(n18), .ZN(N696)
         );
  INR2D1BWP30P140LVT U1439 ( .A1(o_data_forward_reg[353]), .B1(n18), .ZN(N695)
         );
  INR2D1BWP30P140LVT U1440 ( .A1(o_data_forward_reg[360]), .B1(n49), .ZN(N702)
         );
  INR2D1BWP30P140LVT U1441 ( .A1(o_data_forward_reg[415]), .B1(n18), .ZN(N589)
         );
  INR2D1BWP30P140LVT U1442 ( .A1(o_data_forward_reg[361]), .B1(n49), .ZN(N703)
         );
  INR2D1BWP30P140LVT U1443 ( .A1(o_data_forward_reg[357]), .B1(n49), .ZN(N699)
         );
  INR2D1BWP30P140LVT U1444 ( .A1(o_data_forward_reg[362]), .B1(n18), .ZN(N704)
         );
  INR2D1BWP30P140LVT U1445 ( .A1(o_data_forward_reg[343]), .B1(n18), .ZN(N853)
         );
  INR2D1BWP30P140LVT U1446 ( .A1(o_data_forward_reg[347]), .B1(n49), .ZN(N857)
         );
  INR2D1BWP30P140LVT U1447 ( .A1(o_data_forward_reg[342]), .B1(n49), .ZN(N852)
         );
  INR2D1BWP30P140LVT U1448 ( .A1(o_data_forward_reg[348]), .B1(n18), .ZN(N858)
         );
  INR2D1BWP30P140LVT U1449 ( .A1(o_data_forward_reg[349]), .B1(n49), .ZN(N859)
         );
  INR2D1BWP30P140LVT U1450 ( .A1(o_data_forward_reg[344]), .B1(n18), .ZN(N854)
         );
  INR2D1BWP30P140LVT U1451 ( .A1(o_data_forward_reg[345]), .B1(n18), .ZN(N855)
         );
  INR2D1BWP30P140LVT U1452 ( .A1(o_data_forward_reg[346]), .B1(n18), .ZN(N856)
         );
  INR2D1BWP30P140LVT U1453 ( .A1(o_data_forward_reg[339]), .B1(n49), .ZN(N849)
         );
  INR2D1BWP30P140LVT U1454 ( .A1(o_data_forward_reg[340]), .B1(n18), .ZN(N850)
         );
  INR2D1BWP30P140LVT U1455 ( .A1(o_data_forward_reg[341]), .B1(n18), .ZN(N851)
         );
  INR2D1BWP30P140LVT U1456 ( .A1(o_data_forward_reg[338]), .B1(n49), .ZN(N848)
         );
  INR2D1BWP30P140LVT U1457 ( .A1(o_data_forward_reg[191]), .B1(n18), .ZN(N1541) );
  INR2D1BWP30P140LVT U1458 ( .A1(o_data_forward_reg[350]), .B1(n18), .ZN(N860)
         );
  INR2D1BWP30P140LVT U1459 ( .A1(o_data_forward_reg[128]), .B1(n49), .ZN(N1646) );
  INR2D1BWP30P140LVT U1460 ( .A1(o_data_forward_reg[129]), .B1(n49), .ZN(N1647) );
  INR2D1BWP30P140LVT U1461 ( .A1(o_data_forward_reg[299]), .B1(n49), .ZN(N977)
         );
  INR2D1BWP30P140LVT U1462 ( .A1(o_data_forward_reg[298]), .B1(n49), .ZN(N976)
         );
  INR2D1BWP30P140LVT U1463 ( .A1(o_data_forward_reg[297]), .B1(n49), .ZN(N975)
         );
  INR2D1BWP30P140LVT U1464 ( .A1(o_data_forward_reg[296]), .B1(n18), .ZN(N974)
         );
  INR2D1BWP30P140LVT U1465 ( .A1(o_data_forward_reg[295]), .B1(n18), .ZN(N973)
         );
  INR2D1BWP30P140LVT U1466 ( .A1(o_data_forward_reg[294]), .B1(n18), .ZN(N972)
         );
  INR2D1BWP30P140LVT U1467 ( .A1(o_data_forward_reg[293]), .B1(n18), .ZN(N971)
         );
  INR2D1BWP30P140LVT U1468 ( .A1(o_data_forward_reg[291]), .B1(n18), .ZN(N969)
         );
  INR2D1BWP30P140LVT U1469 ( .A1(o_data_forward_reg[290]), .B1(n18), .ZN(N968)
         );
  INR2D1BWP30P140LVT U1470 ( .A1(o_data_forward_reg[289]), .B1(n18), .ZN(N967)
         );
  INR2D1BWP30P140LVT U1471 ( .A1(o_data_forward_reg[288]), .B1(n18), .ZN(N966)
         );
  INR2D1BWP30P140LVT U1472 ( .A1(o_data_forward_reg[130]), .B1(n18), .ZN(N1648) );
  INR2D1BWP30P140LVT U1473 ( .A1(o_data_forward_reg[131]), .B1(n18), .ZN(N1649) );
  INR2D1BWP30P140LVT U1474 ( .A1(o_data_forward_reg[132]), .B1(n18), .ZN(N1650) );
  INR2D1BWP30P140LVT U1475 ( .A1(o_data_forward_reg[133]), .B1(n18), .ZN(N1651) );
  INR2D1BWP30P140LVT U1476 ( .A1(o_data_forward_reg[134]), .B1(n18), .ZN(N1652) );
  INR2D1BWP30P140LVT U1477 ( .A1(o_data_forward_reg[173]), .B1(n18), .ZN(N1523) );
  INR2D1BWP30P140LVT U1478 ( .A1(o_data_forward_reg[174]), .B1(n18), .ZN(N1524) );
  INR2D1BWP30P140LVT U1479 ( .A1(o_data_forward_reg[175]), .B1(n18), .ZN(N1525) );
  INR2D1BWP30P140LVT U1480 ( .A1(o_data_forward_reg[176]), .B1(n18), .ZN(N1526) );
  INR2D1BWP30P140LVT U1481 ( .A1(o_data_forward_reg[177]), .B1(n18), .ZN(N1527) );
  INR2D1BWP30P140LVT U1482 ( .A1(o_data_forward_reg[178]), .B1(n18), .ZN(N1528) );
  INR2D1BWP30P140LVT U1483 ( .A1(o_data_forward_reg[179]), .B1(n49), .ZN(N1529) );
  INR2D1BWP30P140LVT U1484 ( .A1(o_data_forward_reg[180]), .B1(n18), .ZN(N1530) );
  INR2D1BWP30P140LVT U1485 ( .A1(o_data_forward_reg[181]), .B1(n18), .ZN(N1531) );
  INR2D1BWP30P140LVT U1486 ( .A1(o_data_forward_reg[182]), .B1(n18), .ZN(N1532) );
  INR2D1BWP30P140LVT U1487 ( .A1(o_data_forward_reg[183]), .B1(n18), .ZN(N1533) );
  INR2D1BWP30P140LVT U1488 ( .A1(o_data_forward_reg[184]), .B1(n18), .ZN(N1534) );
  INR2D1BWP30P140LVT U1489 ( .A1(o_data_forward_reg[185]), .B1(n18), .ZN(N1535) );
  INR2D1BWP30P140LVT U1490 ( .A1(o_data_forward_reg[186]), .B1(n49), .ZN(N1536) );
  INR2D1BWP30P140LVT U1491 ( .A1(o_data_forward_reg[187]), .B1(n18), .ZN(N1537) );
  INR2D1BWP30P140LVT U1492 ( .A1(o_data_forward_reg[188]), .B1(n18), .ZN(N1538) );
  INR2D1BWP30P140LVT U1493 ( .A1(o_data_forward_reg[189]), .B1(n49), .ZN(N1539) );
  INR2D1BWP30P140LVT U1494 ( .A1(o_data_forward_reg[190]), .B1(n18), .ZN(N1540) );
  INR2D1BWP30P140LVT U1495 ( .A1(o_data_forward_reg[292]), .B1(n18), .ZN(N970)
         );
  INR2D1BWP30P140LVT U1496 ( .A1(o_data_forward_reg[351]), .B1(n18), .ZN(N861)
         );
  INR2D1BWP30P140LVT U1497 ( .A1(o_data_forward_reg[100]), .B1(n18), .ZN(N1786) );
  INR2D1BWP30P140LVT U1498 ( .A1(o_data_forward_reg[99]), .B1(n18), .ZN(N1785)
         );
  INR2D1BWP30P140LVT U1499 ( .A1(o_data_forward_reg[98]), .B1(n18), .ZN(N1784)
         );
  INR2D1BWP30P140LVT U1500 ( .A1(o_data_forward_reg[97]), .B1(n18), .ZN(N1783)
         );
  INR2D1BWP30P140LVT U1501 ( .A1(o_data_forward_reg[95]), .B1(n18), .ZN(N1949)
         );
  INR2D1BWP30P140LVT U1502 ( .A1(o_data_forward_reg[94]), .B1(n18), .ZN(N1948)
         );
  INR2D1BWP30P140LVT U1503 ( .A1(o_data_forward_reg[93]), .B1(n18), .ZN(N1947)
         );
  INR2D1BWP30P140LVT U1504 ( .A1(o_data_forward_reg[92]), .B1(n18), .ZN(N1946)
         );
  INR2D1BWP30P140LVT U1505 ( .A1(o_data_forward_reg[91]), .B1(n18), .ZN(N1945)
         );
  INR2D1BWP30P140LVT U1506 ( .A1(o_data_forward_reg[90]), .B1(n49), .ZN(N1944)
         );
  INR2D1BWP30P140LVT U1507 ( .A1(o_data_forward_reg[89]), .B1(n18), .ZN(N1943)
         );
  INR2D1BWP30P140LVT U1508 ( .A1(o_data_forward_reg[88]), .B1(n18), .ZN(N1942)
         );
  INR2D1BWP30P140LVT U1509 ( .A1(o_data_forward_reg[87]), .B1(n49), .ZN(N1941)
         );
  INR2D1BWP30P140LVT U1510 ( .A1(o_data_forward_reg[86]), .B1(n49), .ZN(N1940)
         );
  INR2D1BWP30P140LVT U1511 ( .A1(o_data_forward_reg[85]), .B1(n49), .ZN(N1939)
         );
  INR2D1BWP30P140LVT U1512 ( .A1(o_data_forward_reg[84]), .B1(n49), .ZN(N1938)
         );
  INR2D1BWP30P140LVT U1513 ( .A1(o_data_forward_reg[83]), .B1(n49), .ZN(N1937)
         );
  INR2D1BWP30P140LVT U1514 ( .A1(o_data_forward_reg[82]), .B1(n18), .ZN(N1936)
         );
  INR2D1BWP30P140LVT U1515 ( .A1(o_data_forward_reg[81]), .B1(n18), .ZN(N1935)
         );
  INR2D1BWP30P140LVT U1516 ( .A1(o_data_forward_reg[80]), .B1(n49), .ZN(N1934)
         );
  INR2D1BWP30P140LVT U1517 ( .A1(o_data_forward_reg[79]), .B1(n49), .ZN(N1933)
         );
  INR2D1BWP30P140LVT U1518 ( .A1(o_data_forward_reg[78]), .B1(n18), .ZN(N1932)
         );
  INR2D1BWP30P140LVT U1519 ( .A1(o_data_forward_reg[77]), .B1(n18), .ZN(N1931)
         );
  INR2D1BWP30P140LVT U1520 ( .A1(o_data_forward_reg[76]), .B1(n18), .ZN(N1930)
         );
  INR2D1BWP30P140LVT U1521 ( .A1(o_data_forward_reg[101]), .B1(n18), .ZN(N1787) );
  INR2D1BWP30P140LVT U1522 ( .A1(o_data_forward_reg[102]), .B1(n18), .ZN(N1788) );
  INR2D1BWP30P140LVT U1523 ( .A1(o_data_forward_reg[103]), .B1(n18), .ZN(N1789) );
  INR2D1BWP30P140LVT U1524 ( .A1(o_data_forward_reg[104]), .B1(n18), .ZN(N1790) );
  INR2D1BWP30P140LVT U1525 ( .A1(o_data_forward_reg[105]), .B1(n49), .ZN(N1791) );
  INR2D1BWP30P140LVT U1526 ( .A1(o_data_forward_reg[106]), .B1(n18), .ZN(N1792) );
  INR2D1BWP30P140LVT U1527 ( .A1(o_data_forward_reg[107]), .B1(n18), .ZN(N1793) );
  INR2D1BWP30P140LVT U1528 ( .A1(o_data_forward_reg[108]), .B1(n18), .ZN(N1794) );
  INR2D1BWP30P140LVT U1529 ( .A1(o_data_forward_reg[109]), .B1(n49), .ZN(N1795) );
  INR2D1BWP30P140LVT U1530 ( .A1(o_data_forward_reg[110]), .B1(n18), .ZN(N1796) );
  INR2D1BWP30P140LVT U1531 ( .A1(o_data_forward_reg[111]), .B1(n49), .ZN(N1797) );
  INR2D1BWP30P140LVT U1532 ( .A1(o_data_forward_reg[112]), .B1(n18), .ZN(N1798) );
  INR2D1BWP30P140LVT U1533 ( .A1(o_data_forward_reg[113]), .B1(n18), .ZN(N1799) );
  INR2D1BWP30P140LVT U1534 ( .A1(o_data_forward_reg[114]), .B1(n18), .ZN(N1800) );
  INR2D1BWP30P140LVT U1535 ( .A1(o_data_forward_reg[115]), .B1(n18), .ZN(N1801) );
  INR2D1BWP30P140LVT U1536 ( .A1(o_data_forward_reg[116]), .B1(n18), .ZN(N1802) );
  INR2D1BWP30P140LVT U1537 ( .A1(o_data_forward_reg[117]), .B1(n18), .ZN(N1803) );
  INR2D1BWP30P140LVT U1538 ( .A1(o_data_forward_reg[118]), .B1(n18), .ZN(N1804) );
  INR2D1BWP30P140LVT U1539 ( .A1(o_data_forward_reg[119]), .B1(n18), .ZN(N1805) );
  INR2D1BWP30P140LVT U1540 ( .A1(o_data_forward_reg[120]), .B1(n18), .ZN(N1806) );
  INR2D1BWP30P140LVT U1541 ( .A1(o_data_forward_reg[121]), .B1(n49), .ZN(N1807) );
  INR2D1BWP30P140LVT U1542 ( .A1(o_data_forward_reg[122]), .B1(n18), .ZN(N1808) );
  INR2D1BWP30P140LVT U1543 ( .A1(o_data_forward_reg[123]), .B1(n18), .ZN(N1809) );
  INR2D1BWP30P140LVT U1544 ( .A1(o_data_forward_reg[124]), .B1(n18), .ZN(N1810) );
  INR2D1BWP30P140LVT U1545 ( .A1(o_data_forward_reg[125]), .B1(n49), .ZN(N1811) );
  INR2D1BWP30P140LVT U1546 ( .A1(o_data_forward_reg[126]), .B1(n18), .ZN(N1812) );
  INR2D1BWP30P140LVT U1547 ( .A1(o_data_forward_reg[127]), .B1(n18), .ZN(N1813) );
  INR2D1BWP30P140LVT U1548 ( .A1(o_data_forward_reg[75]), .B1(n49), .ZN(N1929)
         );
  INR2D1BWP30P140LVT U1549 ( .A1(o_data_forward_reg[74]), .B1(n18), .ZN(N1928)
         );
  INR2D1BWP30P140LVT U1550 ( .A1(o_data_forward_reg[73]), .B1(n18), .ZN(N1927)
         );
  INR2D1BWP30P140LVT U1551 ( .A1(o_data_forward_reg[72]), .B1(n18), .ZN(N1926)
         );
  INR2D1BWP30P140LVT U1552 ( .A1(o_data_forward_reg[71]), .B1(n18), .ZN(N1925)
         );
  INR2D1BWP30P140LVT U1553 ( .A1(o_data_forward_reg[70]), .B1(n49), .ZN(N1924)
         );
  INR2D1BWP30P140LVT U1554 ( .A1(o_data_forward_reg[69]), .B1(n18), .ZN(N1923)
         );
  INR2D1BWP30P140LVT U1555 ( .A1(o_data_forward_reg[68]), .B1(n49), .ZN(N1922)
         );
  INR2D1BWP30P140LVT U1556 ( .A1(o_data_forward_reg[67]), .B1(n18), .ZN(N1921)
         );
  INR2D1BWP30P140LVT U1557 ( .A1(o_data_forward_reg[66]), .B1(n49), .ZN(N1920)
         );
  INR2D1BWP30P140LVT U1558 ( .A1(o_data_forward_reg[65]), .B1(n18), .ZN(N1919)
         );
  INR2D1BWP30P140LVT U1559 ( .A1(o_data_forward_reg[64]), .B1(n18), .ZN(N1918)
         );
  INR2D1BWP30P140LVT U1560 ( .A1(o_data_forward_reg[58]), .B1(n18), .ZN(N2080)
         );
  INR2D1BWP30P140LVT U1561 ( .A1(o_data_forward_reg[57]), .B1(n49), .ZN(N2079)
         );
  INR2D1BWP30P140LVT U1562 ( .A1(o_data_forward_reg[56]), .B1(n18), .ZN(N2078)
         );
  INR2D1BWP30P140LVT U1563 ( .A1(o_data_forward_reg[55]), .B1(n18), .ZN(N2077)
         );
  INR2D1BWP30P140LVT U1564 ( .A1(o_data_forward_reg[54]), .B1(n49), .ZN(N2076)
         );
  INR2D1BWP30P140LVT U1565 ( .A1(o_data_forward_reg[53]), .B1(n18), .ZN(N2075)
         );
  INR2D1BWP30P140LVT U1566 ( .A1(o_data_forward_reg[52]), .B1(n18), .ZN(N2074)
         );
  INR2D1BWP30P140LVT U1567 ( .A1(o_data_forward_reg[51]), .B1(n18), .ZN(N2073)
         );
  INR2D1BWP30P140LVT U1568 ( .A1(o_data_forward_reg[50]), .B1(n18), .ZN(N2072)
         );
  INR2D1BWP30P140LVT U1569 ( .A1(o_data_forward_reg[49]), .B1(n49), .ZN(N2071)
         );
  INR2D1BWP30P140LVT U1570 ( .A1(o_data_forward_reg[48]), .B1(n18), .ZN(N2070)
         );
  INR2D1BWP30P140LVT U1571 ( .A1(o_data_forward_reg[47]), .B1(n18), .ZN(N2069)
         );
  INR2D1BWP30P140LVT U1572 ( .A1(o_data_forward_reg[46]), .B1(n49), .ZN(N2068)
         );
  INR2D1BWP30P140LVT U1573 ( .A1(o_data_forward_reg[45]), .B1(n18), .ZN(N2067)
         );
  INR2D1BWP30P140LVT U1574 ( .A1(o_data_forward_reg[44]), .B1(n18), .ZN(N2066)
         );
  INR2D1BWP30P140LVT U1575 ( .A1(o_data_forward_reg[43]), .B1(n18), .ZN(N2065)
         );
  INR2D1BWP30P140LVT U1576 ( .A1(o_data_forward_reg[42]), .B1(n18), .ZN(N2064)
         );
  INR2D1BWP30P140LVT U1577 ( .A1(o_data_forward_reg[41]), .B1(n18), .ZN(N2063)
         );
  INR2D1BWP30P140LVT U1578 ( .A1(o_data_forward_reg[40]), .B1(n18), .ZN(N2062)
         );
  INR2D1BWP30P140LVT U1579 ( .A1(o_data_forward_reg[39]), .B1(n18), .ZN(N2061)
         );
  INR2D1BWP30P140LVT U1580 ( .A1(o_data_forward_reg[38]), .B1(n18), .ZN(N2060)
         );
  INR2D1BWP30P140LVT U1581 ( .A1(o_data_forward_reg[37]), .B1(n18), .ZN(N2059)
         );
  INR2D1BWP30P140LVT U1582 ( .A1(o_data_forward_reg[36]), .B1(n49), .ZN(N2058)
         );
  INR2D1BWP30P140LVT U1583 ( .A1(o_data_forward_reg[35]), .B1(n49), .ZN(N2057)
         );
  INR2D1BWP30P140LVT U1584 ( .A1(o_data_forward_reg[34]), .B1(n18), .ZN(N2056)
         );
  INR2D1BWP30P140LVT U1585 ( .A1(o_data_forward_reg[33]), .B1(n18), .ZN(N2055)
         );
  INR2D1BWP30P140LVT U1586 ( .A1(o_data_forward_reg[32]), .B1(n18), .ZN(N2054)
         );
  INR2D1BWP30P140LVT U1587 ( .A1(o_cmd_forward_reg[59]), .B1(n18), .ZN(N322)
         );
  INR2D1BWP30P140LVT U1588 ( .A1(o_cmd_forward_reg[55]), .B1(n18), .ZN(N458)
         );
  INR2D1BWP30P140LVT U1589 ( .A1(o_cmd_forward_reg[45]), .B1(n18), .ZN(N728)
         );
  INR2D1BWP30P140LVT U1590 ( .A1(o_cmd_forward_reg[47]), .B1(n18), .ZN(N730)
         );
  INR2D1BWP30P140LVT U1591 ( .A1(o_data_forward_reg[324]), .B1(n18), .ZN(N834)
         );
  INR2D1BWP30P140LVT U1592 ( .A1(o_data_forward_reg[381]), .B1(n18), .ZN(N723)
         );
  INR2D1BWP30P140LVT U1593 ( .A1(o_data_forward_reg[323]), .B1(n18), .ZN(N833)
         );
  INR2D1BWP30P140LVT U1594 ( .A1(o_data_forward_reg[378]), .B1(n18), .ZN(N720)
         );
  INR2D1BWP30P140LVT U1595 ( .A1(o_data_forward_reg[377]), .B1(n18), .ZN(N719)
         );
  INR2D1BWP30P140LVT U1596 ( .A1(o_data_forward_reg[382]), .B1(n18), .ZN(N724)
         );
  INR2D1BWP30P140LVT U1597 ( .A1(o_data_forward_reg[383]), .B1(n18), .ZN(N725)
         );
  INR2D1BWP30P140LVT U1598 ( .A1(o_data_forward_reg[379]), .B1(n18), .ZN(N721)
         );
  INR2D1BWP30P140LVT U1599 ( .A1(o_data_forward_reg[321]), .B1(n18), .ZN(N831)
         );
  INR2D1BWP30P140LVT U1600 ( .A1(o_data_forward_reg[322]), .B1(n18), .ZN(N832)
         );
  INR2D1BWP30P140LVT U1601 ( .A1(o_data_forward_reg[380]), .B1(n18), .ZN(N722)
         );
  INR2D1BWP30P140LVT U1602 ( .A1(o_data_forward_reg[320]), .B1(n18), .ZN(N830)
         );
  INR2D1BWP30P140LVT U1603 ( .A1(o_data_forward_reg[475]), .B1(n18), .ZN(N313)
         );
  INR2D1BWP30P140LVT U1604 ( .A1(o_data_forward_reg[468]), .B1(n18), .ZN(N306)
         );
  INR2D1BWP30P140LVT U1605 ( .A1(o_data_forward_reg[477]), .B1(n18), .ZN(N315)
         );
  INR2D1BWP30P140LVT U1606 ( .A1(o_data_forward_reg[470]), .B1(n18), .ZN(N308)
         );
  INR2D1BWP30P140LVT U1607 ( .A1(o_data_forward_reg[474]), .B1(n18), .ZN(N312)
         );
  INR2D1BWP30P140LVT U1608 ( .A1(o_data_forward_reg[466]), .B1(n18), .ZN(N304)
         );
  INR2D1BWP30P140LVT U1609 ( .A1(o_data_forward_reg[478]), .B1(n18), .ZN(N316)
         );
  INR2D1BWP30P140LVT U1610 ( .A1(o_data_forward_reg[476]), .B1(n18), .ZN(N314)
         );
  INR2D1BWP30P140LVT U1611 ( .A1(o_data_forward_reg[472]), .B1(n18), .ZN(N310)
         );
  INR2D1BWP30P140LVT U1612 ( .A1(o_data_forward_reg[467]), .B1(n18), .ZN(N305)
         );
  INR2D1BWP30P140LVT U1613 ( .A1(o_data_forward_reg[473]), .B1(n18), .ZN(N311)
         );
  INR2D1BWP30P140LVT U1614 ( .A1(o_data_forward_reg[471]), .B1(n18), .ZN(N309)
         );
  INR2D1BWP30P140LVT U1615 ( .A1(o_data_forward_reg[469]), .B1(n18), .ZN(N307)
         );
  INR2D1BWP30P140LVT U1616 ( .A1(o_cmd_forward_reg[51]), .B1(n18), .ZN(N594)
         );
  INR2D1BWP30P140LVT U1617 ( .A1(o_data_forward_reg[386]), .B1(n18), .ZN(N560)
         );
  INR2D1BWP30P140LVT U1618 ( .A1(o_data_forward_reg[447]), .B1(n18), .ZN(N453)
         );
  INR2D1BWP30P140LVT U1619 ( .A1(o_data_forward_reg[444]), .B1(n18), .ZN(N450)
         );
  INR2D1BWP30P140LVT U1620 ( .A1(o_data_forward_reg[384]), .B1(n18), .ZN(N558)
         );
  INR2D1BWP30P140LVT U1621 ( .A1(o_data_forward_reg[443]), .B1(n18), .ZN(N449)
         );
  INR2D1BWP30P140LVT U1622 ( .A1(o_data_forward_reg[445]), .B1(n18), .ZN(N451)
         );
  INR2D1BWP30P140LVT U1623 ( .A1(o_data_forward_reg[387]), .B1(n18), .ZN(N561)
         );
  INR2D1BWP30P140LVT U1624 ( .A1(o_data_forward_reg[385]), .B1(n49), .ZN(N559)
         );
  INR2D1BWP30P140LVT U1625 ( .A1(o_data_forward_reg[442]), .B1(n49), .ZN(N448)
         );
  INR2D1BWP30P140LVT U1626 ( .A1(o_data_forward_reg[441]), .B1(n18), .ZN(N447)
         );
  INR2D1BWP30P140LVT U1627 ( .A1(o_data_forward_reg[446]), .B1(n18), .ZN(N452)
         );
  INR2D1BWP30P140LVT U1628 ( .A1(o_data_forward_reg[388]), .B1(n18), .ZN(N562)
         );
  INR2D1BWP30P140LVT U1629 ( .A1(o_data_forward_reg[448]), .B1(n49), .ZN(N286)
         );
  INR2D1BWP30P140LVT U1630 ( .A1(o_data_forward_reg[449]), .B1(n49), .ZN(N287)
         );
  INR2D1BWP30P140LVT U1631 ( .A1(o_data_forward_reg[450]), .B1(n49), .ZN(N288)
         );
  INR2D1BWP30P140LVT U1632 ( .A1(o_data_forward_reg[452]), .B1(n49), .ZN(N290)
         );
  INR2D1BWP30P140LVT U1633 ( .A1(o_data_forward_reg[451]), .B1(n49), .ZN(N289)
         );
  INR2D1BWP30P140LVT U1634 ( .A1(o_data_forward_reg[156]), .B1(n49), .ZN(N1674) );
  INR2D1BWP30P140LVT U1635 ( .A1(o_data_forward_reg[157]), .B1(n49), .ZN(N1675) );
  INR2D1BWP30P140LVT U1636 ( .A1(o_data_forward_reg[148]), .B1(n18), .ZN(N1666) );
  INR2D1BWP30P140LVT U1637 ( .A1(o_data_forward_reg[149]), .B1(n18), .ZN(N1667) );
  INR2D1BWP30P140LVT U1638 ( .A1(o_data_forward_reg[158]), .B1(n18), .ZN(N1676) );
  INR2D1BWP30P140LVT U1639 ( .A1(o_data_forward_reg[159]), .B1(n18), .ZN(N1677) );
  INR2D1BWP30P140LVT U1640 ( .A1(o_data_forward_reg[151]), .B1(n18), .ZN(N1669) );
  INR2D1BWP30P140LVT U1641 ( .A1(o_data_forward_reg[154]), .B1(n18), .ZN(N1672) );
  INR2D1BWP30P140LVT U1642 ( .A1(o_data_forward_reg[155]), .B1(n18), .ZN(N1673) );
  INR2D1BWP30P140LVT U1643 ( .A1(o_data_forward_reg[152]), .B1(n49), .ZN(N1670) );
  INR2D1BWP30P140LVT U1644 ( .A1(o_data_forward_reg[153]), .B1(n18), .ZN(N1671) );
  INR2D1BWP30P140LVT U1645 ( .A1(o_data_forward_reg[96]), .B1(n49), .ZN(N1782)
         );
  INR2D1BWP30P140LVT U1646 ( .A1(o_data_forward_reg[150]), .B1(n18), .ZN(N1668) );
  INR2D1BWP30P140LVT U1647 ( .A1(o_data_forward_reg[365]), .B1(n18), .ZN(N707)
         );
  INR2D1BWP30P140LVT U1648 ( .A1(o_data_forward_reg[366]), .B1(n18), .ZN(N708)
         );
  INR2D1BWP30P140LVT U1649 ( .A1(o_data_forward_reg[367]), .B1(n18), .ZN(N709)
         );
  INR2D1BWP30P140LVT U1650 ( .A1(o_data_forward_reg[368]), .B1(n18), .ZN(N710)
         );
  INR2D1BWP30P140LVT U1651 ( .A1(o_data_forward_reg[369]), .B1(n18), .ZN(N711)
         );
  INR2D1BWP30P140LVT U1652 ( .A1(o_data_forward_reg[370]), .B1(n18), .ZN(N712)
         );
  INR2D1BWP30P140LVT U1653 ( .A1(o_data_forward_reg[373]), .B1(n18), .ZN(N715)
         );
  INR2D1BWP30P140LVT U1654 ( .A1(o_data_forward_reg[376]), .B1(n18), .ZN(N718)
         );
  INR2D1BWP30P140LVT U1655 ( .A1(o_data_forward_reg[374]), .B1(n18), .ZN(N716)
         );
  INR2D1BWP30P140LVT U1656 ( .A1(o_data_forward_reg[364]), .B1(n18), .ZN(N706)
         );
  INR2D1BWP30P140LVT U1657 ( .A1(o_data_forward_reg[372]), .B1(n18), .ZN(N714)
         );
  INR2D1BWP30P140LVT U1658 ( .A1(o_data_forward_reg[375]), .B1(n18), .ZN(N717)
         );
  INR2D1BWP30P140LVT U1659 ( .A1(o_data_forward_reg[371]), .B1(n18), .ZN(N713)
         );
  INR2D1BWP30P140LVT U1660 ( .A1(o_cmd_forward_reg[29]), .B1(n49), .ZN(N1272)
         );
  INR2D1BWP30P140LVT U1661 ( .A1(o_data_forward_reg[318]), .B1(n18), .ZN(N996)
         );
  INR2D1BWP30P140LVT U1662 ( .A1(o_data_forward_reg[317]), .B1(n18), .ZN(N995)
         );
  INR2D1BWP30P140LVT U1663 ( .A1(o_data_forward_reg[165]), .B1(n18), .ZN(N1515) );
  INR2D1BWP30P140LVT U1664 ( .A1(o_data_forward_reg[162]), .B1(n18), .ZN(N1512) );
  INR2D1BWP30P140LVT U1665 ( .A1(o_data_forward_reg[163]), .B1(n18), .ZN(N1513) );
  INR2D1BWP30P140LVT U1666 ( .A1(o_data_forward_reg[160]), .B1(n18), .ZN(N1510) );
  INR2D1BWP30P140LVT U1667 ( .A1(o_data_forward_reg[161]), .B1(n18), .ZN(N1511) );
  INR2D1BWP30P140LVT U1668 ( .A1(o_data_forward_reg[315]), .B1(n18), .ZN(N993)
         );
  INR2D1BWP30P140LVT U1669 ( .A1(o_data_forward_reg[314]), .B1(n49), .ZN(N992)
         );
  INR2D1BWP30P140LVT U1670 ( .A1(o_data_forward_reg[313]), .B1(n18), .ZN(N991)
         );
  INR2D1BWP30P140LVT U1671 ( .A1(o_data_forward_reg[166]), .B1(n18), .ZN(N1516) );
  INR2D1BWP30P140LVT U1672 ( .A1(o_data_forward_reg[256]), .B1(n18), .ZN(N1102) );
  INR2D1BWP30P140LVT U1673 ( .A1(o_data_forward_reg[164]), .B1(n18), .ZN(N1514) );
  INR2D1BWP30P140LVT U1674 ( .A1(o_data_forward_reg[258]), .B1(n18), .ZN(N1104) );
  INR2D1BWP30P140LVT U1675 ( .A1(o_data_forward_reg[259]), .B1(n18), .ZN(N1105) );
  INR2D1BWP30P140LVT U1676 ( .A1(o_data_forward_reg[260]), .B1(n18), .ZN(N1106) );
  INR2D1BWP30P140LVT U1677 ( .A1(o_data_forward_reg[257]), .B1(n18), .ZN(N1103) );
  INR2D1BWP30P140LVT U1678 ( .A1(o_data_forward_reg[316]), .B1(n49), .ZN(N994)
         );
  INR2D1BWP30P140LVT U1679 ( .A1(o_data_forward_reg[319]), .B1(n18), .ZN(N997)
         );
  INR2D1BWP30P140LVT U1680 ( .A1(o_data_forward_reg[172]), .B1(n49), .ZN(N1522) );
  INR2D1BWP30P140LVT U1681 ( .A1(o_data_forward_reg[171]), .B1(n18), .ZN(N1521) );
  INR2D1BWP30P140LVT U1682 ( .A1(o_data_forward_reg[170]), .B1(n18), .ZN(N1520) );
  INR2D1BWP30P140LVT U1683 ( .A1(o_data_forward_reg[169]), .B1(n18), .ZN(N1519) );
  INR2D1BWP30P140LVT U1684 ( .A1(o_data_forward_reg[168]), .B1(n18), .ZN(N1518) );
  INR2D1BWP30P140LVT U1685 ( .A1(o_data_forward_reg[167]), .B1(n18), .ZN(N1517) );
  INR2D1BWP30P140LVT U1686 ( .A1(o_data_forward_reg[312]), .B1(n18), .ZN(N990)
         );
  INR2D1BWP30P140LVT U1687 ( .A1(o_data_forward_reg[311]), .B1(n18), .ZN(N989)
         );
  INR2D1BWP30P140LVT U1688 ( .A1(o_data_forward_reg[284]), .B1(n49), .ZN(N1130) );
  INR2D1BWP30P140LVT U1689 ( .A1(o_data_forward_reg[309]), .B1(n49), .ZN(N987)
         );
  INR2D1BWP30P140LVT U1690 ( .A1(o_data_forward_reg[308]), .B1(n49), .ZN(N986)
         );
  INR2D1BWP30P140LVT U1691 ( .A1(o_data_forward_reg[307]), .B1(n49), .ZN(N985)
         );
  INR2D1BWP30P140LVT U1692 ( .A1(o_data_forward_reg[306]), .B1(n49), .ZN(N984)
         );
  INR2D1BWP30P140LVT U1693 ( .A1(o_data_forward_reg[305]), .B1(n18), .ZN(N983)
         );
  INR2D1BWP30P140LVT U1694 ( .A1(o_data_forward_reg[304]), .B1(n18), .ZN(N982)
         );
  INR2D1BWP30P140LVT U1695 ( .A1(o_data_forward_reg[303]), .B1(n18), .ZN(N981)
         );
  INR2D1BWP30P140LVT U1696 ( .A1(o_data_forward_reg[302]), .B1(n49), .ZN(N980)
         );
  INR2D1BWP30P140LVT U1697 ( .A1(o_data_forward_reg[301]), .B1(n18), .ZN(N979)
         );
  INR2D1BWP30P140LVT U1698 ( .A1(o_data_forward_reg[300]), .B1(n18), .ZN(N978)
         );
  INR2D1BWP30P140LVT U1699 ( .A1(o_data_forward_reg[310]), .B1(n18), .ZN(N988)
         );
  INR2D1BWP30P140LVT U1700 ( .A1(o_data_forward_reg[287]), .B1(n18), .ZN(N1133) );
  INR2D1BWP30P140LVT U1701 ( .A1(o_data_forward_reg[286]), .B1(n18), .ZN(N1132) );
  INR2D1BWP30P140LVT U1702 ( .A1(o_data_forward_reg[285]), .B1(n18), .ZN(N1131) );
  INR2D1BWP30P140LVT U1703 ( .A1(o_data_forward_reg[263]), .B1(n18), .ZN(N1109) );
  INR2D1BWP30P140LVT U1704 ( .A1(o_data_forward_reg[210]), .B1(n18), .ZN(N1392) );
  INR2D1BWP30P140LVT U1705 ( .A1(o_data_forward_reg[261]), .B1(n18), .ZN(N1107) );
  INR2D1BWP30P140LVT U1706 ( .A1(o_data_forward_reg[264]), .B1(n18), .ZN(N1110) );
  INR2D1BWP30P140LVT U1707 ( .A1(o_data_forward_reg[255]), .B1(n18), .ZN(N1269) );
  INR2D1BWP30P140LVT U1708 ( .A1(o_data_forward_reg[254]), .B1(n18), .ZN(N1268) );
  INR2D1BWP30P140LVT U1709 ( .A1(o_data_forward_reg[253]), .B1(n18), .ZN(N1267) );
  INR2D1BWP30P140LVT U1710 ( .A1(o_data_forward_reg[252]), .B1(n18), .ZN(N1266) );
  INR2D1BWP30P140LVT U1711 ( .A1(o_data_forward_reg[251]), .B1(n18), .ZN(N1265) );
  INR2D1BWP30P140LVT U1712 ( .A1(o_data_forward_reg[250]), .B1(n49), .ZN(N1264) );
  INR2D1BWP30P140LVT U1713 ( .A1(o_data_forward_reg[249]), .B1(n18), .ZN(N1263) );
  INR2D1BWP30P140LVT U1714 ( .A1(o_data_forward_reg[248]), .B1(n49), .ZN(N1262) );
  INR2D1BWP30P140LVT U1715 ( .A1(o_data_forward_reg[262]), .B1(n18), .ZN(N1108) );
  INR2D1BWP30P140LVT U1716 ( .A1(o_data_forward_reg[246]), .B1(n49), .ZN(N1260) );
  INR2D1BWP30P140LVT U1717 ( .A1(o_data_forward_reg[245]), .B1(n18), .ZN(N1259) );
  INR2D1BWP30P140LVT U1718 ( .A1(o_data_forward_reg[244]), .B1(n18), .ZN(N1258) );
  INR2D1BWP30P140LVT U1719 ( .A1(o_data_forward_reg[243]), .B1(n49), .ZN(N1257) );
  INR2D1BWP30P140LVT U1720 ( .A1(o_data_forward_reg[242]), .B1(n49), .ZN(N1256) );
  INR2D1BWP30P140LVT U1721 ( .A1(o_data_forward_reg[241]), .B1(n49), .ZN(N1255) );
  INR2D1BWP30P140LVT U1722 ( .A1(o_data_forward_reg[240]), .B1(n18), .ZN(N1254) );
  INR2D1BWP30P140LVT U1723 ( .A1(o_data_forward_reg[239]), .B1(n18), .ZN(N1253) );
  INR2D1BWP30P140LVT U1724 ( .A1(o_data_forward_reg[238]), .B1(n18), .ZN(N1252) );
  INR2D1BWP30P140LVT U1725 ( .A1(o_data_forward_reg[237]), .B1(n49), .ZN(N1251) );
  INR2D1BWP30P140LVT U1726 ( .A1(o_data_forward_reg[236]), .B1(n18), .ZN(N1250) );
  INR2D1BWP30P140LVT U1727 ( .A1(o_data_forward_reg[235]), .B1(n18), .ZN(N1249) );
  INR2D1BWP30P140LVT U1728 ( .A1(o_data_forward_reg[234]), .B1(n18), .ZN(N1248) );
  INR2D1BWP30P140LVT U1729 ( .A1(o_data_forward_reg[233]), .B1(n18), .ZN(N1247) );
  INR2D1BWP30P140LVT U1730 ( .A1(o_data_forward_reg[232]), .B1(n18), .ZN(N1246) );
  INR2D1BWP30P140LVT U1731 ( .A1(o_data_forward_reg[231]), .B1(n18), .ZN(N1245) );
  INR2D1BWP30P140LVT U1732 ( .A1(o_data_forward_reg[230]), .B1(n18), .ZN(N1244) );
  INR2D1BWP30P140LVT U1733 ( .A1(o_data_forward_reg[229]), .B1(n49), .ZN(N1243) );
  INR2D1BWP30P140LVT U1734 ( .A1(o_data_forward_reg[228]), .B1(n18), .ZN(N1242) );
  INR2D1BWP30P140LVT U1735 ( .A1(o_data_forward_reg[227]), .B1(n18), .ZN(N1241) );
  INR2D1BWP30P140LVT U1736 ( .A1(o_data_forward_reg[226]), .B1(n18), .ZN(N1240) );
  INR2D1BWP30P140LVT U1737 ( .A1(o_data_forward_reg[225]), .B1(n18), .ZN(N1239) );
  INR2D1BWP30P140LVT U1738 ( .A1(o_data_forward_reg[224]), .B1(n18), .ZN(N1238) );
  INR2D1BWP30P140LVT U1739 ( .A1(o_data_forward_reg[223]), .B1(n18), .ZN(N1405) );
  INR2D1BWP30P140LVT U1740 ( .A1(o_data_forward_reg[222]), .B1(n18), .ZN(N1404) );
  INR2D1BWP30P140LVT U1741 ( .A1(o_data_forward_reg[221]), .B1(n49), .ZN(N1403) );
  INR2D1BWP30P140LVT U1742 ( .A1(o_data_forward_reg[220]), .B1(n49), .ZN(N1402) );
  INR2D1BWP30P140LVT U1743 ( .A1(o_data_forward_reg[219]), .B1(n49), .ZN(N1401) );
  INR2D1BWP30P140LVT U1744 ( .A1(o_data_forward_reg[218]), .B1(n18), .ZN(N1400) );
  INR2D1BWP30P140LVT U1745 ( .A1(o_data_forward_reg[217]), .B1(n18), .ZN(N1399) );
  INR2D1BWP30P140LVT U1746 ( .A1(o_data_forward_reg[216]), .B1(n18), .ZN(N1398) );
  INR2D1BWP30P140LVT U1747 ( .A1(o_data_forward_reg[215]), .B1(n18), .ZN(N1397) );
  INR2D1BWP30P140LVT U1748 ( .A1(o_data_forward_reg[214]), .B1(n18), .ZN(N1396) );
  INR2D1BWP30P140LVT U1749 ( .A1(o_data_forward_reg[213]), .B1(n49), .ZN(N1395) );
  INR2D1BWP30P140LVT U1750 ( .A1(o_data_forward_reg[212]), .B1(n18), .ZN(N1394) );
  INR2D1BWP30P140LVT U1751 ( .A1(o_data_forward_reg[211]), .B1(n18), .ZN(N1393) );
  INR2D1BWP30P140LVT U1752 ( .A1(o_data_forward_reg[209]), .B1(n18), .ZN(N1391) );
  INR2D1BWP30P140LVT U1753 ( .A1(o_data_forward_reg[208]), .B1(n18), .ZN(N1390) );
  INR2D1BWP30P140LVT U1754 ( .A1(o_data_forward_reg[207]), .B1(n18), .ZN(N1389) );
  INR2D1BWP30P140LVT U1755 ( .A1(o_data_forward_reg[206]), .B1(n18), .ZN(N1388) );
  INR2D1BWP30P140LVT U1756 ( .A1(o_data_forward_reg[205]), .B1(n18), .ZN(N1387) );
  INR2D1BWP30P140LVT U1757 ( .A1(o_data_forward_reg[247]), .B1(n49), .ZN(N1261) );
  INR2D1BWP30P140LVT U1758 ( .A1(o_data_forward_reg[273]), .B1(n49), .ZN(N1119) );
  INR2D1BWP30P140LVT U1759 ( .A1(o_data_forward_reg[196]), .B1(n18), .ZN(N1378) );
  INR2D1BWP30P140LVT U1760 ( .A1(o_data_forward_reg[204]), .B1(n18), .ZN(N1386) );
  INR2D1BWP30P140LVT U1761 ( .A1(o_data_forward_reg[203]), .B1(n49), .ZN(N1385) );
  INR2D1BWP30P140LVT U1762 ( .A1(o_data_forward_reg[202]), .B1(n18), .ZN(N1384) );
  INR2D1BWP30P140LVT U1763 ( .A1(o_data_forward_reg[192]), .B1(n49), .ZN(N1374) );
  INR2D1BWP30P140LVT U1764 ( .A1(o_data_forward_reg[201]), .B1(n49), .ZN(N1383) );
  INR2D1BWP30P140LVT U1765 ( .A1(o_data_forward_reg[200]), .B1(n18), .ZN(N1382) );
  INR2D1BWP30P140LVT U1766 ( .A1(o_data_forward_reg[199]), .B1(n49), .ZN(N1381) );
  INR2D1BWP30P140LVT U1767 ( .A1(o_data_forward_reg[281]), .B1(n18), .ZN(N1127) );
  INR2D1BWP30P140LVT U1768 ( .A1(o_data_forward_reg[267]), .B1(n18), .ZN(N1113) );
  INR2D1BWP30P140LVT U1769 ( .A1(o_data_forward_reg[198]), .B1(n18), .ZN(N1380) );
  INR2D1BWP30P140LVT U1770 ( .A1(o_data_forward_reg[193]), .B1(n18), .ZN(N1375) );
  INR2D1BWP30P140LVT U1771 ( .A1(o_data_forward_reg[197]), .B1(n49), .ZN(N1379) );
  INR2D1BWP30P140LVT U1772 ( .A1(o_data_forward_reg[270]), .B1(n18), .ZN(N1116) );
  INR2D1BWP30P140LVT U1773 ( .A1(o_data_forward_reg[195]), .B1(n18), .ZN(N1377) );
  INR2D1BWP30P140LVT U1774 ( .A1(o_data_forward_reg[194]), .B1(n18), .ZN(N1376) );
  INR2D1BWP30P140LVT U1775 ( .A1(o_data_forward_reg[274]), .B1(n18), .ZN(N1120) );
  INR2D1BWP30P140LVT U1776 ( .A1(o_data_forward_reg[279]), .B1(n18), .ZN(N1125) );
  INR2D1BWP30P140LVT U1777 ( .A1(o_data_forward_reg[282]), .B1(n18), .ZN(N1128) );
  INR2D1BWP30P140LVT U1778 ( .A1(o_data_forward_reg[265]), .B1(n18), .ZN(N1111) );
  INR2D1BWP30P140LVT U1779 ( .A1(o_data_forward_reg[266]), .B1(n18), .ZN(N1112) );
  INR2D1BWP30P140LVT U1780 ( .A1(o_data_forward_reg[283]), .B1(n18), .ZN(N1129) );
  INR2D1BWP30P140LVT U1781 ( .A1(o_data_forward_reg[271]), .B1(n18), .ZN(N1117) );
  INR2D1BWP30P140LVT U1782 ( .A1(o_data_forward_reg[268]), .B1(n18), .ZN(N1114) );
  INR2D1BWP30P140LVT U1783 ( .A1(o_data_forward_reg[278]), .B1(n49), .ZN(N1124) );
  INR2D1BWP30P140LVT U1784 ( .A1(o_data_forward_reg[269]), .B1(n18), .ZN(N1115) );
  INR2D1BWP30P140LVT U1785 ( .A1(o_data_forward_reg[280]), .B1(n49), .ZN(N1126) );
  INR2D1BWP30P140LVT U1786 ( .A1(o_data_forward_reg[275]), .B1(n49), .ZN(N1121) );
  INR2D1BWP30P140LVT U1787 ( .A1(o_data_forward_reg[272]), .B1(n18), .ZN(N1118) );
  INR2D1BWP30P140LVT U1788 ( .A1(o_data_forward_reg[276]), .B1(n18), .ZN(N1122) );
  INR2D1BWP30P140LVT U1789 ( .A1(o_data_forward_reg[277]), .B1(n18), .ZN(N1123) );
  INR2D1BWP30P140LVT U1790 ( .A1(o_data_forward_reg[61]), .B1(n18), .ZN(N2083)
         );
  INR2D1BWP30P140LVT U1791 ( .A1(o_data_forward_reg[59]), .B1(n18), .ZN(N2081)
         );
  INR2D1BWP30P140LVT U1792 ( .A1(o_data_forward_reg[140]), .B1(n18), .ZN(N1658) );
  INR2D1BWP30P140LVT U1793 ( .A1(o_data_forward_reg[137]), .B1(n49), .ZN(N1655) );
  INR2D1BWP30P140LVT U1794 ( .A1(o_data_forward_reg[147]), .B1(n18), .ZN(N1665) );
  INR2D1BWP30P140LVT U1795 ( .A1(o_data_forward_reg[60]), .B1(n18), .ZN(N2082)
         );
  INR2D1BWP30P140LVT U1796 ( .A1(o_data_forward_reg[136]), .B1(n18), .ZN(N1654) );
  INR2D1BWP30P140LVT U1797 ( .A1(o_data_forward_reg[142]), .B1(n49), .ZN(N1660) );
  INR2D1BWP30P140LVT U1798 ( .A1(o_data_forward_reg[143]), .B1(n18), .ZN(N1661) );
  INR2D1BWP30P140LVT U1799 ( .A1(o_data_forward_reg[63]), .B1(n18), .ZN(N2085)
         );
  INR2D1BWP30P140LVT U1800 ( .A1(o_data_forward_reg[138]), .B1(n18), .ZN(N1656) );
  INR2D1BWP30P140LVT U1801 ( .A1(o_data_forward_reg[145]), .B1(n49), .ZN(N1663) );
  INR2D1BWP30P140LVT U1802 ( .A1(o_data_forward_reg[139]), .B1(n18), .ZN(N1657) );
  INR2D1BWP30P140LVT U1803 ( .A1(o_data_forward_reg[135]), .B1(n49), .ZN(N1653) );
  INR2D1BWP30P140LVT U1804 ( .A1(o_data_forward_reg[144]), .B1(n18), .ZN(N1662) );
  INR2D1BWP30P140LVT U1805 ( .A1(o_data_forward_reg[62]), .B1(n18), .ZN(N2084)
         );
  INR2D1BWP30P140LVT U1806 ( .A1(o_data_forward_reg[146]), .B1(n18), .ZN(N1664) );
  INR2D1BWP30P140LVT U1807 ( .A1(o_data_forward_reg[141]), .B1(n49), .ZN(N1659) );
  INR2D1BWP30P140LVT U1808 ( .A1(o_cmd_forward_reg[43]), .B1(n18), .ZN(N866)
         );
  INR2D1BWP30P140LVT U1809 ( .A1(o_cmd_forward_reg[58]), .B1(n49), .ZN(N321)
         );
  INR2D1BWP30P140LVT U1810 ( .A1(o_cmd_forward_reg[54]), .B1(n49), .ZN(N457)
         );
  INR2D1BWP30P140LVT U1811 ( .A1(o_cmd_forward_reg[39]), .B1(n49), .ZN(N1002)
         );
  INR2D1BWP30P140LVT U1812 ( .A1(o_cmd_forward_reg[30]), .B1(n18), .ZN(N1273)
         );
  INR2D1BWP30P140LVT U1813 ( .A1(o_cmd_forward_reg[32]), .B1(n18), .ZN(N1135)
         );
  INR2D1BWP30P140LVT U1814 ( .A1(o_cmd_forward_reg[8]), .B1(n18), .ZN(N1951)
         );
  INR2D1BWP30P140LVT U1815 ( .A1(o_cmd_forward_reg[16]), .B1(n18), .ZN(N1679)
         );
  INR2D1BWP30P140LVT U1816 ( .A1(o_cmd_forward_reg[13]), .B1(n18), .ZN(N1816)
         );
  INR2D1BWP30P140LVT U1817 ( .A1(o_cmd_forward_reg[22]), .B1(n18), .ZN(N1545)
         );
  INR2D1BWP30P140LVT U1818 ( .A1(o_cmd_forward_reg[5]), .B1(n18), .ZN(N2088)
         );
  INR2D1BWP30P140LVT U1819 ( .A1(o_cmd_forward_reg[33]), .B1(n18), .ZN(N1136)
         );
  INR2D1BWP30P140LVT U1820 ( .A1(o_valid_forward_reg[5]), .B1(n18), .ZN(N998)
         );
  INR2D1BWP30P140LVT U1821 ( .A1(o_cmd_forward_reg[48]), .B1(n49), .ZN(N591)
         );
  INR2D1BWP30P140LVT U1822 ( .A1(o_cmd_forward_reg[26]), .B1(n18), .ZN(N1409)
         );
  INR2D1BWP30P140LVT U1823 ( .A1(o_cmd_forward_reg[21]), .B1(n49), .ZN(N1544)
         );
  INR2D1BWP30P140LVT U1824 ( .A1(o_cmd_forward_reg[14]), .B1(n18), .ZN(N1817)
         );
  INR2D1BWP30P140LVT U1825 ( .A1(i_cmd[2]), .B1(n49), .ZN(N185) );
  INR2D1BWP30P140LVT U1826 ( .A1(i_cmd[3]), .B1(n18), .ZN(N186) );
  INR2D1BWP30P140LVT U1827 ( .A1(i_cmd[1]), .B1(n49), .ZN(N184) );
  CKAN2D1BWP30P140LVT U1828 ( .A1(i_data_bus[26]), .A2(n48), .Z(n204) );
  CKAN2D1BWP30P140LVT U1829 ( .A1(i_data_bus[28]), .A2(n48), .Z(n206) );
  CKAN2D1BWP30P140LVT U1830 ( .A1(i_data_bus[29]), .A2(n48), .Z(n207) );
  CKAN2D1BWP30P140LVT U1831 ( .A1(i_data_bus[30]), .A2(n48), .Z(n208) );
  CKAN2D1BWP30P140LVT U1832 ( .A1(n275), .A2(o_data_forward_reg[0]), .Z(n210)
         );
  CKAN2D1BWP30P140LVT U1833 ( .A1(n275), .A2(o_data_forward_reg[1]), .Z(n211)
         );
  CKAN2D1BWP30P140LVT U1834 ( .A1(n275), .A2(o_data_forward_reg[2]), .Z(n212)
         );
  CKAN2D1BWP30P140LVT U1835 ( .A1(n275), .A2(o_data_forward_reg[3]), .Z(n213)
         );
  CKAN2D1BWP30P140LVT U1836 ( .A1(n275), .A2(o_data_forward_reg[4]), .Z(n214)
         );
  CKAN2D1BWP30P140LVT U1837 ( .A1(n275), .A2(o_data_forward_reg[5]), .Z(n215)
         );
  CKAN2D1BWP30P140LVT U1838 ( .A1(n275), .A2(o_data_forward_reg[6]), .Z(n216)
         );
  CKAN2D1BWP30P140LVT U1839 ( .A1(n275), .A2(o_data_forward_reg[7]), .Z(n217)
         );
  CKAN2D1BWP30P140LVT U1840 ( .A1(n275), .A2(o_data_forward_reg[8]), .Z(n218)
         );
  CKAN2D1BWP30P140LVT U1841 ( .A1(n275), .A2(o_data_forward_reg[9]), .Z(n219)
         );
  CKAN2D1BWP30P140LVT U1842 ( .A1(n275), .A2(o_data_forward_reg[10]), .Z(n220)
         );
  CKAN2D1BWP30P140LVT U1843 ( .A1(n275), .A2(o_data_forward_reg[11]), .Z(n221)
         );
  CKAN2D1BWP30P140LVT U1844 ( .A1(n275), .A2(o_data_forward_reg[12]), .Z(n222)
         );
  CKAN2D1BWP30P140LVT U1845 ( .A1(n275), .A2(o_data_forward_reg[13]), .Z(n223)
         );
  CKAN2D1BWP30P140LVT U1846 ( .A1(n275), .A2(o_data_forward_reg[14]), .Z(n224)
         );
  CKAN2D1BWP30P140LVT U1847 ( .A1(n275), .A2(o_data_forward_reg[15]), .Z(n225)
         );
  CKAN2D1BWP30P140LVT U1848 ( .A1(n275), .A2(o_data_forward_reg[16]), .Z(n226)
         );
  CKAN2D1BWP30P140LVT U1849 ( .A1(n275), .A2(o_data_forward_reg[17]), .Z(n227)
         );
  CKAN2D1BWP30P140LVT U1850 ( .A1(n275), .A2(o_data_forward_reg[18]), .Z(n228)
         );
  CKAN2D1BWP30P140LVT U1851 ( .A1(n275), .A2(o_data_forward_reg[19]), .Z(n229)
         );
  CKAN2D1BWP30P140LVT U1852 ( .A1(n275), .A2(o_data_forward_reg[20]), .Z(n230)
         );
  CKAN2D1BWP30P140LVT U1853 ( .A1(n275), .A2(o_data_forward_reg[21]), .Z(n231)
         );
  CKAN2D1BWP30P140LVT U1854 ( .A1(n275), .A2(o_data_forward_reg[22]), .Z(n232)
         );
  CKAN2D1BWP30P140LVT U1855 ( .A1(n275), .A2(o_data_forward_reg[23]), .Z(n233)
         );
  CKAN2D1BWP30P140LVT U1856 ( .A1(n275), .A2(o_data_forward_reg[24]), .Z(n234)
         );
  CKAN2D1BWP30P140LVT U1857 ( .A1(n275), .A2(o_data_forward_reg[25]), .Z(n235)
         );
  CKAN2D1BWP30P140LVT U1858 ( .A1(n274), .A2(i_data_bus[0]), .Z(n236) );
  CKAN2D1BWP30P140LVT U1859 ( .A1(n274), .A2(i_data_bus[1]), .Z(n237) );
  CKAN2D1BWP30P140LVT U1860 ( .A1(n274), .A2(i_data_bus[2]), .Z(n238) );
  CKAN2D1BWP30P140LVT U1861 ( .A1(n274), .A2(i_data_bus[3]), .Z(n239) );
  CKAN2D1BWP30P140LVT U1862 ( .A1(n274), .A2(i_data_bus[4]), .Z(n240) );
  CKAN2D1BWP30P140LVT U1863 ( .A1(n274), .A2(i_data_bus[5]), .Z(n241) );
  CKAN2D1BWP30P140LVT U1864 ( .A1(n274), .A2(i_data_bus[6]), .Z(n242) );
  CKAN2D1BWP30P140LVT U1865 ( .A1(n274), .A2(i_data_bus[7]), .Z(n243) );
  CKAN2D1BWP30P140LVT U1866 ( .A1(n274), .A2(i_data_bus[8]), .Z(n244) );
  CKAN2D1BWP30P140LVT U1867 ( .A1(n274), .A2(i_data_bus[9]), .Z(n245) );
  CKAN2D1BWP30P140LVT U1868 ( .A1(n274), .A2(i_data_bus[10]), .Z(n246) );
  CKAN2D1BWP30P140LVT U1869 ( .A1(n274), .A2(i_data_bus[11]), .Z(n247) );
  CKAN2D1BWP30P140LVT U1870 ( .A1(n274), .A2(i_data_bus[12]), .Z(n248) );
  CKAN2D1BWP30P140LVT U1871 ( .A1(n274), .A2(i_data_bus[13]), .Z(n249) );
  CKAN2D1BWP30P140LVT U1872 ( .A1(n274), .A2(i_data_bus[14]), .Z(n250) );
  CKAN2D1BWP30P140LVT U1873 ( .A1(n274), .A2(i_data_bus[15]), .Z(n251) );
  CKAN2D1BWP30P140LVT U1874 ( .A1(n274), .A2(i_data_bus[16]), .Z(n252) );
  CKAN2D1BWP30P140LVT U1875 ( .A1(n274), .A2(i_data_bus[17]), .Z(n253) );
  CKAN2D1BWP30P140LVT U1876 ( .A1(n274), .A2(i_data_bus[18]), .Z(n254) );
  CKAN2D1BWP30P140LVT U1877 ( .A1(n274), .A2(i_data_bus[19]), .Z(n255) );
  CKAN2D1BWP30P140LVT U1878 ( .A1(n274), .A2(i_data_bus[20]), .Z(n256) );
  CKAN2D1BWP30P140LVT U1879 ( .A1(n274), .A2(i_data_bus[21]), .Z(n257) );
  CKAN2D1BWP30P140LVT U1880 ( .A1(n274), .A2(i_data_bus[22]), .Z(n258) );
  CKAN2D1BWP30P140LVT U1881 ( .A1(n274), .A2(i_data_bus[23]), .Z(n259) );
  CKAN2D1BWP30P140LVT U1882 ( .A1(n274), .A2(i_data_bus[24]), .Z(n260) );
  CKAN2D1BWP30P140LVT U1883 ( .A1(n274), .A2(i_data_bus[25]), .Z(n261) );
  CKAN2D1BWP30P140LVT U1884 ( .A1(n275), .A2(o_data_forward_reg[26]), .Z(n262)
         );
  CKAN2D1BWP30P140LVT U1885 ( .A1(n275), .A2(o_data_forward_reg[27]), .Z(n263)
         );
  CKAN2D1BWP30P140LVT U1886 ( .A1(n275), .A2(o_data_forward_reg[28]), .Z(n264)
         );
  CKAN2D1BWP30P140LVT U1887 ( .A1(n275), .A2(o_data_forward_reg[29]), .Z(n265)
         );
  CKAN2D1BWP30P140LVT U1888 ( .A1(n275), .A2(o_data_forward_reg[30]), .Z(n266)
         );
  CKAN2D1BWP30P140LVT U1889 ( .A1(n275), .A2(o_data_forward_reg[31]), .Z(n267)
         );
  CKAN2D1BWP30P140LVT U1890 ( .A1(n274), .A2(i_data_bus[26]), .Z(n268) );
  CKAN2D1BWP30P140LVT U1891 ( .A1(n274), .A2(i_data_bus[27]), .Z(n269) );
  CKAN2D1BWP30P140LVT U1892 ( .A1(n274), .A2(i_data_bus[28]), .Z(n270) );
  CKAN2D1BWP30P140LVT U1893 ( .A1(n274), .A2(i_data_bus[29]), .Z(n271) );
  CKAN2D1BWP30P140LVT U1894 ( .A1(n274), .A2(i_data_bus[30]), .Z(n272) );
  CKAN2D1BWP30P140LVT U1895 ( .A1(n274), .A2(i_data_bus[31]), .Z(n273) );
  CKAN2D1BWP30P140LVT U1896 ( .A1(n294), .A2(o_data_forward_reg[448]), .Z(N254) );
  CKAN2D1BWP30P140LVT U1897 ( .A1(n294), .A2(o_data_forward_reg[449]), .Z(N255) );
  CKAN2D1BWP30P140LVT U1898 ( .A1(n294), .A2(o_data_forward_reg[450]), .Z(N256) );
  CKAN2D1BWP30P140LVT U1899 ( .A1(n294), .A2(o_data_forward_reg[451]), .Z(N257) );
  CKAN2D1BWP30P140LVT U1900 ( .A1(n294), .A2(o_data_forward_reg[452]), .Z(N258) );
  CKAN2D1BWP30P140LVT U1901 ( .A1(n294), .A2(o_data_forward_reg[453]), .Z(N259) );
  CKAN2D1BWP30P140LVT U1902 ( .A1(n294), .A2(o_data_forward_reg[454]), .Z(N260) );
  CKAN2D1BWP30P140LVT U1903 ( .A1(n294), .A2(o_data_forward_reg[455]), .Z(N261) );
  CKAN2D1BWP30P140LVT U1904 ( .A1(n294), .A2(o_data_forward_reg[456]), .Z(N262) );
  CKAN2D1BWP30P140LVT U1905 ( .A1(n294), .A2(o_data_forward_reg[457]), .Z(N263) );
  CKAN2D1BWP30P140LVT U1906 ( .A1(n294), .A2(o_data_forward_reg[458]), .Z(N264) );
  CKAN2D1BWP30P140LVT U1907 ( .A1(n294), .A2(o_data_forward_reg[459]), .Z(N265) );
  CKAN2D1BWP30P140LVT U1908 ( .A1(n294), .A2(o_data_forward_reg[460]), .Z(N266) );
  CKAN2D1BWP30P140LVT U1909 ( .A1(n294), .A2(o_data_forward_reg[461]), .Z(N267) );
  CKAN2D1BWP30P140LVT U1910 ( .A1(n294), .A2(o_data_forward_reg[462]), .Z(N268) );
  CKAN2D1BWP30P140LVT U1911 ( .A1(n294), .A2(o_data_forward_reg[463]), .Z(N269) );
  CKAN2D1BWP30P140LVT U1912 ( .A1(n294), .A2(o_data_forward_reg[464]), .Z(N270) );
  CKAN2D1BWP30P140LVT U1913 ( .A1(n294), .A2(o_data_forward_reg[465]), .Z(N271) );
  CKAN2D1BWP30P140LVT U1914 ( .A1(n294), .A2(o_data_forward_reg[466]), .Z(N272) );
  CKAN2D1BWP30P140LVT U1915 ( .A1(n294), .A2(o_data_forward_reg[467]), .Z(N273) );
  CKAN2D1BWP30P140LVT U1916 ( .A1(n294), .A2(o_data_forward_reg[468]), .Z(N274) );
  CKAN2D1BWP30P140LVT U1917 ( .A1(n294), .A2(o_data_forward_reg[469]), .Z(N275) );
  CKAN2D1BWP30P140LVT U1918 ( .A1(n294), .A2(o_data_forward_reg[470]), .Z(N276) );
  CKAN2D1BWP30P140LVT U1919 ( .A1(n294), .A2(o_data_forward_reg[471]), .Z(N277) );
  CKAN2D1BWP30P140LVT U1920 ( .A1(n294), .A2(o_data_forward_reg[472]), .Z(N278) );
  CKAN2D1BWP30P140LVT U1921 ( .A1(n294), .A2(o_data_forward_reg[473]), .Z(N279) );
  CKAN2D1BWP30P140LVT U1922 ( .A1(n294), .A2(o_data_forward_reg[474]), .Z(N280) );
  CKAN2D1BWP30P140LVT U1923 ( .A1(n294), .A2(o_data_forward_reg[475]), .Z(N281) );
  CKAN2D1BWP30P140LVT U1924 ( .A1(n294), .A2(o_data_forward_reg[476]), .Z(N282) );
  CKAN2D1BWP30P140LVT U1925 ( .A1(n294), .A2(o_data_forward_reg[477]), .Z(N283) );
  CKAN2D1BWP30P140LVT U1926 ( .A1(n294), .A2(o_data_forward_reg[478]), .Z(N284) );
  CKAN2D1BWP30P140LVT U1927 ( .A1(n294), .A2(o_data_forward_reg[479]), .Z(N285) );
  CKAN2D1BWP30P140LVT U1928 ( .A1(n292), .A2(o_data_forward_reg[416]), .Z(N390) );
  CKAN2D1BWP30P140LVT U1929 ( .A1(n292), .A2(o_data_forward_reg[417]), .Z(N391) );
  CKAN2D1BWP30P140LVT U1930 ( .A1(n292), .A2(o_data_forward_reg[418]), .Z(N392) );
  CKAN2D1BWP30P140LVT U1931 ( .A1(n292), .A2(o_data_forward_reg[419]), .Z(N393) );
  CKAN2D1BWP30P140LVT U1932 ( .A1(n292), .A2(o_data_forward_reg[420]), .Z(N394) );
  CKAN2D1BWP30P140LVT U1933 ( .A1(n292), .A2(o_data_forward_reg[421]), .Z(N395) );
  CKAN2D1BWP30P140LVT U1934 ( .A1(n292), .A2(o_data_forward_reg[422]), .Z(N396) );
  CKAN2D1BWP30P140LVT U1935 ( .A1(n292), .A2(o_data_forward_reg[423]), .Z(N397) );
  CKAN2D1BWP30P140LVT U1936 ( .A1(n292), .A2(o_data_forward_reg[424]), .Z(N398) );
  CKAN2D1BWP30P140LVT U1937 ( .A1(n292), .A2(o_data_forward_reg[425]), .Z(N399) );
  CKAN2D1BWP30P140LVT U1938 ( .A1(n292), .A2(o_data_forward_reg[426]), .Z(N400) );
  CKAN2D1BWP30P140LVT U1939 ( .A1(n292), .A2(o_data_forward_reg[427]), .Z(N401) );
  CKAN2D1BWP30P140LVT U1940 ( .A1(n292), .A2(o_data_forward_reg[428]), .Z(N402) );
  CKAN2D1BWP30P140LVT U1941 ( .A1(n292), .A2(o_data_forward_reg[429]), .Z(N403) );
  CKAN2D1BWP30P140LVT U1942 ( .A1(n292), .A2(o_data_forward_reg[430]), .Z(N404) );
  CKAN2D1BWP30P140LVT U1943 ( .A1(n292), .A2(o_data_forward_reg[431]), .Z(N405) );
  CKAN2D1BWP30P140LVT U1944 ( .A1(n292), .A2(o_data_forward_reg[432]), .Z(N406) );
  CKAN2D1BWP30P140LVT U1945 ( .A1(n292), .A2(o_data_forward_reg[433]), .Z(N407) );
  CKAN2D1BWP30P140LVT U1946 ( .A1(n292), .A2(o_data_forward_reg[434]), .Z(N408) );
  CKAN2D1BWP30P140LVT U1947 ( .A1(n292), .A2(o_data_forward_reg[435]), .Z(N409) );
  CKAN2D1BWP30P140LVT U1948 ( .A1(n292), .A2(o_data_forward_reg[436]), .Z(N410) );
  CKAN2D1BWP30P140LVT U1949 ( .A1(n292), .A2(o_data_forward_reg[437]), .Z(N411) );
  CKAN2D1BWP30P140LVT U1950 ( .A1(n292), .A2(o_data_forward_reg[438]), .Z(N412) );
  CKAN2D1BWP30P140LVT U1951 ( .A1(n292), .A2(o_data_forward_reg[439]), .Z(N413) );
  CKAN2D1BWP30P140LVT U1952 ( .A1(n292), .A2(o_data_forward_reg[440]), .Z(N414) );
  CKAN2D1BWP30P140LVT U1953 ( .A1(n292), .A2(o_data_forward_reg[441]), .Z(N415) );
  CKAN2D1BWP30P140LVT U1954 ( .A1(n292), .A2(o_data_forward_reg[442]), .Z(N416) );
  CKAN2D1BWP30P140LVT U1955 ( .A1(n292), .A2(o_data_forward_reg[443]), .Z(N417) );
  CKAN2D1BWP30P140LVT U1956 ( .A1(n292), .A2(o_data_forward_reg[444]), .Z(N418) );
  CKAN2D1BWP30P140LVT U1957 ( .A1(n292), .A2(o_data_forward_reg[445]), .Z(N419) );
  CKAN2D1BWP30P140LVT U1958 ( .A1(n292), .A2(o_data_forward_reg[446]), .Z(N420) );
  CKAN2D1BWP30P140LVT U1959 ( .A1(n292), .A2(o_data_forward_reg[447]), .Z(N421) );
  CKAN2D1BWP30P140LVT U1960 ( .A1(n291), .A2(o_data_forward_reg[384]), .Z(N526) );
  CKAN2D1BWP30P140LVT U1961 ( .A1(n291), .A2(o_data_forward_reg[385]), .Z(N527) );
  CKAN2D1BWP30P140LVT U1962 ( .A1(n291), .A2(o_data_forward_reg[386]), .Z(N528) );
  CKAN2D1BWP30P140LVT U1963 ( .A1(n291), .A2(o_data_forward_reg[387]), .Z(N529) );
  CKAN2D1BWP30P140LVT U1964 ( .A1(n291), .A2(o_data_forward_reg[388]), .Z(N530) );
  CKAN2D1BWP30P140LVT U1965 ( .A1(n291), .A2(o_data_forward_reg[389]), .Z(N531) );
  CKAN2D1BWP30P140LVT U1966 ( .A1(n291), .A2(o_data_forward_reg[390]), .Z(N532) );
  CKAN2D1BWP30P140LVT U1967 ( .A1(n291), .A2(o_data_forward_reg[391]), .Z(N533) );
  CKAN2D1BWP30P140LVT U1968 ( .A1(n291), .A2(o_data_forward_reg[392]), .Z(N534) );
  CKAN2D1BWP30P140LVT U1969 ( .A1(n291), .A2(o_data_forward_reg[393]), .Z(N535) );
  CKAN2D1BWP30P140LVT U1970 ( .A1(n291), .A2(o_data_forward_reg[394]), .Z(N536) );
  CKAN2D1BWP30P140LVT U1971 ( .A1(n291), .A2(o_data_forward_reg[395]), .Z(N537) );
  CKAN2D1BWP30P140LVT U1972 ( .A1(n291), .A2(o_data_forward_reg[396]), .Z(N538) );
  CKAN2D1BWP30P140LVT U1973 ( .A1(n291), .A2(o_data_forward_reg[397]), .Z(N539) );
  CKAN2D1BWP30P140LVT U1974 ( .A1(n291), .A2(o_data_forward_reg[398]), .Z(N540) );
  CKAN2D1BWP30P140LVT U1975 ( .A1(n291), .A2(o_data_forward_reg[399]), .Z(N541) );
  CKAN2D1BWP30P140LVT U1976 ( .A1(n291), .A2(o_data_forward_reg[400]), .Z(N542) );
  CKAN2D1BWP30P140LVT U1977 ( .A1(n291), .A2(o_data_forward_reg[401]), .Z(N543) );
  CKAN2D1BWP30P140LVT U1978 ( .A1(n291), .A2(o_data_forward_reg[402]), .Z(N544) );
  CKAN2D1BWP30P140LVT U1979 ( .A1(n291), .A2(o_data_forward_reg[403]), .Z(N545) );
  CKAN2D1BWP30P140LVT U1980 ( .A1(n291), .A2(o_data_forward_reg[404]), .Z(N546) );
  CKAN2D1BWP30P140LVT U1981 ( .A1(n291), .A2(o_data_forward_reg[405]), .Z(N547) );
  CKAN2D1BWP30P140LVT U1982 ( .A1(n291), .A2(o_data_forward_reg[406]), .Z(N548) );
  CKAN2D1BWP30P140LVT U1983 ( .A1(n291), .A2(o_data_forward_reg[407]), .Z(N549) );
  CKAN2D1BWP30P140LVT U1984 ( .A1(n291), .A2(o_data_forward_reg[408]), .Z(N550) );
  CKAN2D1BWP30P140LVT U1985 ( .A1(n291), .A2(o_data_forward_reg[409]), .Z(N551) );
  CKAN2D1BWP30P140LVT U1986 ( .A1(n291), .A2(o_data_forward_reg[410]), .Z(N552) );
  CKAN2D1BWP30P140LVT U1987 ( .A1(n291), .A2(o_data_forward_reg[411]), .Z(N553) );
  CKAN2D1BWP30P140LVT U1988 ( .A1(n291), .A2(o_data_forward_reg[412]), .Z(N554) );
  CKAN2D1BWP30P140LVT U1989 ( .A1(n291), .A2(o_data_forward_reg[413]), .Z(N555) );
  CKAN2D1BWP30P140LVT U1990 ( .A1(n291), .A2(o_data_forward_reg[414]), .Z(N556) );
  CKAN2D1BWP30P140LVT U1991 ( .A1(n291), .A2(o_data_forward_reg[415]), .Z(N557) );
  CKAN2D1BWP30P140LVT U1992 ( .A1(n289), .A2(o_data_forward_reg[352]), .Z(N662) );
  CKAN2D1BWP30P140LVT U1993 ( .A1(n289), .A2(o_data_forward_reg[353]), .Z(N663) );
  CKAN2D1BWP30P140LVT U1994 ( .A1(n289), .A2(o_data_forward_reg[354]), .Z(N664) );
  CKAN2D1BWP30P140LVT U1995 ( .A1(n289), .A2(o_data_forward_reg[355]), .Z(N665) );
  CKAN2D1BWP30P140LVT U1996 ( .A1(n289), .A2(o_data_forward_reg[356]), .Z(N666) );
  CKAN2D1BWP30P140LVT U1997 ( .A1(n289), .A2(o_data_forward_reg[357]), .Z(N667) );
  CKAN2D1BWP30P140LVT U1998 ( .A1(n289), .A2(o_data_forward_reg[358]), .Z(N668) );
  CKAN2D1BWP30P140LVT U1999 ( .A1(n289), .A2(o_data_forward_reg[359]), .Z(N669) );
  CKAN2D1BWP30P140LVT U2000 ( .A1(n289), .A2(o_data_forward_reg[360]), .Z(N670) );
  CKAN2D1BWP30P140LVT U2001 ( .A1(n289), .A2(o_data_forward_reg[361]), .Z(N671) );
  CKAN2D1BWP30P140LVT U2002 ( .A1(n289), .A2(o_data_forward_reg[362]), .Z(N672) );
  CKAN2D1BWP30P140LVT U2003 ( .A1(n289), .A2(o_data_forward_reg[363]), .Z(N673) );
  CKAN2D1BWP30P140LVT U2004 ( .A1(n289), .A2(o_data_forward_reg[364]), .Z(N674) );
  CKAN2D1BWP30P140LVT U2005 ( .A1(n289), .A2(o_data_forward_reg[365]), .Z(N675) );
  CKAN2D1BWP30P140LVT U2006 ( .A1(n289), .A2(o_data_forward_reg[366]), .Z(N676) );
  CKAN2D1BWP30P140LVT U2007 ( .A1(n289), .A2(o_data_forward_reg[367]), .Z(N677) );
  CKAN2D1BWP30P140LVT U2008 ( .A1(n289), .A2(o_data_forward_reg[368]), .Z(N678) );
  CKAN2D1BWP30P140LVT U2009 ( .A1(n289), .A2(o_data_forward_reg[369]), .Z(N679) );
  CKAN2D1BWP30P140LVT U2010 ( .A1(n289), .A2(o_data_forward_reg[370]), .Z(N680) );
  CKAN2D1BWP30P140LVT U2011 ( .A1(n289), .A2(o_data_forward_reg[371]), .Z(N681) );
  CKAN2D1BWP30P140LVT U2012 ( .A1(n289), .A2(o_data_forward_reg[372]), .Z(N682) );
  CKAN2D1BWP30P140LVT U2013 ( .A1(n289), .A2(o_data_forward_reg[373]), .Z(N683) );
  CKAN2D1BWP30P140LVT U2014 ( .A1(n289), .A2(o_data_forward_reg[374]), .Z(N684) );
  CKAN2D1BWP30P140LVT U2015 ( .A1(n289), .A2(o_data_forward_reg[375]), .Z(N685) );
  CKAN2D1BWP30P140LVT U2016 ( .A1(n289), .A2(o_data_forward_reg[376]), .Z(N686) );
  CKAN2D1BWP30P140LVT U2017 ( .A1(n289), .A2(o_data_forward_reg[377]), .Z(N687) );
  CKAN2D1BWP30P140LVT U2018 ( .A1(n289), .A2(o_data_forward_reg[378]), .Z(N688) );
  CKAN2D1BWP30P140LVT U2019 ( .A1(n289), .A2(o_data_forward_reg[379]), .Z(N689) );
  CKAN2D1BWP30P140LVT U2020 ( .A1(n289), .A2(o_data_forward_reg[380]), .Z(N690) );
  CKAN2D1BWP30P140LVT U2021 ( .A1(n289), .A2(o_data_forward_reg[381]), .Z(N691) );
  CKAN2D1BWP30P140LVT U2022 ( .A1(n289), .A2(o_data_forward_reg[382]), .Z(N692) );
  CKAN2D1BWP30P140LVT U2023 ( .A1(n289), .A2(o_data_forward_reg[383]), .Z(N693) );
  CKAN2D1BWP30P140LVT U2024 ( .A1(n286), .A2(o_data_forward_reg[288]), .Z(N934) );
  CKAN2D1BWP30P140LVT U2025 ( .A1(n286), .A2(o_data_forward_reg[289]), .Z(N935) );
  CKAN2D1BWP30P140LVT U2026 ( .A1(n286), .A2(o_data_forward_reg[290]), .Z(N936) );
  CKAN2D1BWP30P140LVT U2027 ( .A1(n286), .A2(o_data_forward_reg[291]), .Z(N937) );
  CKAN2D1BWP30P140LVT U2028 ( .A1(n286), .A2(o_data_forward_reg[292]), .Z(N938) );
  CKAN2D1BWP30P140LVT U2029 ( .A1(n286), .A2(o_data_forward_reg[293]), .Z(N939) );
  CKAN2D1BWP30P140LVT U2030 ( .A1(n286), .A2(o_data_forward_reg[294]), .Z(N940) );
  CKAN2D1BWP30P140LVT U2031 ( .A1(n286), .A2(o_data_forward_reg[295]), .Z(N941) );
  CKAN2D1BWP30P140LVT U2032 ( .A1(n286), .A2(o_data_forward_reg[296]), .Z(N942) );
  CKAN2D1BWP30P140LVT U2033 ( .A1(n286), .A2(o_data_forward_reg[297]), .Z(N943) );
  CKAN2D1BWP30P140LVT U2034 ( .A1(n286), .A2(o_data_forward_reg[298]), .Z(N944) );
  CKAN2D1BWP30P140LVT U2035 ( .A1(n286), .A2(o_data_forward_reg[299]), .Z(N945) );
  CKAN2D1BWP30P140LVT U2036 ( .A1(n286), .A2(o_data_forward_reg[300]), .Z(N946) );
  CKAN2D1BWP30P140LVT U2037 ( .A1(n286), .A2(o_data_forward_reg[301]), .Z(N947) );
  CKAN2D1BWP30P140LVT U2038 ( .A1(n286), .A2(o_data_forward_reg[302]), .Z(N948) );
  CKAN2D1BWP30P140LVT U2039 ( .A1(n286), .A2(o_data_forward_reg[303]), .Z(N949) );
  CKAN2D1BWP30P140LVT U2040 ( .A1(n286), .A2(o_data_forward_reg[304]), .Z(N950) );
  CKAN2D1BWP30P140LVT U2041 ( .A1(n286), .A2(o_data_forward_reg[305]), .Z(N951) );
  CKAN2D1BWP30P140LVT U2042 ( .A1(n286), .A2(o_data_forward_reg[306]), .Z(N952) );
  CKAN2D1BWP30P140LVT U2043 ( .A1(n286), .A2(o_data_forward_reg[307]), .Z(N953) );
  CKAN2D1BWP30P140LVT U2044 ( .A1(n286), .A2(o_data_forward_reg[308]), .Z(N954) );
  CKAN2D1BWP30P140LVT U2045 ( .A1(n286), .A2(o_data_forward_reg[309]), .Z(N955) );
  CKAN2D1BWP30P140LVT U2046 ( .A1(n286), .A2(o_data_forward_reg[310]), .Z(N956) );
  CKAN2D1BWP30P140LVT U2047 ( .A1(n286), .A2(o_data_forward_reg[311]), .Z(N957) );
  CKAN2D1BWP30P140LVT U2048 ( .A1(n286), .A2(o_data_forward_reg[312]), .Z(N958) );
  CKAN2D1BWP30P140LVT U2049 ( .A1(n286), .A2(o_data_forward_reg[313]), .Z(N959) );
  CKAN2D1BWP30P140LVT U2050 ( .A1(n286), .A2(o_data_forward_reg[314]), .Z(N960) );
  CKAN2D1BWP30P140LVT U2051 ( .A1(n286), .A2(o_data_forward_reg[315]), .Z(N961) );
  CKAN2D1BWP30P140LVT U2052 ( .A1(n286), .A2(o_data_forward_reg[316]), .Z(N962) );
  CKAN2D1BWP30P140LVT U2053 ( .A1(n286), .A2(o_data_forward_reg[317]), .Z(N963) );
  CKAN2D1BWP30P140LVT U2054 ( .A1(n286), .A2(o_data_forward_reg[318]), .Z(N964) );
  CKAN2D1BWP30P140LVT U2055 ( .A1(n286), .A2(o_data_forward_reg[319]), .Z(N965) );
  CKAN2D1BWP30P140LVT U2056 ( .A1(n19), .A2(o_data_forward_reg[256]), .Z(N1070) );
  CKAN2D1BWP30P140LVT U2057 ( .A1(n19), .A2(o_data_forward_reg[257]), .Z(N1071) );
  CKAN2D1BWP30P140LVT U2058 ( .A1(n19), .A2(o_data_forward_reg[258]), .Z(N1072) );
  CKAN2D1BWP30P140LVT U2059 ( .A1(n19), .A2(o_data_forward_reg[259]), .Z(N1073) );
  CKAN2D1BWP30P140LVT U2060 ( .A1(n19), .A2(o_data_forward_reg[260]), .Z(N1074) );
  CKAN2D1BWP30P140LVT U2061 ( .A1(n19), .A2(o_data_forward_reg[261]), .Z(N1075) );
  CKAN2D1BWP30P140LVT U2062 ( .A1(n19), .A2(o_data_forward_reg[262]), .Z(N1076) );
  CKAN2D1BWP30P140LVT U2063 ( .A1(n19), .A2(o_data_forward_reg[263]), .Z(N1077) );
  CKAN2D1BWP30P140LVT U2064 ( .A1(n19), .A2(o_data_forward_reg[264]), .Z(N1078) );
  CKAN2D1BWP30P140LVT U2065 ( .A1(n19), .A2(o_data_forward_reg[265]), .Z(N1079) );
  CKAN2D1BWP30P140LVT U2066 ( .A1(n19), .A2(o_data_forward_reg[266]), .Z(N1080) );
  CKAN2D1BWP30P140LVT U2067 ( .A1(n19), .A2(o_data_forward_reg[267]), .Z(N1081) );
  CKAN2D1BWP30P140LVT U2068 ( .A1(n19), .A2(o_data_forward_reg[268]), .Z(N1082) );
  CKAN2D1BWP30P140LVT U2069 ( .A1(n19), .A2(o_data_forward_reg[269]), .Z(N1083) );
  CKAN2D1BWP30P140LVT U2070 ( .A1(n19), .A2(o_data_forward_reg[270]), .Z(N1084) );
  CKAN2D1BWP30P140LVT U2071 ( .A1(n19), .A2(o_data_forward_reg[271]), .Z(N1085) );
  CKAN2D1BWP30P140LVT U2072 ( .A1(n19), .A2(o_data_forward_reg[272]), .Z(N1086) );
  CKAN2D1BWP30P140LVT U2073 ( .A1(n19), .A2(o_data_forward_reg[273]), .Z(N1087) );
  CKAN2D1BWP30P140LVT U2074 ( .A1(n19), .A2(o_data_forward_reg[274]), .Z(N1088) );
  CKAN2D1BWP30P140LVT U2075 ( .A1(n19), .A2(o_data_forward_reg[275]), .Z(N1089) );
  CKAN2D1BWP30P140LVT U2076 ( .A1(n19), .A2(o_data_forward_reg[276]), .Z(N1090) );
  CKAN2D1BWP30P140LVT U2077 ( .A1(n19), .A2(o_data_forward_reg[277]), .Z(N1091) );
  CKAN2D1BWP30P140LVT U2078 ( .A1(n19), .A2(o_data_forward_reg[278]), .Z(N1092) );
  CKAN2D1BWP30P140LVT U2079 ( .A1(n19), .A2(o_data_forward_reg[279]), .Z(N1093) );
  CKAN2D1BWP30P140LVT U2080 ( .A1(n19), .A2(o_data_forward_reg[280]), .Z(N1094) );
  CKAN2D1BWP30P140LVT U2081 ( .A1(n19), .A2(o_data_forward_reg[281]), .Z(N1095) );
  CKAN2D1BWP30P140LVT U2082 ( .A1(n19), .A2(o_data_forward_reg[282]), .Z(N1096) );
  CKAN2D1BWP30P140LVT U2083 ( .A1(n19), .A2(o_data_forward_reg[283]), .Z(N1097) );
  CKAN2D1BWP30P140LVT U2084 ( .A1(n19), .A2(o_data_forward_reg[284]), .Z(N1098) );
  CKAN2D1BWP30P140LVT U2085 ( .A1(n19), .A2(o_data_forward_reg[285]), .Z(N1099) );
  CKAN2D1BWP30P140LVT U2086 ( .A1(n19), .A2(o_data_forward_reg[286]), .Z(N1100) );
  CKAN2D1BWP30P140LVT U2087 ( .A1(n19), .A2(o_data_forward_reg[287]), .Z(N1101) );
  CKAN2D1BWP30P140LVT U2088 ( .A1(n283), .A2(o_data_forward_reg[224]), .Z(
        N1206) );
  CKAN2D1BWP30P140LVT U2089 ( .A1(n283), .A2(o_data_forward_reg[225]), .Z(
        N1207) );
  CKAN2D1BWP30P140LVT U2090 ( .A1(n283), .A2(o_data_forward_reg[226]), .Z(
        N1208) );
  CKAN2D1BWP30P140LVT U2091 ( .A1(n283), .A2(o_data_forward_reg[227]), .Z(
        N1209) );
  CKAN2D1BWP30P140LVT U2092 ( .A1(n283), .A2(o_data_forward_reg[228]), .Z(
        N1210) );
  CKAN2D1BWP30P140LVT U2093 ( .A1(n283), .A2(o_data_forward_reg[229]), .Z(
        N1211) );
  CKAN2D1BWP30P140LVT U2094 ( .A1(n283), .A2(o_data_forward_reg[230]), .Z(
        N1212) );
  CKAN2D1BWP30P140LVT U2095 ( .A1(n283), .A2(o_data_forward_reg[231]), .Z(
        N1213) );
  CKAN2D1BWP30P140LVT U2096 ( .A1(n283), .A2(o_data_forward_reg[232]), .Z(
        N1214) );
  CKAN2D1BWP30P140LVT U2097 ( .A1(n283), .A2(o_data_forward_reg[233]), .Z(
        N1215) );
  CKAN2D1BWP30P140LVT U2098 ( .A1(n283), .A2(o_data_forward_reg[234]), .Z(
        N1216) );
  CKAN2D1BWP30P140LVT U2099 ( .A1(n283), .A2(o_data_forward_reg[235]), .Z(
        N1217) );
  CKAN2D1BWP30P140LVT U2100 ( .A1(n283), .A2(o_data_forward_reg[236]), .Z(
        N1218) );
  CKAN2D1BWP30P140LVT U2101 ( .A1(n283), .A2(o_data_forward_reg[237]), .Z(
        N1219) );
  CKAN2D1BWP30P140LVT U2102 ( .A1(n283), .A2(o_data_forward_reg[238]), .Z(
        N1220) );
  CKAN2D1BWP30P140LVT U2103 ( .A1(n283), .A2(o_data_forward_reg[239]), .Z(
        N1221) );
  CKAN2D1BWP30P140LVT U2104 ( .A1(n283), .A2(o_data_forward_reg[240]), .Z(
        N1222) );
  CKAN2D1BWP30P140LVT U2105 ( .A1(n283), .A2(o_data_forward_reg[241]), .Z(
        N1223) );
  CKAN2D1BWP30P140LVT U2106 ( .A1(n283), .A2(o_data_forward_reg[242]), .Z(
        N1224) );
  CKAN2D1BWP30P140LVT U2107 ( .A1(n283), .A2(o_data_forward_reg[243]), .Z(
        N1225) );
  CKAN2D1BWP30P140LVT U2108 ( .A1(n283), .A2(o_data_forward_reg[244]), .Z(
        N1226) );
  CKAN2D1BWP30P140LVT U2109 ( .A1(n283), .A2(o_data_forward_reg[245]), .Z(
        N1227) );
  CKAN2D1BWP30P140LVT U2110 ( .A1(n283), .A2(o_data_forward_reg[246]), .Z(
        N1228) );
  CKAN2D1BWP30P140LVT U2111 ( .A1(n283), .A2(o_data_forward_reg[247]), .Z(
        N1229) );
  CKAN2D1BWP30P140LVT U2112 ( .A1(n283), .A2(o_data_forward_reg[248]), .Z(
        N1230) );
  CKAN2D1BWP30P140LVT U2113 ( .A1(n283), .A2(o_data_forward_reg[249]), .Z(
        N1231) );
  CKAN2D1BWP30P140LVT U2114 ( .A1(n283), .A2(o_data_forward_reg[250]), .Z(
        N1232) );
  CKAN2D1BWP30P140LVT U2115 ( .A1(n283), .A2(o_data_forward_reg[251]), .Z(
        N1233) );
  CKAN2D1BWP30P140LVT U2116 ( .A1(n283), .A2(o_data_forward_reg[252]), .Z(
        N1234) );
  CKAN2D1BWP30P140LVT U2117 ( .A1(n283), .A2(o_data_forward_reg[253]), .Z(
        N1235) );
  CKAN2D1BWP30P140LVT U2118 ( .A1(n283), .A2(o_data_forward_reg[254]), .Z(
        N1236) );
  CKAN2D1BWP30P140LVT U2119 ( .A1(n283), .A2(o_data_forward_reg[255]), .Z(
        N1237) );
  CKAN2D1BWP30P140LVT U2120 ( .A1(n21), .A2(o_data_forward_reg[160]), .Z(N1478) );
  CKAN2D1BWP30P140LVT U2121 ( .A1(n21), .A2(o_data_forward_reg[161]), .Z(N1479) );
  CKAN2D1BWP30P140LVT U2122 ( .A1(n21), .A2(o_data_forward_reg[162]), .Z(N1480) );
  CKAN2D1BWP30P140LVT U2123 ( .A1(n21), .A2(o_data_forward_reg[163]), .Z(N1481) );
  CKAN2D1BWP30P140LVT U2124 ( .A1(n21), .A2(o_data_forward_reg[164]), .Z(N1482) );
  CKAN2D1BWP30P140LVT U2125 ( .A1(n21), .A2(o_data_forward_reg[165]), .Z(N1483) );
  CKAN2D1BWP30P140LVT U2126 ( .A1(n21), .A2(o_data_forward_reg[166]), .Z(N1484) );
  CKAN2D1BWP30P140LVT U2127 ( .A1(n21), .A2(o_data_forward_reg[167]), .Z(N1485) );
  CKAN2D1BWP30P140LVT U2128 ( .A1(n21), .A2(o_data_forward_reg[168]), .Z(N1486) );
  CKAN2D1BWP30P140LVT U2129 ( .A1(n21), .A2(o_data_forward_reg[169]), .Z(N1487) );
  CKAN2D1BWP30P140LVT U2130 ( .A1(n21), .A2(o_data_forward_reg[170]), .Z(N1488) );
  CKAN2D1BWP30P140LVT U2131 ( .A1(n21), .A2(o_data_forward_reg[171]), .Z(N1489) );
  CKAN2D1BWP30P140LVT U2132 ( .A1(n21), .A2(o_data_forward_reg[172]), .Z(N1490) );
  CKAN2D1BWP30P140LVT U2133 ( .A1(n21), .A2(o_data_forward_reg[173]), .Z(N1491) );
  CKAN2D1BWP30P140LVT U2134 ( .A1(n21), .A2(o_data_forward_reg[174]), .Z(N1492) );
  CKAN2D1BWP30P140LVT U2135 ( .A1(n21), .A2(o_data_forward_reg[175]), .Z(N1493) );
  CKAN2D1BWP30P140LVT U2136 ( .A1(n21), .A2(o_data_forward_reg[176]), .Z(N1494) );
  CKAN2D1BWP30P140LVT U2137 ( .A1(n21), .A2(o_data_forward_reg[177]), .Z(N1495) );
  CKAN2D1BWP30P140LVT U2138 ( .A1(n21), .A2(o_data_forward_reg[178]), .Z(N1496) );
  CKAN2D1BWP30P140LVT U2139 ( .A1(n21), .A2(o_data_forward_reg[179]), .Z(N1497) );
  CKAN2D1BWP30P140LVT U2140 ( .A1(n21), .A2(o_data_forward_reg[180]), .Z(N1498) );
  CKAN2D1BWP30P140LVT U2141 ( .A1(n21), .A2(o_data_forward_reg[181]), .Z(N1499) );
  CKAN2D1BWP30P140LVT U2142 ( .A1(n21), .A2(o_data_forward_reg[182]), .Z(N1500) );
  CKAN2D1BWP30P140LVT U2143 ( .A1(n21), .A2(o_data_forward_reg[183]), .Z(N1501) );
  CKAN2D1BWP30P140LVT U2144 ( .A1(n21), .A2(o_data_forward_reg[184]), .Z(N1502) );
  CKAN2D1BWP30P140LVT U2145 ( .A1(n21), .A2(o_data_forward_reg[185]), .Z(N1503) );
  CKAN2D1BWP30P140LVT U2146 ( .A1(n21), .A2(o_data_forward_reg[186]), .Z(N1504) );
  CKAN2D1BWP30P140LVT U2147 ( .A1(n21), .A2(o_data_forward_reg[187]), .Z(N1505) );
  CKAN2D1BWP30P140LVT U2148 ( .A1(n21), .A2(o_data_forward_reg[188]), .Z(N1506) );
  CKAN2D1BWP30P140LVT U2149 ( .A1(n21), .A2(o_data_forward_reg[189]), .Z(N1507) );
  CKAN2D1BWP30P140LVT U2150 ( .A1(n21), .A2(o_data_forward_reg[190]), .Z(N1508) );
  CKAN2D1BWP30P140LVT U2151 ( .A1(n21), .A2(o_data_forward_reg[191]), .Z(N1509) );
  CKAN2D1BWP30P140LVT U2152 ( .A1(n20), .A2(o_data_forward_reg[96]), .Z(N1750)
         );
  CKAN2D1BWP30P140LVT U2153 ( .A1(n20), .A2(o_data_forward_reg[97]), .Z(N1751)
         );
  CKAN2D1BWP30P140LVT U2154 ( .A1(n20), .A2(o_data_forward_reg[98]), .Z(N1752)
         );
  CKAN2D1BWP30P140LVT U2155 ( .A1(n20), .A2(o_data_forward_reg[99]), .Z(N1753)
         );
  CKAN2D1BWP30P140LVT U2156 ( .A1(n20), .A2(o_data_forward_reg[100]), .Z(N1754) );
  CKAN2D1BWP30P140LVT U2157 ( .A1(n20), .A2(o_data_forward_reg[101]), .Z(N1755) );
  CKAN2D1BWP30P140LVT U2158 ( .A1(n20), .A2(o_data_forward_reg[102]), .Z(N1756) );
  CKAN2D1BWP30P140LVT U2159 ( .A1(n20), .A2(o_data_forward_reg[103]), .Z(N1757) );
  CKAN2D1BWP30P140LVT U2160 ( .A1(n20), .A2(o_data_forward_reg[104]), .Z(N1758) );
  CKAN2D1BWP30P140LVT U2161 ( .A1(n20), .A2(o_data_forward_reg[105]), .Z(N1759) );
  CKAN2D1BWP30P140LVT U2162 ( .A1(n20), .A2(o_data_forward_reg[106]), .Z(N1760) );
  CKAN2D1BWP30P140LVT U2163 ( .A1(n20), .A2(o_data_forward_reg[107]), .Z(N1761) );
  CKAN2D1BWP30P140LVT U2164 ( .A1(n20), .A2(o_data_forward_reg[108]), .Z(N1762) );
  CKAN2D1BWP30P140LVT U2165 ( .A1(n20), .A2(o_data_forward_reg[109]), .Z(N1763) );
  CKAN2D1BWP30P140LVT U2166 ( .A1(n20), .A2(o_data_forward_reg[110]), .Z(N1764) );
  CKAN2D1BWP30P140LVT U2167 ( .A1(n20), .A2(o_data_forward_reg[111]), .Z(N1765) );
  CKAN2D1BWP30P140LVT U2168 ( .A1(n20), .A2(o_data_forward_reg[112]), .Z(N1766) );
  CKAN2D1BWP30P140LVT U2169 ( .A1(n20), .A2(o_data_forward_reg[113]), .Z(N1767) );
  CKAN2D1BWP30P140LVT U2170 ( .A1(n20), .A2(o_data_forward_reg[114]), .Z(N1768) );
  CKAN2D1BWP30P140LVT U2171 ( .A1(n20), .A2(o_data_forward_reg[115]), .Z(N1769) );
  CKAN2D1BWP30P140LVT U2172 ( .A1(n20), .A2(o_data_forward_reg[116]), .Z(N1770) );
  CKAN2D1BWP30P140LVT U2173 ( .A1(n20), .A2(o_data_forward_reg[117]), .Z(N1771) );
  CKAN2D1BWP30P140LVT U2174 ( .A1(n20), .A2(o_data_forward_reg[118]), .Z(N1772) );
  CKAN2D1BWP30P140LVT U2175 ( .A1(n20), .A2(o_data_forward_reg[119]), .Z(N1773) );
  CKAN2D1BWP30P140LVT U2176 ( .A1(n20), .A2(o_data_forward_reg[120]), .Z(N1774) );
  CKAN2D1BWP30P140LVT U2177 ( .A1(n20), .A2(o_data_forward_reg[121]), .Z(N1775) );
  CKAN2D1BWP30P140LVT U2178 ( .A1(n20), .A2(o_data_forward_reg[122]), .Z(N1776) );
  CKAN2D1BWP30P140LVT U2179 ( .A1(n20), .A2(o_data_forward_reg[123]), .Z(N1777) );
  CKAN2D1BWP30P140LVT U2180 ( .A1(n20), .A2(o_data_forward_reg[124]), .Z(N1778) );
  CKAN2D1BWP30P140LVT U2181 ( .A1(n20), .A2(o_data_forward_reg[125]), .Z(N1779) );
  CKAN2D1BWP30P140LVT U2182 ( .A1(n20), .A2(o_data_forward_reg[126]), .Z(N1780) );
  CKAN2D1BWP30P140LVT U2183 ( .A1(n20), .A2(o_data_forward_reg[127]), .Z(N1781) );
  INR2D1BWP30P140LVT U2184 ( .A1(o_cmd_forward_reg[4]), .B1(n18), .ZN(N2087)
         );
  INR2D1BWP30P140LVT U2185 ( .A1(o_cmd_forward_reg[7]), .B1(n18), .ZN(N2090)
         );
  INR2D1BWP30P140LVT U2186 ( .A1(o_valid_forward_reg[13]), .B1(n18), .ZN(N2086) );
  INR2D1BWP30P140LVT U2187 ( .A1(o_cmd_forward_reg[9]), .B1(n49), .ZN(N1952)
         );
  INR2D1BWP30P140LVT U2188 ( .A1(o_cmd_forward_reg[10]), .B1(n18), .ZN(N1953)
         );
  INR2D1BWP30P140LVT U2189 ( .A1(o_valid_forward_reg[12]), .B1(n18), .ZN(N1950) );
  INR2D1BWP30P140LVT U2190 ( .A1(o_cmd_forward_reg[12]), .B1(n49), .ZN(N1815)
         );
  INR2D1BWP30P140LVT U2191 ( .A1(o_valid_forward_reg[11]), .B1(n18), .ZN(N1814) );
  INR2D1BWP30P140LVT U2192 ( .A1(o_cmd_forward_reg[18]), .B1(n18), .ZN(N1681)
         );
  INR2D1BWP30P140LVT U2193 ( .A1(o_cmd_forward_reg[19]), .B1(n18), .ZN(N1682)
         );
  INR2D1BWP30P140LVT U2194 ( .A1(o_valid_forward_reg[10]), .B1(n18), .ZN(N1678) );
  INR2D1BWP30P140LVT U2195 ( .A1(o_cmd_forward_reg[20]), .B1(n49), .ZN(N1543)
         );
  INR2D1BWP30P140LVT U2196 ( .A1(o_valid_forward_reg[9]), .B1(n18), .ZN(N1542)
         );
  INR2D1BWP30P140LVT U2197 ( .A1(o_cmd_forward_reg[25]), .B1(n49), .ZN(N1408)
         );
  INR2D1BWP30P140LVT U2198 ( .A1(o_cmd_forward_reg[27]), .B1(n18), .ZN(N1410)
         );
  INR2D1BWP30P140LVT U2199 ( .A1(o_valid_forward_reg[8]), .B1(n18), .ZN(N1406)
         );
  INR2D1BWP30P140LVT U2200 ( .A1(o_cmd_forward_reg[28]), .B1(n49), .ZN(N1271)
         );
  INR2D1BWP30P140LVT U2201 ( .A1(o_valid_forward_reg[7]), .B1(n49), .ZN(N1270)
         );
  INR2D1BWP30P140LVT U2202 ( .A1(o_cmd_forward_reg[35]), .B1(n18), .ZN(N1138)
         );
  INR2D1BWP30P140LVT U2203 ( .A1(o_valid_forward_reg[6]), .B1(n18), .ZN(N1134)
         );
  INR2D1BWP30P140LVT U2204 ( .A1(o_cmd_forward_reg[36]), .B1(n18), .ZN(N999)
         );
  INR2D1BWP30P140LVT U2205 ( .A1(o_cmd_forward_reg[38]), .B1(n49), .ZN(N1001)
         );
  INR2D1BWP30P140LVT U2206 ( .A1(o_cmd_forward_reg[41]), .B1(n18), .ZN(N864)
         );
  INR2D1BWP30P140LVT U2207 ( .A1(o_cmd_forward_reg[42]), .B1(n49), .ZN(N865)
         );
  INR2D1BWP30P140LVT U2208 ( .A1(o_valid_forward_reg[4]), .B1(n18), .ZN(N862)
         );
  INR2D1BWP30P140LVT U2209 ( .A1(o_cmd_forward_reg[44]), .B1(n18), .ZN(N727)
         );
  INR2D1BWP30P140LVT U2210 ( .A1(o_valid_forward_reg[3]), .B1(n18), .ZN(N726)
         );
  INR2D1BWP30P140LVT U2211 ( .A1(o_cmd_forward_reg[50]), .B1(n49), .ZN(N593)
         );
  INR2D1BWP30P140LVT U2212 ( .A1(o_valid_forward_reg[2]), .B1(n18), .ZN(N590)
         );
  INR2D1BWP30P140LVT U2213 ( .A1(o_cmd_forward_reg[52]), .B1(n18), .ZN(N455)
         );
  INR2D1BWP30P140LVT U2214 ( .A1(o_valid_forward_reg[1]), .B1(n18), .ZN(N454)
         );
  INR2D1BWP30P140LVT U2215 ( .A1(o_cmd_forward_reg[57]), .B1(n18), .ZN(N320)
         );
  INR2D1BWP30P140LVT U2216 ( .A1(o_valid_forward_reg[0]), .B1(n18), .ZN(N318)
         );
  INR2D1BWP30P140LVT U2217 ( .A1(i_cmd[0]), .B1(n18), .ZN(N183) );
endmodule

