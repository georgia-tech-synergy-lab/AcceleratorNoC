
module mux_2x1_simple_seq ( clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, 
        i_en );
  input [1:0] i_valid;
  input [63:0] i_data_bus;
  output [31:0] o_data_bus;
  input clk, rst, i_en;
  output o_valid;
  wire   N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44;
  wire   [63:0] buf_def_0__i_data_o_buf;
  wire   [63:0] buf_def_1__i_data_o_buf;
  wire   [63:0] buf_def_2__i_data_o_buf;
  wire   [63:0] buf_def_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_assign_0__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[0]), .Z(buf_def_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_assign_0__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[0]), .Z(buf_def_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_assign_0__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[0]), .Z(buf_def_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_assign_0__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[0]), .Z(buf_def_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_assign_1__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[1]), .Z(buf_def_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_assign_1__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[1]), .Z(buf_def_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_assign_1__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[1]), .Z(buf_def_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_assign_1__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[1]), .Z(buf_def_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_assign_2__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[2]), .Z(buf_def_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_assign_2__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[2]), .Z(buf_def_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_assign_2__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[2]), .Z(buf_def_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_assign_2__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[2]), .Z(buf_def_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_assign_3__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[3]), .Z(buf_def_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_assign_3__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[3]), .Z(buf_def_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_assign_3__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[3]), .Z(buf_def_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_assign_3__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[3]), .Z(buf_def_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_assign_4__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[4]), .Z(buf_def_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_assign_4__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[4]), .Z(buf_def_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_assign_4__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[4]), .Z(buf_def_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_assign_4__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[4]), .Z(buf_def_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_assign_5__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[5]), .Z(buf_def_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_assign_5__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[5]), .Z(buf_def_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_assign_5__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[5]), .Z(buf_def_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_assign_5__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[5]), .Z(buf_def_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_assign_6__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[6]), .Z(buf_def_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_assign_6__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[6]), .Z(buf_def_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_assign_6__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[6]), .Z(buf_def_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_assign_6__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[6]), .Z(buf_def_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_assign_7__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[7]), .Z(buf_def_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_assign_7__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[7]), .Z(buf_def_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_assign_7__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[7]), .Z(buf_def_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_assign_7__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[7]), .Z(buf_def_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_assign_8__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[8]), .Z(buf_def_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_assign_8__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[8]), .Z(buf_def_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_assign_8__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[8]), .Z(buf_def_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_assign_8__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[8]), .Z(buf_def_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_assign_9__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[9]), .Z(buf_def_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_assign_9__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[9]), .Z(buf_def_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_assign_9__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[9]), .Z(buf_def_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_assign_9__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[9]), .Z(buf_def_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_assign_10__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[10]), .Z(buf_def_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_assign_10__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[10]), .Z(buf_def_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_assign_10__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[10]), .Z(buf_def_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_assign_10__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[10]), .Z(buf_def_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_assign_11__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[11]), .Z(buf_def_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_assign_11__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[11]), .Z(buf_def_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_assign_11__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[11]), .Z(buf_def_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_assign_11__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[11]), .Z(buf_def_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_assign_12__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[12]), .Z(buf_def_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_assign_12__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[12]), .Z(buf_def_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_assign_12__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[12]), .Z(buf_def_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_assign_12__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[12]), .Z(buf_def_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_assign_13__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[13]), .Z(buf_def_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_assign_13__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[13]), .Z(buf_def_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_assign_13__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[13]), .Z(buf_def_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_assign_13__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[13]), .Z(buf_def_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_assign_14__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[14]), .Z(buf_def_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_assign_14__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[14]), .Z(buf_def_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_assign_14__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[14]), .Z(buf_def_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_assign_14__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[14]), .Z(buf_def_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_assign_15__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[15]), .Z(buf_def_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_assign_15__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[15]), .Z(buf_def_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_assign_15__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[15]), .Z(buf_def_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_assign_15__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[15]), .Z(buf_def_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_assign_16__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[16]), .Z(buf_def_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_assign_16__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[16]), .Z(buf_def_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_assign_16__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[16]), .Z(buf_def_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_assign_16__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[16]), .Z(buf_def_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_assign_17__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[17]), .Z(buf_def_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_assign_17__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[17]), .Z(buf_def_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_assign_17__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[17]), .Z(buf_def_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_assign_17__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[17]), .Z(buf_def_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_assign_18__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[18]), .Z(buf_def_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_assign_18__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[18]), .Z(buf_def_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_assign_18__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[18]), .Z(buf_def_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_assign_18__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[18]), .Z(buf_def_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_assign_19__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[19]), .Z(buf_def_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_assign_19__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[19]), .Z(buf_def_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_assign_19__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[19]), .Z(buf_def_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_assign_19__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[19]), .Z(buf_def_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_assign_20__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[20]), .Z(buf_def_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_assign_20__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[20]), .Z(buf_def_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_assign_20__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[20]), .Z(buf_def_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_assign_20__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[20]), .Z(buf_def_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_assign_21__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[21]), .Z(buf_def_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_assign_21__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[21]), .Z(buf_def_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_assign_21__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[21]), .Z(buf_def_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_assign_21__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[21]), .Z(buf_def_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_assign_22__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[22]), .Z(buf_def_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_assign_22__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[22]), .Z(buf_def_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_assign_22__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[22]), .Z(buf_def_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_assign_22__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[22]), .Z(buf_def_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_assign_23__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[23]), .Z(buf_def_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_assign_23__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[23]), .Z(buf_def_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_assign_23__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[23]), .Z(buf_def_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_assign_23__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[23]), .Z(buf_def_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_assign_24__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[24]), .Z(buf_def_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_assign_24__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[24]), .Z(buf_def_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_assign_24__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[24]), .Z(buf_def_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_assign_24__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[24]), .Z(buf_def_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_assign_25__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[25]), .Z(buf_def_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_assign_25__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[25]), .Z(buf_def_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_assign_25__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[25]), .Z(buf_def_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_assign_25__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[25]), .Z(buf_def_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_assign_26__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[26]), .Z(buf_def_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_assign_26__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[26]), .Z(buf_def_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_assign_26__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[26]), .Z(buf_def_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_assign_26__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[26]), .Z(buf_def_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_assign_27__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[27]), .Z(buf_def_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_assign_27__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[27]), .Z(buf_def_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_assign_27__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[27]), .Z(buf_def_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_assign_27__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[27]), .Z(buf_def_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_assign_28__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[28]), .Z(buf_def_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_assign_28__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[28]), .Z(buf_def_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_assign_28__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[28]), .Z(buf_def_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_assign_28__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[28]), .Z(buf_def_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_assign_29__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[29]), .Z(buf_def_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_assign_29__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[29]), .Z(buf_def_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_assign_29__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[29]), .Z(buf_def_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_assign_29__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[29]), .Z(buf_def_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_assign_30__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[30]), .Z(buf_def_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_assign_30__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[30]), .Z(buf_def_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_assign_30__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[30]), .Z(buf_def_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_assign_30__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[30]), .Z(buf_def_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_assign_31__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[31]), .Z(buf_def_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_assign_31__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[31]), .Z(buf_def_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_assign_31__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[31]), .Z(buf_def_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_assign_31__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[31]), .Z(buf_def_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_assign_32__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[32]), .Z(buf_def_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_assign_32__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[32]), .Z(buf_def_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_assign_32__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[32]), .Z(buf_def_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_assign_32__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[32]), .Z(buf_def_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_assign_33__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[33]), .Z(buf_def_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_assign_33__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[33]), .Z(buf_def_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_assign_33__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[33]), .Z(buf_def_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_assign_33__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[33]), .Z(buf_def_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_assign_34__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[34]), .Z(buf_def_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_assign_34__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[34]), .Z(buf_def_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_assign_34__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[34]), .Z(buf_def_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_assign_34__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[34]), .Z(buf_def_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_assign_35__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[35]), .Z(buf_def_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_assign_35__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[35]), .Z(buf_def_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_assign_35__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[35]), .Z(buf_def_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_assign_35__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[35]), .Z(buf_def_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_assign_36__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[36]), .Z(buf_def_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_assign_36__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[36]), .Z(buf_def_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_assign_36__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[36]), .Z(buf_def_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_assign_36__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[36]), .Z(buf_def_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_assign_37__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[37]), .Z(buf_def_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_assign_37__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[37]), .Z(buf_def_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_assign_37__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[37]), .Z(buf_def_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_assign_37__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[37]), .Z(buf_def_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_assign_38__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[38]), .Z(buf_def_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_assign_38__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[38]), .Z(buf_def_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_assign_38__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[38]), .Z(buf_def_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_assign_38__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[38]), .Z(buf_def_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_assign_39__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[39]), .Z(buf_def_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_assign_39__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[39]), .Z(buf_def_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_assign_39__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[39]), .Z(buf_def_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_assign_39__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[39]), .Z(buf_def_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_assign_40__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[40]), .Z(buf_def_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_assign_40__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[40]), .Z(buf_def_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_assign_40__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[40]), .Z(buf_def_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_assign_40__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[40]), .Z(buf_def_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_assign_41__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[41]), .Z(buf_def_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_assign_41__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[41]), .Z(buf_def_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_assign_41__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[41]), .Z(buf_def_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_assign_41__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[41]), .Z(buf_def_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_assign_42__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[42]), .Z(buf_def_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_assign_42__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[42]), .Z(buf_def_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_assign_42__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[42]), .Z(buf_def_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_assign_42__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[42]), .Z(buf_def_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_assign_43__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[43]), .Z(buf_def_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_assign_43__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[43]), .Z(buf_def_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_assign_43__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[43]), .Z(buf_def_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_assign_43__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[43]), .Z(buf_def_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_assign_44__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[44]), .Z(buf_def_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_assign_44__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[44]), .Z(buf_def_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_assign_44__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[44]), .Z(buf_def_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_assign_44__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[44]), .Z(buf_def_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_assign_45__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[45]), .Z(buf_def_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_assign_45__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[45]), .Z(buf_def_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_assign_45__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[45]), .Z(buf_def_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_assign_45__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[45]), .Z(buf_def_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_assign_46__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[46]), .Z(buf_def_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_assign_46__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[46]), .Z(buf_def_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_assign_46__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[46]), .Z(buf_def_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_assign_46__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[46]), .Z(buf_def_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_assign_47__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[47]), .Z(buf_def_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_assign_47__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[47]), .Z(buf_def_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_assign_47__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[47]), .Z(buf_def_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_assign_47__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[47]), .Z(buf_def_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_assign_48__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[48]), .Z(buf_def_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_assign_48__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[48]), .Z(buf_def_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_assign_48__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[48]), .Z(buf_def_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_assign_48__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[48]), .Z(buf_def_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_assign_49__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[49]), .Z(buf_def_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_assign_49__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[49]), .Z(buf_def_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_assign_49__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[49]), .Z(buf_def_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_assign_49__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[49]), .Z(buf_def_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_assign_50__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[50]), .Z(buf_def_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_assign_50__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[50]), .Z(buf_def_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_assign_50__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[50]), .Z(buf_def_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_assign_50__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[50]), .Z(buf_def_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_assign_51__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[51]), .Z(buf_def_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_assign_51__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[51]), .Z(buf_def_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_assign_51__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[51]), .Z(buf_def_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_assign_51__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[51]), .Z(buf_def_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_assign_52__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[52]), .Z(buf_def_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_assign_52__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[52]), .Z(buf_def_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_assign_52__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[52]), .Z(buf_def_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_assign_52__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[52]), .Z(buf_def_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_assign_53__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[53]), .Z(buf_def_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_assign_53__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[53]), .Z(buf_def_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_assign_53__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[53]), .Z(buf_def_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_assign_53__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[53]), .Z(buf_def_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_assign_54__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[54]), .Z(buf_def_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_assign_54__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[54]), .Z(buf_def_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_assign_54__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[54]), .Z(buf_def_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_assign_54__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[54]), .Z(buf_def_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_assign_55__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[55]), .Z(buf_def_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_assign_55__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[55]), .Z(buf_def_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_assign_55__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[55]), .Z(buf_def_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_assign_55__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[55]), .Z(buf_def_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_assign_56__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[56]), .Z(buf_def_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_assign_56__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[56]), .Z(buf_def_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_assign_56__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[56]), .Z(buf_def_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_assign_56__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[56]), .Z(buf_def_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_assign_57__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[57]), .Z(buf_def_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_assign_57__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[57]), .Z(buf_def_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_assign_57__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[57]), .Z(buf_def_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_assign_57__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[57]), .Z(buf_def_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_assign_58__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[58]), .Z(buf_def_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_assign_58__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[58]), .Z(buf_def_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_assign_58__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[58]), .Z(buf_def_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_assign_58__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[58]), .Z(buf_def_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_assign_59__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[59]), .Z(buf_def_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_assign_59__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[59]), .Z(buf_def_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_assign_59__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[59]), .Z(buf_def_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_assign_59__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[59]), .Z(buf_def_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_assign_60__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[60]), .Z(buf_def_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_assign_60__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[60]), .Z(buf_def_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_assign_60__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[60]), .Z(buf_def_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_assign_60__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[60]), .Z(buf_def_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_assign_61__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[61]), .Z(buf_def_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_assign_61__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[61]), .Z(buf_def_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_assign_61__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[61]), .Z(buf_def_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_assign_61__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[61]), .Z(buf_def_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_assign_62__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[62]), .Z(buf_def_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_assign_62__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[62]), .Z(buf_def_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_assign_62__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[62]), .Z(buf_def_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_assign_62__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[62]), .Z(buf_def_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_assign_63__UI_BUF_o_data_bus_first ( .I(
        i_data_bus[63]), .Z(buf_def_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_assign_63__buf_level_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_0__i_data_o_buf[63]), .Z(buf_def_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_assign_63__buf_level_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_1__i_data_o_buf[63]), .Z(buf_def_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_assign_63__buf_level_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_def_2__i_data_o_buf[63]), .Z(buf_def_3__i_data_o_buf[63]) );
  DFQD4BWP30P140LVT o_valid_inner_reg ( .D(N84), .CP(clk), .Q(o_valid) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_31_ ( .D(N116), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_30_ ( .D(N115), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_29_ ( .D(N114), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_28_ ( .D(N113), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_27_ ( .D(N112), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_26_ ( .D(N111), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_25_ ( .D(N110), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_24_ ( .D(N109), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_23_ ( .D(N108), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_22_ ( .D(N107), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_21_ ( .D(N106), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_20_ ( .D(N105), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_19_ ( .D(N104), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_18_ ( .D(N103), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_17_ ( .D(N102), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_16_ ( .D(N101), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_15_ ( .D(N100), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_14_ ( .D(N99), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_13_ ( .D(N98), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_12_ ( .D(N97), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_11_ ( .D(N96), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_10_ ( .D(N95), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_9_ ( .D(N94), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_8_ ( .D(N93), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_7_ ( .D(N92), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_6_ ( .D(N91), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_5_ ( .D(N90), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_4_ ( .D(N89), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_3_ ( .D(N88), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_2_ ( .D(N87), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_1_ ( .D(N86), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140LVT o_data_bus_inner_reg_0_ ( .D(N85), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2D1BWP30P140LVT U40 ( .A1(n6), .A2(i_en), .ZN(n10) );
  NR3OPTPAD2BWP30P140LVT U41 ( .A1(n10), .A2(n9), .A3(i_valid[1]), .ZN(n5) );
  INVD2BWP30P140LVT U42 ( .I(n12), .ZN(n32) );
  XNR2UD1BWP30P140LVT U43 ( .A1(i_valid[1]), .A2(i_valid[0]), .ZN(n7) );
  INVD1BWP30P140LVT U44 ( .I(rst), .ZN(n6) );
  NR2D1BWP30P140LVT U45 ( .A1(n7), .A2(n10), .ZN(N84) );
  INVD1BWP30P140LVT U46 ( .I(n10), .ZN(n8) );
  INVD1BWP30P140LVT U47 ( .I(i_valid[0]), .ZN(n9) );
  AN3D1BWP30P140LVT U48 ( .A1(n8), .A2(i_valid[1]), .A3(n9), .Z(n12) );
  INVD1BWP30P140LVT U49 ( .I(buf_def_3__i_data_o_buf[32]), .ZN(n11) );
  MOAI22D1BWP30P140LVT U50 ( .A1(n32), .A2(n11), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[0]), .ZN(N85) );
  INVD1BWP30P140LVT U51 ( .I(buf_def_3__i_data_o_buf[33]), .ZN(n13) );
  MOAI22D1BWP30P140LVT U52 ( .A1(n32), .A2(n13), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[1]), .ZN(N86) );
  INVD1BWP30P140LVT U53 ( .I(buf_def_3__i_data_o_buf[34]), .ZN(n14) );
  MOAI22D1BWP30P140LVT U54 ( .A1(n32), .A2(n14), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[2]), .ZN(N87) );
  INVD1BWP30P140LVT U55 ( .I(buf_def_3__i_data_o_buf[35]), .ZN(n15) );
  MOAI22D1BWP30P140LVT U56 ( .A1(n32), .A2(n15), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[3]), .ZN(N88) );
  INVD1BWP30P140LVT U57 ( .I(buf_def_3__i_data_o_buf[36]), .ZN(n16) );
  MOAI22D1BWP30P140LVT U58 ( .A1(n32), .A2(n16), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[4]), .ZN(N89) );
  INVD1BWP30P140LVT U59 ( .I(buf_def_3__i_data_o_buf[37]), .ZN(n17) );
  MOAI22D1BWP30P140LVT U60 ( .A1(n32), .A2(n17), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[5]), .ZN(N90) );
  INVD1BWP30P140LVT U61 ( .I(buf_def_3__i_data_o_buf[38]), .ZN(n18) );
  MOAI22D1BWP30P140LVT U62 ( .A1(n32), .A2(n18), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[6]), .ZN(N91) );
  INVD1BWP30P140LVT U63 ( .I(buf_def_3__i_data_o_buf[39]), .ZN(n19) );
  MOAI22D1BWP30P140LVT U64 ( .A1(n32), .A2(n19), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[7]), .ZN(N92) );
  INVD1BWP30P140LVT U65 ( .I(buf_def_3__i_data_o_buf[40]), .ZN(n20) );
  MOAI22D1BWP30P140LVT U66 ( .A1(n32), .A2(n20), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[8]), .ZN(N93) );
  INVD1BWP30P140LVT U67 ( .I(buf_def_3__i_data_o_buf[41]), .ZN(n21) );
  MOAI22D1BWP30P140LVT U68 ( .A1(n32), .A2(n21), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[9]), .ZN(N94) );
  INVD1BWP30P140LVT U69 ( .I(buf_def_3__i_data_o_buf[42]), .ZN(n22) );
  MOAI22D1BWP30P140LVT U70 ( .A1(n32), .A2(n22), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[10]), .ZN(N95) );
  INVD1BWP30P140LVT U71 ( .I(buf_def_3__i_data_o_buf[43]), .ZN(n23) );
  MOAI22D1BWP30P140LVT U72 ( .A1(n32), .A2(n23), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[11]), .ZN(N96) );
  INVD1BWP30P140LVT U73 ( .I(buf_def_3__i_data_o_buf[44]), .ZN(n24) );
  MOAI22D1BWP30P140LVT U74 ( .A1(n32), .A2(n24), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[12]), .ZN(N97) );
  INVD1BWP30P140LVT U75 ( .I(buf_def_3__i_data_o_buf[45]), .ZN(n25) );
  MOAI22D1BWP30P140LVT U76 ( .A1(n32), .A2(n25), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[13]), .ZN(N98) );
  INVD1BWP30P140LVT U77 ( .I(buf_def_3__i_data_o_buf[46]), .ZN(n26) );
  MOAI22D1BWP30P140LVT U78 ( .A1(n32), .A2(n26), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[14]), .ZN(N99) );
  INVD1BWP30P140LVT U79 ( .I(buf_def_3__i_data_o_buf[47]), .ZN(n27) );
  MOAI22D1BWP30P140LVT U80 ( .A1(n32), .A2(n27), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[15]), .ZN(N100) );
  INVD1BWP30P140LVT U81 ( .I(buf_def_3__i_data_o_buf[48]), .ZN(n28) );
  MOAI22D1BWP30P140LVT U82 ( .A1(n32), .A2(n28), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[16]), .ZN(N101) );
  INVD1BWP30P140LVT U83 ( .I(buf_def_3__i_data_o_buf[49]), .ZN(n29) );
  MOAI22D1BWP30P140LVT U84 ( .A1(n32), .A2(n29), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[17]), .ZN(N102) );
  INVD1BWP30P140LVT U85 ( .I(buf_def_3__i_data_o_buf[50]), .ZN(n30) );
  MOAI22D1BWP30P140LVT U86 ( .A1(n32), .A2(n30), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[18]), .ZN(N103) );
  INVD1BWP30P140LVT U87 ( .I(buf_def_3__i_data_o_buf[51]), .ZN(n31) );
  MOAI22D1BWP30P140LVT U88 ( .A1(n32), .A2(n31), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[19]), .ZN(N104) );
  INVD1BWP30P140LVT U89 ( .I(buf_def_3__i_data_o_buf[52]), .ZN(n33) );
  MOAI22D1BWP30P140LVT U90 ( .A1(n32), .A2(n33), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[20]), .ZN(N105) );
  INVD1BWP30P140LVT U91 ( .I(buf_def_3__i_data_o_buf[53]), .ZN(n34) );
  MOAI22D1BWP30P140LVT U92 ( .A1(n32), .A2(n34), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[21]), .ZN(N106) );
  INVD1BWP30P140LVT U93 ( .I(buf_def_3__i_data_o_buf[54]), .ZN(n35) );
  MOAI22D1BWP30P140LVT U94 ( .A1(n32), .A2(n35), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[22]), .ZN(N107) );
  INVD1BWP30P140LVT U95 ( .I(buf_def_3__i_data_o_buf[55]), .ZN(n36) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n32), .A2(n36), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[23]), .ZN(N108) );
  INVD1BWP30P140LVT U97 ( .I(buf_def_3__i_data_o_buf[56]), .ZN(n37) );
  MOAI22D1BWP30P140LVT U98 ( .A1(n32), .A2(n37), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[24]), .ZN(N109) );
  INVD1BWP30P140LVT U99 ( .I(buf_def_3__i_data_o_buf[57]), .ZN(n38) );
  MOAI22D1BWP30P140LVT U100 ( .A1(n32), .A2(n38), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[25]), .ZN(N110) );
  INVD1BWP30P140LVT U101 ( .I(buf_def_3__i_data_o_buf[58]), .ZN(n39) );
  MOAI22D1BWP30P140LVT U102 ( .A1(n32), .A2(n39), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[26]), .ZN(N111) );
  INVD1BWP30P140LVT U103 ( .I(buf_def_3__i_data_o_buf[59]), .ZN(n40) );
  MOAI22D1BWP30P140LVT U104 ( .A1(n32), .A2(n40), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[27]), .ZN(N112) );
  INVD1BWP30P140LVT U105 ( .I(buf_def_3__i_data_o_buf[60]), .ZN(n41) );
  MOAI22D1BWP30P140LVT U106 ( .A1(n32), .A2(n41), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[28]), .ZN(N113) );
  INVD1BWP30P140LVT U107 ( .I(buf_def_3__i_data_o_buf[61]), .ZN(n42) );
  MOAI22D1BWP30P140LVT U108 ( .A1(n32), .A2(n42), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[29]), .ZN(N114) );
  INVD1BWP30P140LVT U109 ( .I(buf_def_3__i_data_o_buf[62]), .ZN(n43) );
  MOAI22D1BWP30P140LVT U110 ( .A1(n32), .A2(n43), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[30]), .ZN(N115) );
  INVD1BWP30P140LVT U111 ( .I(buf_def_3__i_data_o_buf[63]), .ZN(n44) );
  MOAI22D1BWP30P140LVT U112 ( .A1(n32), .A2(n44), .B1(n5), .B2(
        buf_def_3__i_data_o_buf[31]), .ZN(N116) );
endmodule

