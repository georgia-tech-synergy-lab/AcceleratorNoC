`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

//module controller_integrated(CLK, reset, boot_up, boot_up_local, boot_up_table_update, start, init_sram, direct_tap, table_parse, input_valid, glob_scen_noc_input_valid, delay_matrix_element, obj_id_element, scenario_update, hardware_latency1, hardware_latency2, scenario_len, data_in, final_out_0, final_out_1, final_out_2);//, final_out_3);

//module controller_integrated(CLK, reset, boot_up, boot_up_local, boot_up_table_update, start, init_sram, direct_tap, table_parse, input_valid, glob_scen_noc_input_valid, delay_matrix_element, obj_id_element, scenario_update, hardware_latency1, hardware_latency2, scenario_len, data_in, coe, interp_coe, sel1,sel2,sel3,sel4,output_real_with_multi_1, output_real_with_multi_2, output_real_with_multi_3, output_img_with_multi_1, output_img_with_multi_2, output_img_with_multi_3);

//module controller_integrated(CLK, reset, boot_up, boot_up_local, boot_up_table_update, start, init_sram, direct_tap, table_parse, input_valid, glob_scen_noc_input_valid, delay_matrix_element, obj_id_element, hardware_latency1, hardware_latency2, scenario_len, data_in, coe, interp_coe, sel1,sel2,sel3,sel4,out1_real,out1_img,out2_real,out2_img,out3_real,out3_img, din, scen_ch, doppler_dft_clk, scenario_update_input_block, input_block_latency, input_block_scen_pipeline, load_same_scenario, pe_controller_latency, interp_time_block_latency, doppler_time_block_latency,scenario_update_rx, input_latency, loc_controller_latency, ddnoc_latency,pre_cycle_doppler);

module controller_integrated(CLK, reset, boot_up_ext, boot_up_local_ext, boot_up_table_update_ext, start_ext, init_sram_ext, direct_tap, table_parse_ext, dft_clk_out, delay_matrix_element, obj_id_element, hardware_latency1, hardware_latency2, scenario_len, data_in, coe, interp_coe, sel1,sel2,out1_real,out1_img,out2_real,out2_img,out3_real,out3_img, din, doppler_dft_clk, scenario_update_input_block, scenario_update_input_block2,input_block_latency, input_block_scen_pipeline, load_same_scenario, pe_controller_latency, interp_time_block_latency, doppler_time_block_latency,scenario_update_rx, input_latency, loc_controller_latency, ddnoc_latency,pre_cycle_doppler,scenario_global_latency2, scenario_interp_latency2, dft_program_delay, scen_del_pe_config, scenario_del_global_internal_config);


    // parameter
    	parameter N_sample = 1024;
	parameter datawidth = 16;
	parameter address_vector_width = 4; //4; //can be 200 or 8: 8 for small tapeout
	parameter full_address_vector_width = 8; //4; //can be 200 or 8: 8 for small tapeout
	parameter N_obj = 4; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 4; // 16 local controllers in subscaled system
	parameter sample_address_width = 10; /// assuming 256 words: needs to change if arrangement is different
	parameter pe_sample_address_width = 8; /// assuming 256 words: needs to change if arrangement is different
	parameter packet_width = 2+2*datawidth + full_address_vector_width;
	parameter delay_length = 14; // log(id_width*N_sample)
	parameter obj_id_width = 2; // log(N_obj)
	parameter tapping_loc_packet_width = sample_address_width + obj_id_width; // log(N_obj)
	parameter scen_len_width = 14;   //needs to be revised
	parameter noc_output_half = 8;   //needs to be revised
	parameter num_loc_controller = 16;	
	parameter num_prefetch_config_width = 25;
	parameter latency_width = 7;

//=== IO Ports ===//

     // Normal Mode Input
    	input CLK; // system clock, generated by VCO
	input reset;
	input start_ext;
	input init_sram_ext;
	input direct_tap;
	input boot_up_ext;
	input boot_up_local_ext;
	input boot_up_table_update_ext;
	input table_parse_ext;
	//input input_valid;
	//input glob_scen_noc_input_valid;
	input dft_clk_out;
	input [delay_length - 1:0] delay_matrix_element;
	input [obj_id_width - 1:0] obj_id_element;
	input [delay_length - 1:0] hardware_latency1;   ///keep as config to be input through spi?
	input [delay_length - 1:0] hardware_latency2;   /// keep as config to be input through spi?
	input [scen_len_width - 1:0] scenario_len;   /// keep as config to be input through spi?
	input [2*datawidth - 1:0] data_in;   
	input [delay_length - 1:0] input_block_latency;
	input [delay_length - 1:0] input_block_scen_pipeline;
	input load_same_scenario;
	//input     sel1,sel2,sel3,sel4;
	input     sel1,sel2;
    	//input     [15:0] data_real1, data_img1,data_real2, data_img2,data_real3, data_img3;
    	input     [15:0] coe;
    	input     [9:0]  interp_coe;
	//output [2*datawidth-1:0] final_out_3;

	//input [15:0] ts_inc;
	//input scen_ch;
	input doppler_dft_clk;

	//input [15:0] din_0,din_1,din_2;
	input [15:0] din;
	input [latency_width - 1:0] scenario_global_latency2;
	input [latency_width - 1:0] scenario_interp_latency2;
	input [latency_width - 1:0] input_latency;
	input [latency_width - 1:0] loc_controller_latency;
	input [latency_width - 1:0] ddnoc_latency;
	input [latency_width - 1:0] pe_controller_latency;
	input [latency_width - 1:0] interp_time_block_latency;
	input [latency_width - 1:0] doppler_time_block_latency;
	input [latency_width - 1:0] scen_del_pe_config;
	input [latency_width - 1:0] scenario_del_global_internal_config;
	input [8:0] pre_cycle_doppler;
	input [5:0] dft_program_delay;


	output [15:0] out1_real,out1_img,out2_real,out2_img,out3_real,out3_img;

	output reg scenario_update_input_block;
	output scenario_update_input_block2;
	output scenario_update_rx;
    // output

	wire [2*datawidth-1:0] final_out_0;
	wire [2*datawidth-1:0] final_out_1;
	wire [2*datawidth-1:0] final_out_2;
    	wire [15:0] output_real_with_multi_1, output_real_with_multi_2, output_real_with_multi_3;
    	wire [15:0] output_img_with_multi_1, output_img_with_multi_2, output_img_with_multi_3;



	wire [address_vector_width - 1:0] from_glob_prefetch_dest;
	wire [sample_address_width - 1:0] from_glob_prefetch_start;
	wire [sample_address_width - 1:0] from_glob_prefetch_stop;
	wire [id_width - 1:0] local_controller_id;
	wire scenario_update_to_loc; 
	wire valid_bit;
	wire prefetch_enable;

        wire [2*datawidth-1:0] noc_out_0;   
        wire [2*datawidth-1:0] noc_out_1;   
        wire [2*datawidth-1:0] noc_out_2;   
        wire [2*datawidth-1:0] noc_out_3;   
        wire [2*datawidth-1:0] noc_out_4;   
        wire [2*datawidth-1:0] noc_out_5;   
        wire [2*datawidth-1:0] noc_out_6;   
        wire [2*datawidth-1:0] noc_out_7;    
        wire [2*datawidth-1:0] noc_out_8;   
        wire [2*datawidth-1:0] noc_out_9;   
        wire [2*datawidth-1:0] noc_out_10;   
        wire [2*datawidth-1:0] noc_out_11;   
        wire [2*datawidth-1:0] noc_out_12;   
        wire [2*datawidth-1:0] noc_out_13;   
        wire [2*datawidth-1:0] noc_out_14;   
        wire [2*datawidth-1:0] noc_out_15;   
	wire [noc_output_half - 1:0] from_noc_output_valid_0;
	wire [noc_output_half - 1:0] from_noc_output_valid_1;

//////////// internal status regs/signals //////////////////////////////////
	wire [2*datawidth - 1:0] h_tree_input_data;
	wire write_flag_0;


	wire boundary_next_0;
	wire boundary_next_1;
	wire boundary_next_2;
	wire boundary_next_3;
	wire boundary_next_4;
	wire boundary_next_5;
	wire boundary_next_6;
	wire boundary_next_7;
	wire boundary_next_8;
	wire boundary_next_9;
	wire boundary_next_10;
	wire boundary_next_11;
	wire boundary_next_12;
	wire boundary_next_13;
	wire boundary_next_14;
	wire boundary_next_15;

	wire [address_vector_width - 1:0] dest_address_0;
	wire [address_vector_width - 1:0] dest_address_1;
	wire [address_vector_width - 1:0] dest_address_2;
	wire [address_vector_width - 1:0] dest_address_3;
	wire [address_vector_width - 1:0] dest_address_4;
	wire [address_vector_width - 1:0] dest_address_5;
	wire [address_vector_width - 1:0] dest_address_6;
	wire [address_vector_width - 1:0] dest_address_7;
	wire [address_vector_width - 1:0] dest_address_8;
	wire [address_vector_width - 1:0] dest_address_9;
	wire [address_vector_width - 1:0] dest_address_10;
	wire [address_vector_width - 1:0] dest_address_11;
	wire [address_vector_width - 1:0] dest_address_12;
	wire [address_vector_width - 1:0] dest_address_13;
	wire [address_vector_width - 1:0] dest_address_14;
	wire [address_vector_width - 1:0] dest_address_15;

	wire [sample_address_width - 1:0] prefetch_stop_address_0;
	wire [sample_address_width - 1:0] prefetch_stop_address_1;
	wire [sample_address_width - 1:0] prefetch_stop_address_2;
	wire [sample_address_width - 1:0] prefetch_stop_address_3;
	wire [sample_address_width - 1:0] prefetch_stop_address_4;
	wire [sample_address_width - 1:0] prefetch_stop_address_5;
	wire [sample_address_width - 1:0] prefetch_stop_address_6;
	wire [sample_address_width - 1:0] prefetch_stop_address_7;
	wire [sample_address_width - 1:0] prefetch_stop_address_8;
	wire [sample_address_width - 1:0] prefetch_stop_address_9;
	wire [sample_address_width - 1:0] prefetch_stop_address_10;
	wire [sample_address_width - 1:0] prefetch_stop_address_11;
	wire [sample_address_width - 1:0] prefetch_stop_address_12;
	wire [sample_address_width - 1:0] prefetch_stop_address_13;
	wire [sample_address_width - 1:0] prefetch_stop_address_14;
	wire [sample_address_width - 1:0] prefetch_stop_address_15;

	wire [address_vector_width - 1:0] prefetch_dest_addr_0;
	wire [address_vector_width - 1:0] prefetch_dest_addr_1;
	wire [address_vector_width - 1:0] prefetch_dest_addr_2;
	wire [address_vector_width - 1:0] prefetch_dest_addr_3;
	wire [address_vector_width - 1:0] prefetch_dest_addr_4;
	wire [address_vector_width - 1:0] prefetch_dest_addr_5;
	wire [address_vector_width - 1:0] prefetch_dest_addr_6;
	wire [address_vector_width - 1:0] prefetch_dest_addr_7;
	wire [address_vector_width - 1:0] prefetch_dest_addr_8;
	wire [address_vector_width - 1:0] prefetch_dest_addr_9;
	wire [address_vector_width - 1:0] prefetch_dest_addr_10;
	wire [address_vector_width - 1:0] prefetch_dest_addr_11;
	wire [address_vector_width - 1:0] prefetch_dest_addr_12;
	wire [address_vector_width - 1:0] prefetch_dest_addr_13;
	wire [address_vector_width - 1:0] prefetch_dest_addr_14;
	wire [address_vector_width - 1:0] prefetch_dest_addr_15;

	wire prefetch_boundary_prev_0;
	wire prefetch_boundary_prev_1;
	wire prefetch_boundary_prev_2;
	wire prefetch_boundary_prev_3;
	wire prefetch_boundary_prev_4;
	wire prefetch_boundary_prev_5;
	wire prefetch_boundary_prev_6;
	wire prefetch_boundary_prev_7;
	wire prefetch_boundary_prev_8;
	wire prefetch_boundary_prev_9;
	wire prefetch_boundary_prev_10;
	wire prefetch_boundary_prev_11;
	wire prefetch_boundary_prev_12;
	wire prefetch_boundary_prev_13;
	wire prefetch_boundary_prev_14;
	wire prefetch_boundary_prev_15;


	wire [2*datawidth - 1:0] D_0;
	wire [2*datawidth - 1:0] D_1;
	wire [2*datawidth - 1:0] D_2;
	wire [2*datawidth - 1:0] D_3;
	wire [2*datawidth - 1:0] D_4;
	wire [2*datawidth - 1:0] D_5;
	wire [2*datawidth - 1:0] D_6;
	wire [2*datawidth - 1:0] D_7;
	wire [2*datawidth - 1:0] D_8;
	wire [2*datawidth - 1:0] D_9;
	wire [2*datawidth - 1:0] D_10;
	wire [2*datawidth - 1:0] D_11;
	wire [2*datawidth - 1:0] D_12;
	wire [2*datawidth - 1:0] D_13;
	wire [2*datawidth - 1:0] D_14;
	wire [2*datawidth - 1:0] D_15;

        wire [packet_width-1:0] packet_out_0;   
        wire [packet_width-1:0] packet_out_1;   
        wire [packet_width-1:0] packet_out_2;   
        wire [packet_width-1:0] packet_out_3;   
        wire [packet_width-1:0] packet_out_4;   
        wire [packet_width-1:0] packet_out_5;   
        wire [packet_width-1:0] packet_out_6;   
        wire [packet_width-1:0] packet_out_7;   
        wire [packet_width-1:0] packet_out_8;   
        wire [packet_width-1:0] packet_out_9;   
        wire [packet_width-1:0] packet_out_10;   
        wire [packet_width-1:0] packet_out_11;   
        wire [packet_width-1:0] packet_out_12;   
        wire [packet_width-1:0] packet_out_13;   
        wire [packet_width-1:0] packet_out_14;   
        wire [packet_width-1:0] packet_out_15;   

////////// to be removed ///////////////////////

	wire write_boundary_next_0;
	wire write_boundary_next_1;
	wire write_boundary_next_2;
	wire write_boundary_next_3;
	wire write_boundary_next_4;
	wire write_boundary_next_5;
	wire write_boundary_next_6;
	wire write_boundary_next_7;
	wire write_boundary_next_8;
	wire write_boundary_next_9;
	wire write_boundary_next_10;
	wire write_boundary_next_11;
	wire write_boundary_next_12;
	wire write_boundary_next_13;
	wire write_boundary_next_14;
	wire write_boundary_next_15;

	wire ready;

	wire [noc_output_half-1:0] from_loc_controller_data_valid_0;
	wire [noc_output_half-1:0] from_loc_controller_data_valid_1;
	wire [2*datawidth*noc_output_half - 1: 0] from_local_controller_data_bus_0;
	wire [2*datawidth*noc_output_half- 1: 0] from_local_controller_data_bus_1;
	wire [2*datawidth*noc_output_half - 1:0] from_noc_output_data_0;
	wire [2*datawidth*noc_output_half - 1:0] from_noc_output_data_1;
	wire [full_address_vector_width*noc_output_half - 1:0] from_local_controller_dest_addr_0;
	wire [full_address_vector_width*noc_output_half - 1:0] from_local_controller_dest_addr_1;
	wire [num_loc_controller - 1:0] from_glob_prefetch_valid;
	wire [num_loc_controller*num_prefetch_config_width - 1:0] from_glob_prefetch_start_stop_dest_en;
	wire [11:0] htree_connected_addr;  //no of bits needs to be fixed once Htree is fixed

	wire scenario_update_input_block_l1;
	reg scenario_update_input_block_l2;
	reg scenario_update_input_block_l3;
	reg scenario_update_input_block_l4;
	reg scenario_update_input_block_l5;
	reg scenario_update_input_block_l6;
	wire scenario_update_interp;
	wire scenario_update_interp2;
	wire scenario_update_doppler_real;

	wire start;
	wire init_sram;
	wire boot_up;
	wire boot_up_local;
	wire boot_up_table_update;
	wire table_parse;


////////////////////// NoC interface ////////////////////////////////////////
	assign from_loc_controller_data_valid_0 = {packet_out_7[41], packet_out_6[41], packet_out_5[41], packet_out_4[41], packet_out_3[41], packet_out_2[41], packet_out_1[41], packet_out_0[41]};
	assign from_loc_controller_data_valid_1 = {packet_out_15[41], packet_out_14[41], packet_out_13[41], packet_out_12[41], packet_out_11[41], packet_out_10[41], packet_out_9[41], packet_out_8[41]};


	assign from_local_controller_data_bus_0 = {packet_out_7[39:8], packet_out_6[39:8], packet_out_5[39:8], packet_out_4[39:8], packet_out_3[39:8], packet_out_2[39:8], packet_out_1[39:8], packet_out_0[39:8]};
	assign from_local_controller_data_bus_1 = {packet_out_15[39:8], packet_out_14[39:8], packet_out_13[39:8], packet_out_12[39:8], packet_out_11[39:8], packet_out_10[39:8], packet_out_9[39:8], packet_out_8[39:8]};

	assign from_local_controller_dest_addr_0 = {packet_out_7[7:0], packet_out_6[7:0], packet_out_5[7:0], packet_out_4[7:0], packet_out_3[7:0], packet_out_2[7:0], packet_out_1[7:0], packet_out_0[7:0]};
	assign from_local_controller_dest_addr_1 = {packet_out_15[7:0], packet_out_14[7:0], packet_out_13[7:0], packet_out_12[7:0], packet_out_11[7:0], packet_out_10[7:0], packet_out_9[7:0], packet_out_8[7:0]};


	


	assign noc_out_0 = from_noc_output_data_0[31:0];
	assign noc_out_1 = from_noc_output_data_0[63:32];
	assign noc_out_2 = from_noc_output_data_0[95:64];
	assign noc_out_3 = from_noc_output_data_0[127:96];
	assign noc_out_4 = from_noc_output_data_0[159:128];
	assign noc_out_5 = from_noc_output_data_0[191:160];
	assign noc_out_6 = from_noc_output_data_0[223:192];
	assign noc_out_7 = from_noc_output_data_0[255:224];
	assign noc_out_8 = from_noc_output_data_1[31:0];
	assign noc_out_9 = from_noc_output_data_1[63:32];
	assign noc_out_10 = from_noc_output_data_1[95:64];
	assign noc_out_11 = from_noc_output_data_1[127:96];
	assign noc_out_12 = from_noc_output_data_1[159:128];
	assign noc_out_13 = from_noc_output_data_1[191:160];
	assign noc_out_14 = from_noc_output_data_1[223:192];
	assign noc_out_15 = from_noc_output_data_1[255:224];


	always @(posedge CLK) begin
		if (reset) begin
			scenario_update_input_block_l2 <= 0;
			scenario_update_input_block_l3 <= 0;
			scenario_update_input_block_l4 <= 0;
			scenario_update_input_block_l5 <= 0;
			scenario_update_input_block_l6 <= 0;
			scenario_update_input_block <= 0;
		end		
		else begin
			scenario_update_input_block_l2 <= scenario_update_input_block_l1;
			scenario_update_input_block_l3 <= scenario_update_input_block_l2;
			scenario_update_input_block_l4 <= scenario_update_input_block_l3;
			scenario_update_input_block_l5 <= scenario_update_input_block_l4;
			scenario_update_input_block_l6 <= scenario_update_input_block_l5;
			scenario_update_input_block <= scenario_update_input_block_l6;
		end		



	end



////// GLOBAL CONTROLLER//////////
    //global_controller DUT_global_controller(.CLK(CLK), .reset(reset), .start(start), .boot_up(boot_up), .boot_up_table_update(boot_up_table_update), .table_parse(table_parse), .input_valid(input_valid), .glob_scen_noc_input_valid(glob_scen_noc_input_valid), .delay_matrix_element(delay_matrix_element), .obj_id_element(obj_id_element),.from_glob_prefetch_start(from_glob_prefetch_start),.from_glob_prefetch_dest(from_glob_prefetch_dest),  .scenario_update(scenario_update_global), .local_controller_id(local_controller_id), .tapping_loc_packet(tapping_loc_packet), .from_glob_prefetch_stop(from_glob_prefetch_stop), .hardware_latency1(hardware_latency1), .hardware_latency2(hardware_latency2), .scenario_len(scenario_len), .prefetch_bypass_dest_addr_int(prefetch_bypass_dest_addr_int), .prefetch_bypass_cycles(prefetch_bypass_cycles), .prefetch_bypass_start_addr(prefetch_bypass_start_addr), .addr(addr), .data_in(data_in), .h_tree_input_data(h_tree_input_data), .h_tree_input_addr(h_tree_input_addr), .prefetch_bypass_path_input_data(prefetch_bypass_path_input_data), .prefetch_bypass_path_input_addr(prefetch_bypass_path_input_addr), .prefetch_bypass_valid(prefetch_bypass_valid), .prefetch_bypass_reqd(prefetch_bypass_reqd), .ready(ready), .scenario_counter(scenario_counter), .scenario_update_loc(scenario_update_to_loc), .scenario_update_global(scenario_update_global), .valid_bit(valid_bit), .prefetch_enable(prefetch_enable), .tapping_loc_valid(tapping_loc_valid),  .real_bypass_dest_addr_int(real_bypass_dest_addr_int), .real_bypass_reqd(real_bypass_reqd), .real_bypass_tap_loc(real_bypass_tap_loc), .real_bypass_path_input_data(real_bypass_path_input_data), .real_bypass_path_input_addr(real_bypass_path_input_addr), .real_bypass_valid(real_bypass_valid), .real_bypass_tap_loc_valid(real_bypass_tap_loc_valid));


	//glob_pe_controller DUT_glob_pe_controller(.CLK(CLK), .reset(reset), .boot_up(boot_up), .boot_up_local(boot_up_local), .boot_up_table_update(boot_up_table_update), .start(start), .init_sram(init_sram), .table_parse(table_parse), .input_valid(input_valid), .glob_scen_noc_input_valid(glob_scen_noc_input_valid), .delay_matrix_element(delay_matrix_element), .obj_id_element(obj_id_element), .from_glob_prefetch_start(from_glob_prefetch_start),  .from_glob_prefetch_dest(from_glob_prefetch_dest), .local_controller_id(local_controller_id), .from_glob_prefetch_stop(from_glob_prefetch_stop), .hardware_latency1(hardware_latency1), .hardware_latency2(hardware_latency2), .scenario_len(scenario_len), .data_in(data_in), .noc_out_0(noc_out_0), .noc_out_1(noc_out_1), .noc_out_2(noc_out_2), .noc_out_3(noc_out_3), .noc_out_4(noc_out_4), .noc_out_5(noc_out_5), .noc_out_6(noc_out_6), .noc_out_7(noc_out_7), .noc_out_8(noc_out_8), .noc_out_9(noc_out_9), .noc_out_10(noc_out_10), .noc_out_11(noc_out_11), .noc_out_12(noc_out_12), .noc_out_13(noc_out_13), .noc_out_14(noc_out_14), .noc_out_15(noc_out_15), .final_out_0(final_out_0), .final_out_1(final_out_1), .final_out_2(final_out_2), .valid_bit(valid_bit), .h_tree_input_data(h_tree_input_data), .htree_connected_addr(htree_connected_addr), .from_noc_output_valid_0(from_noc_output_valid_0), .from_noc_output_valid_1(from_noc_output_valid_1), .scenario_update_to_loc(scenario_update_to_loc), .prefetch_enable(prefetch_enable), .direct_tap(direct_tap), .ready(ready), .input_block_latency(input_block_latency), .scenario_update_global(scenario_update_input_block_l1), .load_same_scenario(load_same_scenario), .input_block_scen_pipeline(input_block_scen_pipeline), .pe_controller_latency(pe_controller_latency), .interp_time_block_latency(interp_time_block_latency), .doppler_time_block_latency(doppler_time_block_latency), .scenario_update_interp(scenario_update_interp), .scenario_update_doppler(scenario_update_doppler), .scenario_update_rx(scenario_update_rx), .input_latency(input_latency), .loc_controller_latency(loc_controller_latency), .ddnoc_latency(ddnoc_latency), .scenario_update_doppler_real(scenario_update_doppler_real), .pre_cycle_doppler(pre_cycle_doppler));
	glob_pe_controller DUT_glob_pe_controller(.CLK(CLK), .reset(reset), .boot_up_ext(boot_up_ext), .boot_up_local_ext(boot_up_local_ext), .boot_up_table_update_ext(boot_up_table_update_ext), .start_ext(start_ext), .init_sram_ext(init_sram_ext), .table_parse_ext(table_parse_ext), .dft_clk_out(dft_clk_out), .delay_matrix_element(delay_matrix_element), .obj_id_element(obj_id_element), .from_glob_prefetch_start(from_glob_prefetch_start),  .from_glob_prefetch_dest(from_glob_prefetch_dest), .local_controller_id(local_controller_id), .from_glob_prefetch_stop(from_glob_prefetch_stop), .hardware_latency1(hardware_latency1), .hardware_latency2(hardware_latency2), .scenario_len(scenario_len), .data_in(data_in), .noc_out_0(noc_out_0), .noc_out_1(noc_out_1), .noc_out_2(noc_out_2), .noc_out_3(noc_out_3), .noc_out_4(noc_out_4), .noc_out_5(noc_out_5), .noc_out_6(noc_out_6), .noc_out_7(noc_out_7), .noc_out_8(noc_out_8), .noc_out_9(noc_out_9), .noc_out_10(noc_out_10), .noc_out_11(noc_out_11), .noc_out_12(noc_out_12), .noc_out_13(noc_out_13), .noc_out_14(noc_out_14), .noc_out_15(noc_out_15), .final_out_0(final_out_0), .final_out_1(final_out_1), .final_out_2(final_out_2), .valid_bit(valid_bit), .h_tree_input_data(h_tree_input_data), .htree_connected_addr(htree_connected_addr), .from_noc_output_valid_0(from_noc_output_valid_0), .from_noc_output_valid_1(from_noc_output_valid_1), .scenario_update_to_loc(scenario_update_to_loc), .prefetch_enable(prefetch_enable), .direct_tap(direct_tap), .ready(ready), .input_block_latency(input_block_latency), .scenario_update_global(scenario_update_input_block_l1), .scenario_update_global2(scenario_update_input_block2), .load_same_scenario(load_same_scenario), .input_block_scen_pipeline(input_block_scen_pipeline), .pe_controller_latency(pe_controller_latency), .interp_time_block_latency(interp_time_block_latency), .doppler_time_block_latency(doppler_time_block_latency), .scenario_update_interp(scenario_update_interp), .scenario_update_doppler(scenario_update_doppler), .scenario_update_rx(scenario_update_rx), .input_latency(input_latency), .loc_controller_latency(loc_controller_latency), .ddnoc_latency(ddnoc_latency), .scenario_update_doppler_real(scenario_update_doppler_real), .pre_cycle_doppler(pre_cycle_doppler), .scenario_global_latency2(scenario_global_latency2), .scenario_update_interp2(scenario_update_interp2), .scenario_interp_latency2(scenario_interp_latency2), .boot_up(boot_up), .boot_up_local(boot_up_local), .boot_up_table_update(boot_up_table_update), .start(start), .init_sram(init_sram), .table_parse(table_parse), .dft_program_delay(dft_program_delay), .scen_del_pe_config(scen_del_pe_config), .scenario_del_global_internal_config(scenario_del_global_internal_config));

//////// interpolation ///////////////

       combine_top_level_with_o_addertree_1 DUT_interp( .data_real1(final_out_0[31:16]), .data_img1(final_out_0[15:0]), .data_real2(final_out_1[31:16]), .data_img2(final_out_1[15:0]), .data_real3(final_out_2[31:16]), .data_img3(final_out_2[15:0]), .coe(coe), .interp_coe(interp_coe), .CLK(CLK), .sel1(sel1), .sel2(sel2), .sel3(scenario_update_interp), .sel4(scenario_update_interp2), .Reset(reset), .output_real_with_multi_1(output_real_with_multi_1), .output_real_with_multi_2(output_real_with_multi_2), .output_real_with_multi_3(output_real_with_multi_3), .output_img_with_multi_1(output_img_with_multi_1), .output_img_with_multi_2(output_img_with_multi_2), .output_img_with_multi_3(output_img_with_multi_3));




///////////////////// Doppler module /////////////////////////

	//top_mod_cm_1 DUT_doppler(.CLK(CLK), .scen_ch(scen_ch), .reset(reset), .ts_inc(ts_inc), .din_0(din_0), .din_1(din_1), .din_2(din_2), .int1_real(output_real_with_multi_1), .int1_img(output_img_with_multi_1), .int2_real(output_real_with_multi_2), .int2_img(output_img_with_multi_2), .int3_real(output_real_with_multi_3), .int3_img(output_img_with_multi_3), .out1_real(out1_real), .out1_img(out1_img), .out2_real(out2_real), .out2_img(out2_img), .out3_real(out3_real), .out3_img(out3_img));

	top_mod_cm_1 DUT_doppler( .doppler_dft_clk(doppler_dft_clk), .CLK(CLK), .scen_ch(scenario_update_doppler_real), .reset(reset), .din(din), .int1_real(output_real_with_multi_1), .int1_img(output_img_with_multi_1), .int2_real(output_real_with_multi_2), .int2_img(output_img_with_multi_2), .int3_real(output_real_with_multi_3), .int3_img(output_img_with_multi_3), .out1_real(out1_real), .out1_img(out1_img), .out2_real(out2_real), .out2_img(out2_img), .out3_real(out3_real), .out3_img(out3_img) );


////////// H TREE //////////////
    Htree_Flat_clockedHiFeq_16 DUT_htree( .CLK(CLK), .addr(htree_connected_addr), .en(ready), .data_in(h_tree_input_data),  .en_sub_0(write_flag_0),  .data_in_sub_0(D_0), .data_in_sub_1(D_1), .data_in_sub_2(D_2), .data_in_sub_3(D_3),  .data_in_sub_4(D_4), .data_in_sub_5(D_5), .data_in_sub_6(D_6), .data_in_sub_7(D_7),  .data_in_sub_8(D_8), .data_in_sub_9(D_9), .data_in_sub_10(D_10), .data_in_sub_11(D_11), .data_in_sub_12(D_12), .data_in_sub_13(D_13), .data_in_sub_14(D_14), .data_in_sub_15(D_15) );

/////////// DDNOC////////////
 crossbar_one_hot_seq DUT_ddnoc_0(.CLK(CLK), .rst(reset), .i_valid(from_loc_controller_data_valid_0), .i_data_bus(from_local_controller_data_bus_0), .o_valid(from_noc_output_valid_0), .o_data_bus(from_noc_output_data_0), .i_en(ready), .i_cmd(from_local_controller_dest_addr_0) );
 
crossbar_one_hot_seq DUT_ddnoc_1(.CLK(CLK), .rst(reset), .i_valid(from_loc_controller_data_valid_1), .i_data_bus(from_local_controller_data_bus_1), .o_valid(from_noc_output_valid_1), .o_data_bus(from_noc_output_data_1), .i_en(ready), .i_cmd(from_local_controller_dest_addr_1) );

///////////PE CONTROLLER //////



////////////// LINEAR NOC FROM GLOBAL CONTROLLER TO LOCAL CONTROLLER ///////

 linear_network_unicast_seq_1_16 DUT_linNoc_1_16(.CLK(CLK), .rst(reset), .i_valid(valid_bit), .i_data_bus({from_glob_prefetch_start,from_glob_prefetch_stop,from_glob_prefetch_dest,prefetch_enable}), .o_valid(from_glob_prefetch_valid), .o_data_bus(from_glob_prefetch_start_stop_dest_en), .i_en(1'b1), .i_cmd(local_controller_id) );



///////// LOCAL CONTROLLER ///////// 
    local_controller_prefetch_full DUT_local_controller_0(.CLK(CLK), .reset(reset), .boot_up(boot_up_local), .start(start),     .input_boundary_flag(boundary_next_15), .prev_dest_address(dest_address_15),.packet_out(packet_out_0), .boundary_next(boundary_next_0), .dest_address(dest_address_0), .D(D_0),.write_flag(write_flag_0), .from_glob_prefetch_valid(from_glob_prefetch_valid[0]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[24:15]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[14:5]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[4:1]),  .write_boundary_next(write_boundary_next_0), .input_write_boundary(write_boundary_next_15), .prefetch_next_dest_addr(prefetch_dest_addr_1), .prefetch_next_stop_address(prefetch_stop_address_1), .prefetch_boundary_prev(prefetch_boundary_prev_0), .input_prefetch_boundary_flag(prefetch_boundary_prev_1), .prefetch_stop_address(prefetch_stop_address_0), .prefetch_dest_addr(prefetch_dest_addr_0),.scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[0]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_1(.CLK(CLK), .reset(reset),  .boot_up(boot_up_local), .start(start),     .input_boundary_flag(boundary_next_0), .prev_dest_address(dest_address_0), .packet_out(packet_out_1), .boundary_next(boundary_next_1), .dest_address(dest_address_1), .D(D_1),  .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[1]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[49:40]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[39:30]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[29:26]),   .write_boundary_next(write_boundary_next_1), .input_write_boundary(write_boundary_next_0), .prefetch_next_dest_addr(prefetch_dest_addr_2), .prefetch_next_stop_address(prefetch_stop_address_2), .prefetch_boundary_prev(prefetch_boundary_prev_1), .input_prefetch_boundary_flag(prefetch_boundary_prev_2), .prefetch_stop_address(prefetch_stop_address_1), .prefetch_dest_addr(prefetch_dest_addr_1), .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[25]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_2(.CLK(CLK), .reset(reset),  .boot_up(boot_up_local), .start(start),    .input_boundary_flag(boundary_next_1), .prev_dest_address(dest_address_1), .packet_out(packet_out_2), .boundary_next(boundary_next_2), .dest_address(dest_address_2), .D(D_2), .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[2]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[74:65]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[64:55]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[54:51]),  .write_boundary_next(write_boundary_next_2), .input_write_boundary(write_boundary_next_1), .prefetch_next_dest_addr(prefetch_dest_addr_3), .prefetch_next_stop_address(prefetch_stop_address_3), .prefetch_boundary_prev(prefetch_boundary_prev_2), .input_prefetch_boundary_flag(prefetch_boundary_prev_3), .prefetch_stop_address(prefetch_stop_address_2), .prefetch_dest_addr(prefetch_dest_addr_2),  .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[50]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_3(.CLK(CLK), .reset(reset),  .boot_up(boot_up_local), .start(start),   .input_boundary_flag(boundary_next_2), .prev_dest_address(dest_address_2),  .packet_out(packet_out_3), .boundary_next(boundary_next_3), .dest_address(dest_address_3), .D(D_3),  .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[3]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[99:90]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[89:80]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[79:76]),  .write_boundary_next(write_boundary_next_3), .input_write_boundary(write_boundary_next_2), .prefetch_next_dest_addr(prefetch_dest_addr_4), .prefetch_next_stop_address(prefetch_stop_address_4), .prefetch_boundary_prev(prefetch_boundary_prev_3), .input_prefetch_boundary_flag(prefetch_boundary_prev_4), .prefetch_stop_address(prefetch_stop_address_3), .prefetch_dest_addr(prefetch_dest_addr_3),  .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[75]), .init_sram(init_sram));


///////////////////////////////////////////////////////////



    local_controller_prefetch_full DUT_local_controller_4(.CLK(CLK), .reset(reset), .boot_up(boot_up_local), .start(start),     .input_boundary_flag(boundary_next_3), .prev_dest_address(dest_address_3),.packet_out(packet_out_4), .boundary_next(boundary_next_4), .dest_address(dest_address_4), .D(D_4),.write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[4]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[124:115]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[114:105]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[104:101]),  .write_boundary_next(write_boundary_next_4), .input_write_boundary(write_boundary_next_3), .prefetch_next_dest_addr(prefetch_dest_addr_5), .prefetch_next_stop_address(prefetch_stop_address_5), .prefetch_boundary_prev(prefetch_boundary_prev_4), .input_prefetch_boundary_flag(prefetch_boundary_prev_5), .prefetch_stop_address(prefetch_stop_address_4), .prefetch_dest_addr(prefetch_dest_addr_4),.scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[100]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_5(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),     .input_boundary_flag(boundary_next_4), .prev_dest_address(dest_address_4), .packet_out(packet_out_5), .boundary_next(boundary_next_5), .dest_address(dest_address_5), .D(D_5),  .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[5]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[149:140]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[139:130]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[129:126]),   .write_boundary_next(write_boundary_next_5), .input_write_boundary(write_boundary_next_4), .prefetch_next_dest_addr(prefetch_dest_addr_6), .prefetch_next_stop_address(prefetch_stop_address_6), .prefetch_boundary_prev(prefetch_boundary_prev_5), .input_prefetch_boundary_flag(prefetch_boundary_prev_6), .prefetch_stop_address(prefetch_stop_address_5), .prefetch_dest_addr(prefetch_dest_addr_5), .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[125]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_6(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),    .input_boundary_flag(boundary_next_5), .prev_dest_address(dest_address_5), .packet_out(packet_out_6), .boundary_next(boundary_next_6), .dest_address(dest_address_6), .D(D_6), .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[6]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[174:165]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[164:155]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[154:151]), .write_boundary_next(write_boundary_next_6), .input_write_boundary(write_boundary_next_5), .prefetch_next_dest_addr(prefetch_dest_addr_7), .prefetch_next_stop_address(prefetch_stop_address_7), .prefetch_boundary_prev(prefetch_boundary_prev_6), .input_prefetch_boundary_flag(prefetch_boundary_prev_7), .prefetch_stop_address(prefetch_stop_address_6), .prefetch_dest_addr(prefetch_dest_addr_6),  .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[150]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_7(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),   .input_boundary_flag(boundary_next_6), .prev_dest_address(dest_address_6),  .packet_out(packet_out_7), .boundary_next(boundary_next_7), .dest_address(dest_address_7), .D(D_7),  .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[7]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[199:190]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[189:180]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[179:176]),  .write_boundary_next(write_boundary_next_7), .input_write_boundary(write_boundary_next_6), .prefetch_next_dest_addr(prefetch_dest_addr_8), .prefetch_next_stop_address(prefetch_stop_address_8), .prefetch_boundary_prev(prefetch_boundary_prev_7), .input_prefetch_boundary_flag(prefetch_boundary_prev_8), .prefetch_stop_address(prefetch_stop_address_7), .prefetch_dest_addr(prefetch_dest_addr_7),  .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[175]), .init_sram(init_sram));

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

    local_controller_prefetch_full DUT_local_controller_8(.CLK(CLK), .reset(reset), .boot_up(boot_up_local), .start(start),     .input_boundary_flag(boundary_next_7), .prev_dest_address(dest_address_7),.packet_out(packet_out_8), .boundary_next(boundary_next_8), .dest_address(dest_address_8), .D(D_8),.write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[8]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[224:215]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[214:205]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[204:201]),  .write_boundary_next(write_boundary_next_8), .input_write_boundary(write_boundary_next_7), .prefetch_next_dest_addr(prefetch_dest_addr_9), .prefetch_next_stop_address(prefetch_stop_address_9), .prefetch_boundary_prev(prefetch_boundary_prev_8), .input_prefetch_boundary_flag(prefetch_boundary_prev_9), .prefetch_stop_address(prefetch_stop_address_8), .prefetch_dest_addr(prefetch_dest_addr_8),.scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[200]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_9(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),     .input_boundary_flag(boundary_next_8), .prev_dest_address(dest_address_8), .packet_out(packet_out_9), .boundary_next(boundary_next_9), .dest_address(dest_address_9), .D(D_9),  .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[9]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[249:240]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[239:230]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[229:226]),   .write_boundary_next(write_boundary_next_9), .input_write_boundary(write_boundary_next_8), .prefetch_next_dest_addr(prefetch_dest_addr_10), .prefetch_next_stop_address(prefetch_stop_address_10), .prefetch_boundary_prev(prefetch_boundary_prev_9), .input_prefetch_boundary_flag(prefetch_boundary_prev_10), .prefetch_stop_address(prefetch_stop_address_9), .prefetch_dest_addr(prefetch_dest_addr_9), .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[225]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_10(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),    .input_boundary_flag(boundary_next_9), .prev_dest_address(dest_address_9), .packet_out(packet_out_10), .boundary_next(boundary_next_10), .dest_address(dest_address_10), .D(D_10), .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[10]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[274:265]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[264:255]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[254:251]),  .write_boundary_next(write_boundary_next_10), .input_write_boundary(write_boundary_next_9), .prefetch_next_dest_addr(prefetch_dest_addr_11), .prefetch_next_stop_address(prefetch_stop_address_11), .prefetch_boundary_prev(prefetch_boundary_prev_10), .input_prefetch_boundary_flag(prefetch_boundary_prev_11), .prefetch_stop_address(prefetch_stop_address_10), .prefetch_dest_addr(prefetch_dest_addr_10),  .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[250]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_11(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),   .input_boundary_flag(boundary_next_10), .prev_dest_address(dest_address_10),  .packet_out(packet_out_11), .boundary_next(boundary_next_11), .dest_address(dest_address_11), .D(D_11),  .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[11]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[299:290]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[289:280]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[279:276]),  .write_boundary_next(write_boundary_next_11), .input_write_boundary(write_boundary_next_10), .prefetch_next_dest_addr(prefetch_dest_addr_12), .prefetch_next_stop_address(prefetch_stop_address_12), .prefetch_boundary_prev(prefetch_boundary_prev_11), .input_prefetch_boundary_flag(prefetch_boundary_prev_12), .prefetch_stop_address(prefetch_stop_address_11), .prefetch_dest_addr(prefetch_dest_addr_11),  .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[275]), .init_sram(init_sram));


///////////////////////////////////////////////////////////



    local_controller_prefetch_full DUT_local_controller_12(.CLK(CLK), .reset(reset), .boot_up(boot_up_local), .start(start),     .input_boundary_flag(boundary_next_11), .prev_dest_address(dest_address_11),.packet_out(packet_out_12), .boundary_next(boundary_next_12), .dest_address(dest_address_12), .D(D_12),.write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[12]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[324:315]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[314:305]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[304:301]),  .write_boundary_next(write_boundary_next_12), .input_write_boundary(write_boundary_next_11), .prefetch_next_dest_addr(prefetch_dest_addr_13), .prefetch_next_stop_address(prefetch_stop_address_13), .prefetch_boundary_prev(prefetch_boundary_prev_12), .input_prefetch_boundary_flag(prefetch_boundary_prev_13), .prefetch_stop_address(prefetch_stop_address_12), .prefetch_dest_addr(prefetch_dest_addr_12),.scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[300]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_13(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),     .input_boundary_flag(boundary_next_12), .prev_dest_address(dest_address_12), .packet_out(packet_out_13), .boundary_next(boundary_next_13), .dest_address(dest_address_13), .D(D_13),  .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[13]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[349:340]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[339:330]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[329:326]),   .write_boundary_next(write_boundary_next_13), .input_write_boundary(write_boundary_next_12), .prefetch_next_dest_addr(prefetch_dest_addr_14), .prefetch_next_stop_address(prefetch_stop_address_14), .prefetch_boundary_prev(prefetch_boundary_prev_13), .input_prefetch_boundary_flag(prefetch_boundary_prev_14), .prefetch_stop_address(prefetch_stop_address_13), .prefetch_dest_addr(prefetch_dest_addr_13), .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[325]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_14(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),    .input_boundary_flag(boundary_next_13), .prev_dest_address(dest_address_13), .packet_out(packet_out_14), .boundary_next(boundary_next_14), .dest_address(dest_address_14), .D(D_14), .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[14]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[374:365]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[364:355]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[354:351]), .write_boundary_next(write_boundary_next_14), .input_write_boundary(write_boundary_next_13), .prefetch_next_dest_addr(prefetch_dest_addr_15), .prefetch_next_stop_address(prefetch_stop_address_15), .prefetch_boundary_prev(prefetch_boundary_prev_14), .input_prefetch_boundary_flag(prefetch_boundary_prev_15), .prefetch_stop_address(prefetch_stop_address_14), .prefetch_dest_addr(prefetch_dest_addr_14),  .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[350]), .init_sram(init_sram));

    local_controller_prefetch_full DUT_local_controller_15(.CLK(CLK), .reset(reset),   .boot_up(boot_up_local), .start(start),   .input_boundary_flag(boundary_next_14), .prev_dest_address(dest_address_14),  .packet_out(packet_out_15), .boundary_next(boundary_next_15), .dest_address(dest_address_15), .D(D_15),  .write_flag(1'b0), .from_glob_prefetch_valid(from_glob_prefetch_valid[15]), .from_glob_prefetch_start(from_glob_prefetch_start_stop_dest_en[399:390]), .from_glob_prefetch_stop(from_glob_prefetch_start_stop_dest_en[389:380]), .from_glob_prefetch_dest(from_glob_prefetch_start_stop_dest_en[379:376]),  .write_boundary_next(write_boundary_next_15), .input_write_boundary(write_boundary_next_14), .prefetch_next_dest_addr(prefetch_dest_addr_0), .prefetch_next_stop_address(prefetch_stop_address_0), .prefetch_boundary_prev(prefetch_boundary_prev_15), .input_prefetch_boundary_flag(prefetch_boundary_prev_0), .prefetch_stop_address(prefetch_stop_address_15), .prefetch_dest_addr(prefetch_dest_addr_15),  .scenario_update(scenario_update_to_loc), .prefetch_enable(from_glob_prefetch_start_stop_dest_en[375]), .init_sram(init_sram));





	 
	 


   
endmodule
    

