

    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_0 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n121), .ZN(n1) );
  INVD6BWP30P140LVT U4 ( .I(n43), .ZN(n2) );
  INVD3BWP30P140LVT U5 ( .I(n42), .ZN(n196) );
  INVD4BWP30P140LVT U6 ( .I(n195), .ZN(n207) );
  OR2D2BWP30P140LVT U7 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .Z(n31) );
  ND2OPTPAD4BWP30P140LVT U8 ( .A1(n11), .A2(n14), .ZN(n195) );
  INVD3BWP30P140LVT U9 ( .I(n120), .ZN(n3) );
  INVD1BWP30P140LVT U10 ( .I(i_cmd[1]), .ZN(n25) );
  ND2D1BWP30P140LVT U11 ( .A1(n22), .A2(n6), .ZN(n7) );
  IOA21D1BWP30P140LVT U12 ( .A1(n210), .A2(i_data_bus[238]), .B(n188), .ZN(
        n189) );
  AOI22D1BWP30P140LVT U13 ( .A1(n208), .A2(i_data_bus[220]), .B1(n207), .B2(
        i_data_bus[188]), .ZN(n140) );
  INVD3BWP30P140LVT U14 ( .I(n30), .ZN(n213) );
  OR2D1BWP30P140LVT U15 ( .A1(n34), .A2(n29), .Z(n30) );
  AOI211D1BWP30P140LVT U16 ( .A1(n210), .A2(i_data_bus[224]), .B(n20), .C(n19), 
        .ZN(n40) );
  AOI21D1BWP30P140LVT U17 ( .A1(n142), .A2(i_data_bus[1]), .B(n58), .ZN(n61)
         );
  AOI21D1BWP30P140LVT U18 ( .A1(n142), .A2(i_data_bus[25]), .B(n119), .ZN(n124) );
  OR2D1BWP30P140LVT U19 ( .A1(n34), .A2(n26), .Z(n120) );
  OR2D1BWP30P140LVT U20 ( .A1(n34), .A2(n33), .Z(n121) );
  ND2D1BWP30P140LVT U21 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n4) );
  NR3D0P7BWP30P140LVT U22 ( .A1(n4), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n8) );
  NR2D1BWP30P140LVT U23 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n22) );
  INR2D1BWP30P140LVT U24 ( .A1(i_en), .B1(rst), .ZN(n5) );
  INR2D1BWP30P140LVT U25 ( .A1(n5), .B1(i_cmd[3]), .ZN(n6) );
  OR2D4BWP30P140LVT U26 ( .A1(n31), .A2(n7), .Z(n12) );
  INR2D4BWP30P140LVT U27 ( .A1(n8), .B1(n12), .ZN(n210) );
  INVD4BWP30P140LVT U28 ( .I(n12), .ZN(n11) );
  INVD1BWP30P140LVT U29 ( .I(i_cmd[6]), .ZN(n9) );
  INR4D0BWP30P140LVT U30 ( .A1(i_valid[6]), .B1(i_cmd[5]), .B2(i_cmd[7]), .B3(
        n9), .ZN(n10) );
  CKND2D4BWP30P140LVT U31 ( .A1(n11), .A2(n10), .ZN(n42) );
  INVD1BWP30P140LVT U32 ( .I(i_cmd[5]), .ZN(n13) );
  INR4D1BWP30P140LVT U33 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n13), .ZN(n14) );
  INVD4BWP30P140LVT U34 ( .I(n195), .ZN(n102) );
  AO22D1BWP30P140LVT U35 ( .A1(n196), .A2(i_data_bus[192]), .B1(n102), .B2(
        i_data_bus[160]), .Z(n20) );
  OR2D4BWP30P140LVT U36 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n27) );
  NR2D1BWP30P140LVT U37 ( .A1(n27), .A2(i_cmd[1]), .ZN(n17) );
  NR3D0P7BWP30P140LVT U38 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .A3(i_cmd[6]), .ZN(
        n21) );
  IND2D1BWP30P140LVT U39 ( .A1(rst), .B1(i_en), .ZN(n23) );
  INVD1BWP30P140LVT U40 ( .I(n23), .ZN(n15) );
  ND2OPTIBD1BWP30P140LVT U41 ( .A1(n21), .A2(n15), .ZN(n16) );
  INR2D2BWP30P140LVT U42 ( .A1(n17), .B1(n16), .ZN(n36) );
  INR2D1BWP30P140LVT U43 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n18) );
  ND3D2BWP30P140LVT U44 ( .A1(n36), .A2(i_cmd[0]), .A3(n18), .ZN(n41) );
  INR2D1BWP30P140LVT U45 ( .A1(i_data_bus[0]), .B1(n41), .ZN(n19) );
  IND3D1BWP30P140LVT U46 ( .A1(n23), .B1(n22), .B2(n21), .ZN(n34) );
  INVD1BWP30P140LVT U47 ( .I(i_cmd[3]), .ZN(n24) );
  ND4D1BWP30P140LVT U48 ( .A1(n25), .A2(n24), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n26) );
  INVD1BWP30P140LVT U49 ( .I(n27), .ZN(n28) );
  ND3D1BWP30P140LVT U50 ( .A1(n28), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n29)
         );
  AOI22D1BWP30P140LVT U51 ( .A1(n3), .A2(i_data_bus[64]), .B1(n213), .B2(
        i_data_bus[32]), .ZN(n39) );
  INVD0P7BWP30P140LVT U52 ( .I(n31), .ZN(n32) );
  ND3D1BWP30P140LVT U53 ( .A1(n32), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n33)
         );
  IND3D1BWP30P140LVT U54 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n35) );
  INR2D1BWP30P140LVT U55 ( .A1(n36), .B1(n35), .ZN(n37) );
  INVD2BWP30P140LVT U56 ( .I(n37), .ZN(n43) );
  AOI22D1BWP30P140LVT U57 ( .A1(n1), .A2(i_data_bus[96]), .B1(n2), .B2(
        i_data_bus[128]), .ZN(n38) );
  ND3D1BWP30P140LVT U58 ( .A1(n40), .A2(n39), .A3(n38), .ZN(N369) );
  INVD1BWP30P140LVT U59 ( .I(n41), .ZN(n142) );
  INVD3BWP30P140LVT U60 ( .I(n42), .ZN(n208) );
  NR4D0BWP30P140LVT U61 ( .A1(n142), .A2(n210), .A3(n208), .A4(n207), .ZN(n46)
         );
  NR2D1BWP30P140LVT U62 ( .A1(n3), .A2(n213), .ZN(n45) );
  NR2D1BWP30P140LVT U63 ( .A1(n1), .A2(n2), .ZN(n44) );
  ND3D1BWP30P140LVT U64 ( .A1(n46), .A2(n45), .A3(n44), .ZN(N402) );
  AOI22D1BWP30P140LVT U65 ( .A1(n196), .A2(i_data_bus[204]), .B1(n102), .B2(
        i_data_bus[172]), .ZN(n47) );
  IOA21D1BWP30P140LVT U66 ( .A1(n210), .A2(i_data_bus[236]), .B(n47), .ZN(n48)
         );
  AOI21D1BWP30P140LVT U67 ( .A1(n212), .A2(i_data_bus[12]), .B(n48), .ZN(n51)
         );
  AOI22D1BWP30P140LVT U68 ( .A1(n3), .A2(i_data_bus[76]), .B1(n213), .B2(
        i_data_bus[44]), .ZN(n50) );
  AOI22D1BWP30P140LVT U69 ( .A1(n1), .A2(i_data_bus[108]), .B1(n2), .B2(
        i_data_bus[140]), .ZN(n49) );
  ND3D1BWP30P140LVT U70 ( .A1(n51), .A2(n50), .A3(n49), .ZN(N381) );
  AOI22D1BWP30P140LVT U71 ( .A1(n196), .A2(i_data_bus[194]), .B1(n102), .B2(
        i_data_bus[162]), .ZN(n52) );
  IOA21D1BWP30P140LVT U72 ( .A1(n210), .A2(i_data_bus[226]), .B(n52), .ZN(n53)
         );
  AOI21D1BWP30P140LVT U73 ( .A1(n212), .A2(i_data_bus[2]), .B(n53), .ZN(n56)
         );
  AOI22D1BWP30P140LVT U74 ( .A1(n3), .A2(i_data_bus[66]), .B1(n213), .B2(
        i_data_bus[34]), .ZN(n55) );
  AOI22D1BWP30P140LVT U75 ( .A1(n1), .A2(i_data_bus[98]), .B1(n2), .B2(
        i_data_bus[130]), .ZN(n54) );
  ND3D1BWP30P140LVT U76 ( .A1(n56), .A2(n55), .A3(n54), .ZN(N371) );
  AOI22D1BWP30P140LVT U77 ( .A1(n196), .A2(i_data_bus[193]), .B1(n102), .B2(
        i_data_bus[161]), .ZN(n57) );
  IOA21D1BWP30P140LVT U78 ( .A1(n210), .A2(i_data_bus[225]), .B(n57), .ZN(n58)
         );
  AOI22D1BWP30P140LVT U79 ( .A1(n3), .A2(i_data_bus[65]), .B1(n213), .B2(
        i_data_bus[33]), .ZN(n60) );
  AOI22D1BWP30P140LVT U80 ( .A1(n1), .A2(i_data_bus[97]), .B1(n2), .B2(
        i_data_bus[129]), .ZN(n59) );
  ND3D1BWP30P140LVT U81 ( .A1(n61), .A2(n60), .A3(n59), .ZN(N370) );
  AOI22D1BWP30P140LVT U82 ( .A1(n196), .A2(i_data_bus[196]), .B1(n102), .B2(
        i_data_bus[164]), .ZN(n62) );
  IOA21D1BWP30P140LVT U83 ( .A1(n210), .A2(i_data_bus[228]), .B(n62), .ZN(n63)
         );
  AOI21D1BWP30P140LVT U84 ( .A1(n142), .A2(i_data_bus[4]), .B(n63), .ZN(n66)
         );
  AOI22D1BWP30P140LVT U85 ( .A1(n3), .A2(i_data_bus[68]), .B1(n213), .B2(
        i_data_bus[36]), .ZN(n65) );
  AOI22D1BWP30P140LVT U86 ( .A1(n1), .A2(i_data_bus[100]), .B1(n2), .B2(
        i_data_bus[132]), .ZN(n64) );
  ND3D1BWP30P140LVT U87 ( .A1(n66), .A2(n65), .A3(n64), .ZN(N373) );
  AOI22D1BWP30P140LVT U88 ( .A1(n196), .A2(i_data_bus[197]), .B1(n102), .B2(
        i_data_bus[165]), .ZN(n67) );
  IOA21D1BWP30P140LVT U89 ( .A1(n210), .A2(i_data_bus[229]), .B(n67), .ZN(n68)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n212), .A2(i_data_bus[5]), .B(n68), .ZN(n71)
         );
  AOI22D1BWP30P140LVT U91 ( .A1(n3), .A2(i_data_bus[69]), .B1(n213), .B2(
        i_data_bus[37]), .ZN(n70) );
  AOI22D1BWP30P140LVT U92 ( .A1(n1), .A2(i_data_bus[101]), .B1(n2), .B2(
        i_data_bus[133]), .ZN(n69) );
  ND3D1BWP30P140LVT U93 ( .A1(n71), .A2(n70), .A3(n69), .ZN(N374) );
  AOI22D1BWP30P140LVT U94 ( .A1(n196), .A2(i_data_bus[199]), .B1(n102), .B2(
        i_data_bus[167]), .ZN(n72) );
  IOA21D1BWP30P140LVT U95 ( .A1(n210), .A2(i_data_bus[231]), .B(n72), .ZN(n73)
         );
  AOI21D1BWP30P140LVT U96 ( .A1(n212), .A2(i_data_bus[7]), .B(n73), .ZN(n76)
         );
  AOI22D1BWP30P140LVT U97 ( .A1(n3), .A2(i_data_bus[71]), .B1(n213), .B2(
        i_data_bus[39]), .ZN(n75) );
  AOI22D1BWP30P140LVT U98 ( .A1(n1), .A2(i_data_bus[103]), .B1(n2), .B2(
        i_data_bus[135]), .ZN(n74) );
  ND3D1BWP30P140LVT U99 ( .A1(n76), .A2(n75), .A3(n74), .ZN(N376) );
  AOI22D1BWP30P140LVT U100 ( .A1(n196), .A2(i_data_bus[195]), .B1(n102), .B2(
        i_data_bus[163]), .ZN(n77) );
  IOA21D1BWP30P140LVT U101 ( .A1(n210), .A2(i_data_bus[227]), .B(n77), .ZN(n78) );
  AOI21D1BWP30P140LVT U102 ( .A1(n142), .A2(i_data_bus[3]), .B(n78), .ZN(n81)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n3), .A2(i_data_bus[67]), .B1(n213), .B2(
        i_data_bus[35]), .ZN(n80) );
  AOI22D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[99]), .B1(n2), .B2(
        i_data_bus[131]), .ZN(n79) );
  ND3D1BWP30P140LVT U105 ( .A1(n81), .A2(n80), .A3(n79), .ZN(N372) );
  AOI22D1BWP30P140LVT U106 ( .A1(n196), .A2(i_data_bus[201]), .B1(n102), .B2(
        i_data_bus[169]), .ZN(n82) );
  IOA21D1BWP30P140LVT U107 ( .A1(n210), .A2(i_data_bus[233]), .B(n82), .ZN(n83) );
  AOI21D1BWP30P140LVT U108 ( .A1(n212), .A2(i_data_bus[9]), .B(n83), .ZN(n86)
         );
  AOI22D1BWP30P140LVT U109 ( .A1(n3), .A2(i_data_bus[73]), .B1(n213), .B2(
        i_data_bus[41]), .ZN(n85) );
  AOI22D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[105]), .B1(n2), .B2(
        i_data_bus[137]), .ZN(n84) );
  ND3D1BWP30P140LVT U111 ( .A1(n86), .A2(n85), .A3(n84), .ZN(N378) );
  AOI22D1BWP30P140LVT U112 ( .A1(n196), .A2(i_data_bus[202]), .B1(n102), .B2(
        i_data_bus[170]), .ZN(n87) );
  IOA21D1BWP30P140LVT U113 ( .A1(n210), .A2(i_data_bus[234]), .B(n87), .ZN(n88) );
  AOI21D1BWP30P140LVT U114 ( .A1(n212), .A2(i_data_bus[10]), .B(n88), .ZN(n91)
         );
  AOI22D1BWP30P140LVT U115 ( .A1(n3), .A2(i_data_bus[74]), .B1(n213), .B2(
        i_data_bus[42]), .ZN(n90) );
  AOI22D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[106]), .B1(n2), .B2(
        i_data_bus[138]), .ZN(n89) );
  ND3D1BWP30P140LVT U117 ( .A1(n91), .A2(n90), .A3(n89), .ZN(N379) );
  AOI22D1BWP30P140LVT U118 ( .A1(n196), .A2(i_data_bus[203]), .B1(n102), .B2(
        i_data_bus[171]), .ZN(n92) );
  IOA21D1BWP30P140LVT U119 ( .A1(n210), .A2(i_data_bus[235]), .B(n92), .ZN(n93) );
  AOI21D1BWP30P140LVT U120 ( .A1(n142), .A2(i_data_bus[11]), .B(n93), .ZN(n96)
         );
  AOI22D1BWP30P140LVT U121 ( .A1(n3), .A2(i_data_bus[75]), .B1(n213), .B2(
        i_data_bus[43]), .ZN(n95) );
  AOI22D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[107]), .B1(n2), .B2(
        i_data_bus[139]), .ZN(n94) );
  ND3D1BWP30P140LVT U123 ( .A1(n96), .A2(n95), .A3(n94), .ZN(N380) );
  AOI22D1BWP30P140LVT U124 ( .A1(n196), .A2(i_data_bus[200]), .B1(n102), .B2(
        i_data_bus[168]), .ZN(n97) );
  IOA21D1BWP30P140LVT U125 ( .A1(n210), .A2(i_data_bus[232]), .B(n97), .ZN(n98) );
  AOI21D1BWP30P140LVT U126 ( .A1(n212), .A2(i_data_bus[8]), .B(n98), .ZN(n101)
         );
  AOI22D1BWP30P140LVT U127 ( .A1(n3), .A2(i_data_bus[72]), .B1(n213), .B2(
        i_data_bus[40]), .ZN(n100) );
  AOI22D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[104]), .B1(n2), .B2(
        i_data_bus[136]), .ZN(n99) );
  ND3D1BWP30P140LVT U129 ( .A1(n101), .A2(n100), .A3(n99), .ZN(N377) );
  AOI22D1BWP30P140LVT U130 ( .A1(n196), .A2(i_data_bus[198]), .B1(n102), .B2(
        i_data_bus[166]), .ZN(n103) );
  IOA21D1BWP30P140LVT U131 ( .A1(n210), .A2(i_data_bus[230]), .B(n103), .ZN(
        n104) );
  AOI21D1BWP30P140LVT U132 ( .A1(n212), .A2(i_data_bus[6]), .B(n104), .ZN(n107) );
  AOI22D1BWP30P140LVT U133 ( .A1(n3), .A2(i_data_bus[70]), .B1(n213), .B2(
        i_data_bus[38]), .ZN(n106) );
  AOI22D1BWP30P140LVT U134 ( .A1(n1), .A2(i_data_bus[102]), .B1(n2), .B2(
        i_data_bus[134]), .ZN(n105) );
  ND3D1BWP30P140LVT U135 ( .A1(n107), .A2(n106), .A3(n105), .ZN(N375) );
  AOI22D1BWP30P140LVT U136 ( .A1(n208), .A2(i_data_bus[218]), .B1(n207), .B2(
        i_data_bus[186]), .ZN(n108) );
  IOA21D1BWP30P140LVT U137 ( .A1(n210), .A2(i_data_bus[250]), .B(n108), .ZN(
        n109) );
  AOI21D1BWP30P140LVT U138 ( .A1(n142), .A2(i_data_bus[26]), .B(n109), .ZN(
        n112) );
  AOI22D1BWP30P140LVT U139 ( .A1(n3), .A2(i_data_bus[90]), .B1(n213), .B2(
        i_data_bus[58]), .ZN(n111) );
  AOI22D1BWP30P140LVT U140 ( .A1(n1), .A2(i_data_bus[122]), .B1(n2), .B2(
        i_data_bus[154]), .ZN(n110) );
  ND3D1BWP30P140LVT U141 ( .A1(n112), .A2(n111), .A3(n110), .ZN(N395) );
  AOI22D1BWP30P140LVT U142 ( .A1(n208), .A2(i_data_bus[219]), .B1(n207), .B2(
        i_data_bus[187]), .ZN(n113) );
  IOA21D1BWP30P140LVT U143 ( .A1(n210), .A2(i_data_bus[251]), .B(n113), .ZN(
        n114) );
  AOI21D1BWP30P140LVT U144 ( .A1(n142), .A2(i_data_bus[27]), .B(n114), .ZN(
        n117) );
  AOI22D1BWP30P140LVT U145 ( .A1(n3), .A2(i_data_bus[91]), .B1(n213), .B2(
        i_data_bus[59]), .ZN(n116) );
  AOI22D1BWP30P140LVT U146 ( .A1(n1), .A2(i_data_bus[123]), .B1(n2), .B2(
        i_data_bus[155]), .ZN(n115) );
  ND3D1BWP30P140LVT U147 ( .A1(n117), .A2(n116), .A3(n115), .ZN(N396) );
  AOI22D1BWP30P140LVT U148 ( .A1(n208), .A2(i_data_bus[217]), .B1(n207), .B2(
        i_data_bus[185]), .ZN(n118) );
  IOA21D1BWP30P140LVT U149 ( .A1(n210), .A2(i_data_bus[249]), .B(n118), .ZN(
        n119) );
  AOI22D1BWP30P140LVT U150 ( .A1(n3), .A2(i_data_bus[89]), .B1(n213), .B2(
        i_data_bus[57]), .ZN(n123) );
  AOI22D1BWP30P140LVT U151 ( .A1(n1), .A2(i_data_bus[121]), .B1(n2), .B2(
        i_data_bus[153]), .ZN(n122) );
  ND3D1BWP30P140LVT U152 ( .A1(n124), .A2(n123), .A3(n122), .ZN(N394) );
  AOI22D1BWP30P140LVT U153 ( .A1(n208), .A2(i_data_bus[221]), .B1(n207), .B2(
        i_data_bus[189]), .ZN(n125) );
  IOA21D1BWP30P140LVT U154 ( .A1(n210), .A2(i_data_bus[253]), .B(n125), .ZN(
        n126) );
  AOI21D1BWP30P140LVT U155 ( .A1(n142), .A2(i_data_bus[29]), .B(n126), .ZN(
        n129) );
  AOI22D1BWP30P140LVT U156 ( .A1(n3), .A2(i_data_bus[93]), .B1(n213), .B2(
        i_data_bus[61]), .ZN(n128) );
  AOI22D1BWP30P140LVT U157 ( .A1(n1), .A2(i_data_bus[125]), .B1(n2), .B2(
        i_data_bus[157]), .ZN(n127) );
  ND3D1BWP30P140LVT U158 ( .A1(n129), .A2(n128), .A3(n127), .ZN(N398) );
  AOI22D1BWP30P140LVT U159 ( .A1(n208), .A2(i_data_bus[222]), .B1(n207), .B2(
        i_data_bus[190]), .ZN(n130) );
  IOA21D1BWP30P140LVT U160 ( .A1(n210), .A2(i_data_bus[254]), .B(n130), .ZN(
        n131) );
  AOI21D1BWP30P140LVT U161 ( .A1(n142), .A2(i_data_bus[30]), .B(n131), .ZN(
        n134) );
  AOI22D1BWP30P140LVT U162 ( .A1(n3), .A2(i_data_bus[94]), .B1(n213), .B2(
        i_data_bus[62]), .ZN(n133) );
  AOI22D1BWP30P140LVT U163 ( .A1(n1), .A2(i_data_bus[126]), .B1(n2), .B2(
        i_data_bus[158]), .ZN(n132) );
  ND3D1BWP30P140LVT U164 ( .A1(n134), .A2(n133), .A3(n132), .ZN(N399) );
  AOI22D1BWP30P140LVT U165 ( .A1(n208), .A2(i_data_bus[223]), .B1(n207), .B2(
        i_data_bus[191]), .ZN(n135) );
  IOA21D1BWP30P140LVT U166 ( .A1(n210), .A2(i_data_bus[255]), .B(n135), .ZN(
        n136) );
  AOI21D1BWP30P140LVT U167 ( .A1(n142), .A2(i_data_bus[31]), .B(n136), .ZN(
        n139) );
  AOI22D1BWP30P140LVT U168 ( .A1(n3), .A2(i_data_bus[95]), .B1(n213), .B2(
        i_data_bus[63]), .ZN(n138) );
  AOI22D1BWP30P140LVT U169 ( .A1(n1), .A2(i_data_bus[127]), .B1(n2), .B2(
        i_data_bus[159]), .ZN(n137) );
  ND3D1BWP30P140LVT U170 ( .A1(n139), .A2(n138), .A3(n137), .ZN(N400) );
  IOA21D1BWP30P140LVT U171 ( .A1(n210), .A2(i_data_bus[252]), .B(n140), .ZN(
        n141) );
  AOI21D1BWP30P140LVT U172 ( .A1(n142), .A2(i_data_bus[28]), .B(n141), .ZN(
        n145) );
  AOI22D1BWP30P140LVT U173 ( .A1(n3), .A2(i_data_bus[92]), .B1(n213), .B2(
        i_data_bus[60]), .ZN(n144) );
  AOI22D1BWP30P140LVT U174 ( .A1(n1), .A2(i_data_bus[124]), .B1(n2), .B2(
        i_data_bus[156]), .ZN(n143) );
  ND3D1BWP30P140LVT U175 ( .A1(n145), .A2(n144), .A3(n143), .ZN(N397) );
  INVD2BWP30P140LVT U176 ( .I(n41), .ZN(n212) );
  AOI22D1BWP30P140LVT U177 ( .A1(n208), .A2(i_data_bus[208]), .B1(n207), .B2(
        i_data_bus[176]), .ZN(n146) );
  IOA21D1BWP30P140LVT U178 ( .A1(n210), .A2(i_data_bus[240]), .B(n146), .ZN(
        n147) );
  AOI21D1BWP30P140LVT U179 ( .A1(n212), .A2(i_data_bus[16]), .B(n147), .ZN(
        n150) );
  AOI22D1BWP30P140LVT U180 ( .A1(n3), .A2(i_data_bus[80]), .B1(n213), .B2(
        i_data_bus[48]), .ZN(n149) );
  AOI22D1BWP30P140LVT U181 ( .A1(n1), .A2(i_data_bus[112]), .B1(n2), .B2(
        i_data_bus[144]), .ZN(n148) );
  ND3D1BWP30P140LVT U182 ( .A1(n150), .A2(n149), .A3(n148), .ZN(N385) );
  AOI22D1BWP30P140LVT U183 ( .A1(n208), .A2(i_data_bus[211]), .B1(n207), .B2(
        i_data_bus[179]), .ZN(n151) );
  IOA21D1BWP30P140LVT U184 ( .A1(n210), .A2(i_data_bus[243]), .B(n151), .ZN(
        n152) );
  AOI21D1BWP30P140LVT U185 ( .A1(n212), .A2(i_data_bus[19]), .B(n152), .ZN(
        n155) );
  AOI22D1BWP30P140LVT U186 ( .A1(n3), .A2(i_data_bus[83]), .B1(n213), .B2(
        i_data_bus[51]), .ZN(n154) );
  AOI22D1BWP30P140LVT U187 ( .A1(n1), .A2(i_data_bus[115]), .B1(n2), .B2(
        i_data_bus[147]), .ZN(n153) );
  ND3D1BWP30P140LVT U188 ( .A1(n155), .A2(n154), .A3(n153), .ZN(N388) );
  AOI22D1BWP30P140LVT U189 ( .A1(n208), .A2(i_data_bus[210]), .B1(n207), .B2(
        i_data_bus[178]), .ZN(n156) );
  IOA21D1BWP30P140LVT U190 ( .A1(n210), .A2(i_data_bus[242]), .B(n156), .ZN(
        n157) );
  AOI21D1BWP30P140LVT U191 ( .A1(n212), .A2(i_data_bus[18]), .B(n157), .ZN(
        n160) );
  AOI22D1BWP30P140LVT U192 ( .A1(n3), .A2(i_data_bus[82]), .B1(n213), .B2(
        i_data_bus[50]), .ZN(n159) );
  AOI22D1BWP30P140LVT U193 ( .A1(n1), .A2(i_data_bus[114]), .B1(n2), .B2(
        i_data_bus[146]), .ZN(n158) );
  ND3D1BWP30P140LVT U194 ( .A1(n160), .A2(n159), .A3(n158), .ZN(N387) );
  AOI22D1BWP30P140LVT U195 ( .A1(n208), .A2(i_data_bus[215]), .B1(n207), .B2(
        i_data_bus[183]), .ZN(n161) );
  IOA21D1BWP30P140LVT U196 ( .A1(n210), .A2(i_data_bus[247]), .B(n161), .ZN(
        n162) );
  AOI21D1BWP30P140LVT U197 ( .A1(n212), .A2(i_data_bus[23]), .B(n162), .ZN(
        n165) );
  AOI22D1BWP30P140LVT U198 ( .A1(n3), .A2(i_data_bus[87]), .B1(n213), .B2(
        i_data_bus[55]), .ZN(n164) );
  AOI22D1BWP30P140LVT U199 ( .A1(n1), .A2(i_data_bus[119]), .B1(n2), .B2(
        i_data_bus[151]), .ZN(n163) );
  ND3D1BWP30P140LVT U200 ( .A1(n165), .A2(n164), .A3(n163), .ZN(N392) );
  AOI22D1BWP30P140LVT U201 ( .A1(n208), .A2(i_data_bus[216]), .B1(n207), .B2(
        i_data_bus[184]), .ZN(n166) );
  IOA21D1BWP30P140LVT U202 ( .A1(n210), .A2(i_data_bus[248]), .B(n166), .ZN(
        n167) );
  AOI21D1BWP30P140LVT U203 ( .A1(n212), .A2(i_data_bus[24]), .B(n167), .ZN(
        n170) );
  AOI22D1BWP30P140LVT U204 ( .A1(n3), .A2(i_data_bus[88]), .B1(n213), .B2(
        i_data_bus[56]), .ZN(n169) );
  AOI22D1BWP30P140LVT U205 ( .A1(n1), .A2(i_data_bus[120]), .B1(n2), .B2(
        i_data_bus[152]), .ZN(n168) );
  ND3D1BWP30P140LVT U206 ( .A1(n170), .A2(n169), .A3(n168), .ZN(N393) );
  AOI22D1BWP30P140LVT U207 ( .A1(n208), .A2(i_data_bus[209]), .B1(n207), .B2(
        i_data_bus[177]), .ZN(n171) );
  IOA21D1BWP30P140LVT U208 ( .A1(n210), .A2(i_data_bus[241]), .B(n171), .ZN(
        n172) );
  AOI21D1BWP30P140LVT U209 ( .A1(n212), .A2(i_data_bus[17]), .B(n172), .ZN(
        n175) );
  AOI22D1BWP30P140LVT U210 ( .A1(n3), .A2(i_data_bus[81]), .B1(n213), .B2(
        i_data_bus[49]), .ZN(n174) );
  AOI22D1BWP30P140LVT U211 ( .A1(n1), .A2(i_data_bus[113]), .B1(n2), .B2(
        i_data_bus[145]), .ZN(n173) );
  ND3D1BWP30P140LVT U212 ( .A1(n175), .A2(n174), .A3(n173), .ZN(N386) );
  AOI22D1BWP30P140LVT U213 ( .A1(n208), .A2(i_data_bus[212]), .B1(n207), .B2(
        i_data_bus[180]), .ZN(n176) );
  IOA21D1BWP30P140LVT U214 ( .A1(n210), .A2(i_data_bus[244]), .B(n176), .ZN(
        n177) );
  AOI21D1BWP30P140LVT U215 ( .A1(n212), .A2(i_data_bus[20]), .B(n177), .ZN(
        n180) );
  AOI22D1BWP30P140LVT U216 ( .A1(n3), .A2(i_data_bus[84]), .B1(n213), .B2(
        i_data_bus[52]), .ZN(n179) );
  AOI22D1BWP30P140LVT U217 ( .A1(n1), .A2(i_data_bus[116]), .B1(n2), .B2(
        i_data_bus[148]), .ZN(n178) );
  ND3D1BWP30P140LVT U218 ( .A1(n180), .A2(n179), .A3(n178), .ZN(N389) );
  AOI22D1BWP30P140LVT U219 ( .A1(n196), .A2(i_data_bus[207]), .B1(n207), .B2(
        i_data_bus[175]), .ZN(n181) );
  IOA21D1BWP30P140LVT U220 ( .A1(n210), .A2(i_data_bus[239]), .B(n181), .ZN(
        n182) );
  AOI21D1BWP30P140LVT U221 ( .A1(n212), .A2(i_data_bus[15]), .B(n182), .ZN(
        n185) );
  AOI22D1BWP30P140LVT U222 ( .A1(n3), .A2(i_data_bus[79]), .B1(n213), .B2(
        i_data_bus[47]), .ZN(n184) );
  AOI22D1BWP30P140LVT U223 ( .A1(n1), .A2(i_data_bus[111]), .B1(n2), .B2(
        i_data_bus[143]), .ZN(n183) );
  ND3D1BWP30P140LVT U224 ( .A1(n185), .A2(n184), .A3(n183), .ZN(N384) );
  INVD1BWP30P140LVT U225 ( .I(n212), .ZN(n187) );
  INVD1BWP30P140LVT U226 ( .I(i_data_bus[14]), .ZN(n186) );
  NR2D1BWP30P140LVT U227 ( .A1(n187), .A2(n186), .ZN(n190) );
  AOI22D1BWP30P140LVT U228 ( .A1(n196), .A2(i_data_bus[206]), .B1(n207), .B2(
        i_data_bus[174]), .ZN(n188) );
  NR2D1BWP30P140LVT U229 ( .A1(n190), .A2(n189), .ZN(n193) );
  AOI22D1BWP30P140LVT U230 ( .A1(n3), .A2(i_data_bus[78]), .B1(n213), .B2(
        i_data_bus[46]), .ZN(n192) );
  AOI22D1BWP30P140LVT U231 ( .A1(n1), .A2(i_data_bus[110]), .B1(n2), .B2(
        i_data_bus[142]), .ZN(n191) );
  ND3D1BWP30P140LVT U232 ( .A1(n193), .A2(n192), .A3(n191), .ZN(N383) );
  INVD1BWP30P140LVT U233 ( .I(i_data_bus[173]), .ZN(n194) );
  MAOI22D1BWP30P140LVT U234 ( .A1(n196), .A2(i_data_bus[205]), .B1(n195), .B2(
        n194), .ZN(n197) );
  IOA21D1BWP30P140LVT U235 ( .A1(n210), .A2(i_data_bus[237]), .B(n197), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U236 ( .A1(n212), .A2(i_data_bus[13]), .B(n198), .ZN(
        n201) );
  AOI22D1BWP30P140LVT U237 ( .A1(n3), .A2(i_data_bus[77]), .B1(n213), .B2(
        i_data_bus[45]), .ZN(n200) );
  AOI22D1BWP30P140LVT U238 ( .A1(n1), .A2(i_data_bus[109]), .B1(n2), .B2(
        i_data_bus[141]), .ZN(n199) );
  ND3D1BWP30P140LVT U239 ( .A1(n201), .A2(n200), .A3(n199), .ZN(N382) );
  AOI22D1BWP30P140LVT U240 ( .A1(n208), .A2(i_data_bus[213]), .B1(n207), .B2(
        i_data_bus[181]), .ZN(n202) );
  IOA21D1BWP30P140LVT U241 ( .A1(n210), .A2(i_data_bus[245]), .B(n202), .ZN(
        n203) );
  AOI21D1BWP30P140LVT U242 ( .A1(n212), .A2(i_data_bus[21]), .B(n203), .ZN(
        n206) );
  AOI22D1BWP30P140LVT U243 ( .A1(n3), .A2(i_data_bus[85]), .B1(n213), .B2(
        i_data_bus[53]), .ZN(n205) );
  AOI22D1BWP30P140LVT U244 ( .A1(n1), .A2(i_data_bus[117]), .B1(n2), .B2(
        i_data_bus[149]), .ZN(n204) );
  ND3D1BWP30P140LVT U245 ( .A1(n206), .A2(n205), .A3(n204), .ZN(N390) );
  AOI22D1BWP30P140LVT U246 ( .A1(n208), .A2(i_data_bus[214]), .B1(n207), .B2(
        i_data_bus[182]), .ZN(n209) );
  IOA21D1BWP30P140LVT U247 ( .A1(n210), .A2(i_data_bus[246]), .B(n209), .ZN(
        n211) );
  AOI21D1BWP30P140LVT U248 ( .A1(n212), .A2(i_data_bus[22]), .B(n211), .ZN(
        n216) );
  AOI22D1BWP30P140LVT U249 ( .A1(n3), .A2(i_data_bus[86]), .B1(n213), .B2(
        i_data_bus[54]), .ZN(n215) );
  AOI22D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[118]), .B1(n2), .B2(
        i_data_bus[150]), .ZN(n214) );
  ND3D1BWP30P140LVT U251 ( .A1(n216), .A2(n215), .A3(n214), .ZN(N391) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_1 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n141), .ZN(n3) );
  INVD2BWP30P140LVT U4 ( .I(n4), .ZN(n7) );
  INVD2BWP30P140LVT U5 ( .I(n26), .ZN(n66) );
  INR2D1BWP30P140LVT U6 ( .A1(n21), .B1(n25), .ZN(n22) );
  NR2OPTPAD1BWP30P140LVT U7 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .ZN(n8) );
  NR2OPTPAD1BWP30P140LVT U8 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n29) );
  AOI21D1BWP30P140LVT U9 ( .A1(n7), .A2(i_data_bus[14]), .B(n133), .ZN(n137)
         );
  INVD8BWP30P140LVT U10 ( .I(n66), .ZN(n1) );
  INVD4BWP30P140LVT U11 ( .I(n143), .ZN(n2) );
  ND2OPTPAD2BWP30P140LVT U12 ( .A1(n5), .A2(n8), .ZN(n25) );
  NR2OPTPAD1BWP30P140LVT U13 ( .A1(n25), .A2(n24), .ZN(n26) );
  INVD1BWP30P140LVT U14 ( .I(n33), .ZN(n61) );
  ND2OPTIBD1BWP30P140LVT U15 ( .A1(n44), .A2(n43), .ZN(n141) );
  ND3D1BWP30P140LVT U16 ( .A1(n23), .A2(i_cmd[5]), .A3(i_valid[5]), .ZN(n24)
         );
  NR2D1BWP30P140LVT U17 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .ZN(n23) );
  NR2D1BWP30P140LVT U18 ( .A1(n9), .A2(i_cmd[1]), .ZN(n44) );
  AN2D2BWP30P140LVT U19 ( .A1(n37), .A2(n35), .Z(n6) );
  NR2D1BWP30P140LVT U20 ( .A1(n9), .A2(n34), .ZN(n35) );
  ND2D1BWP30P140LVT U21 ( .A1(i_valid[1]), .A2(i_cmd[1]), .ZN(n34) );
  AOI21D1BWP30P140LVT U22 ( .A1(n7), .A2(i_data_bus[26]), .B(n28), .ZN(n47) );
  ND2OPTIBD1BWP30P140LVT U23 ( .A1(n44), .A2(n15), .ZN(n4) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n29), .A2(n18), .Z(n5) );
  INVD1BWP30P140LVT U25 ( .I(n38), .ZN(n143) );
  OR2D1BWP30P140LVT U26 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .Z(n9) );
  NR2OPTPAD2BWP30P140LVT U27 ( .A1(i_cmd[6]), .A2(i_cmd[5]), .ZN(n12) );
  INR2D1BWP30P140LVT U28 ( .A1(i_en), .B1(rst), .ZN(n10) );
  INR2D1BWP30P140LVT U29 ( .A1(n10), .B1(i_cmd[7]), .ZN(n11) );
  ND2OPTIBD2BWP30P140LVT U30 ( .A1(n12), .A2(n11), .ZN(n42) );
  INR2D1BWP30P140LVT U31 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n13) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n13), .A2(i_cmd[0]), .ZN(n14) );
  NR2D1BWP30P140LVT U33 ( .A1(n42), .A2(n14), .ZN(n15) );
  ND2D1BWP30P140LVT U34 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n16) );
  NR3D0P7BWP30P140LVT U35 ( .A1(n16), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n19)
         );
  INR2D1BWP30P140LVT U36 ( .A1(i_en), .B1(rst), .ZN(n17) );
  INR2D1BWP30P140LVT U37 ( .A1(n17), .B1(i_cmd[3]), .ZN(n18) );
  INR2D4BWP30P140LVT U38 ( .A1(n19), .B1(n25), .ZN(n216) );
  INVD1BWP30P140LVT U39 ( .I(i_cmd[6]), .ZN(n20) );
  INR4D0BWP30P140LVT U40 ( .A1(i_valid[6]), .B1(i_cmd[5]), .B2(i_cmd[7]), .B3(
        n20), .ZN(n21) );
  INVD2BWP30P140LVT U41 ( .I(n22), .ZN(n48) );
  INVD3BWP30P140LVT U42 ( .I(n48), .ZN(n152) );
  AOI22D1BWP30P140LVT U43 ( .A1(n152), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n27) );
  IOA21D1BWP30P140LVT U44 ( .A1(n216), .A2(i_data_bus[250]), .B(n27), .ZN(n28)
         );
  INR2D2BWP30P140LVT U45 ( .A1(n29), .B1(n42), .ZN(n37) );
  INVD1BWP30P140LVT U46 ( .I(i_cmd[1]), .ZN(n31) );
  INVD1BWP30P140LVT U47 ( .I(i_cmd[3]), .ZN(n30) );
  ND4D1BWP30P140LVT U48 ( .A1(n31), .A2(n30), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n32) );
  INR2D1BWP30P140LVT U49 ( .A1(n37), .B1(n32), .ZN(n33) );
  INVD1BWP30P140LVT U50 ( .I(n61), .ZN(n155) );
  AOI22D1BWP30P140LVT U51 ( .A1(n155), .A2(i_data_bus[90]), .B1(n6), .B2(
        i_data_bus[58]), .ZN(n46) );
  ND3D1BWP30P140LVT U52 ( .A1(n8), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n36) );
  INR2D1BWP30P140LVT U53 ( .A1(n37), .B1(n36), .ZN(n38) );
  INVD1BWP30P140LVT U54 ( .I(i_cmd[0]), .ZN(n39) );
  ND2OPTIBD1BWP30P140LVT U55 ( .A1(n39), .A2(i_cmd[4]), .ZN(n41) );
  INVD1BWP30P140LVT U56 ( .I(i_valid[4]), .ZN(n40) );
  NR3D0P7BWP30P140LVT U57 ( .A1(n42), .A2(n41), .A3(n40), .ZN(n43) );
  AOI22D1BWP30P140LVT U58 ( .A1(n2), .A2(i_data_bus[122]), .B1(n3), .B2(
        i_data_bus[154]), .ZN(n45) );
  ND3D1BWP30P140LVT U59 ( .A1(n47), .A2(n46), .A3(n45), .ZN(N395) );
  INVD1BWP30P140LVT U60 ( .I(n216), .ZN(n52) );
  INVD1BWP30P140LVT U61 ( .I(i_data_bus[224]), .ZN(n51) );
  INVD3BWP30P140LVT U62 ( .I(n48), .ZN(n214) );
  AOI22D1BWP30P140LVT U63 ( .A1(n214), .A2(i_data_bus[192]), .B1(n1), .B2(
        i_data_bus[160]), .ZN(n50) );
  ND2D1BWP30P140LVT U64 ( .A1(i_data_bus[0]), .A2(n7), .ZN(n49) );
  OA211D1BWP30P140LVT U65 ( .A1(n52), .A2(n51), .B(n50), .C(n49), .Z(n55) );
  INVD2BWP30P140LVT U66 ( .I(n61), .ZN(n218) );
  AOI22D1BWP30P140LVT U67 ( .A1(n218), .A2(i_data_bus[64]), .B1(n6), .B2(
        i_data_bus[32]), .ZN(n54) );
  AOI22D1BWP30P140LVT U68 ( .A1(n2), .A2(i_data_bus[96]), .B1(n3), .B2(
        i_data_bus[128]), .ZN(n53) );
  ND3D1BWP30P140LVT U69 ( .A1(n55), .A2(n54), .A3(n53), .ZN(N369) );
  NR4D0BWP30P140LVT U70 ( .A1(n7), .A2(n216), .A3(n152), .A4(n1), .ZN(n58) );
  NR2D1BWP30P140LVT U71 ( .A1(n155), .A2(n6), .ZN(n57) );
  NR2D1BWP30P140LVT U72 ( .A1(n2), .A2(n3), .ZN(n56) );
  ND3D1BWP30P140LVT U73 ( .A1(n58), .A2(n57), .A3(n56), .ZN(N402) );
  AOI22D1BWP30P140LVT U74 ( .A1(n152), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n59) );
  IOA21D1BWP30P140LVT U75 ( .A1(n216), .A2(i_data_bus[247]), .B(n59), .ZN(n60)
         );
  AOI21D1BWP30P140LVT U76 ( .A1(n7), .A2(i_data_bus[23]), .B(n60), .ZN(n64) );
  INVD2BWP30P140LVT U77 ( .I(n61), .ZN(n134) );
  AOI22D1BWP30P140LVT U78 ( .A1(n134), .A2(i_data_bus[87]), .B1(n6), .B2(
        i_data_bus[55]), .ZN(n63) );
  AOI22D1BWP30P140LVT U79 ( .A1(n2), .A2(i_data_bus[119]), .B1(n3), .B2(
        i_data_bus[151]), .ZN(n62) );
  ND3D1BWP30P140LVT U80 ( .A1(n64), .A2(n63), .A3(n62), .ZN(N392) );
  INVD1BWP30P140LVT U81 ( .I(i_data_bus[173]), .ZN(n65) );
  MAOI22D1BWP30P140LVT U82 ( .A1(n214), .A2(i_data_bus[205]), .B1(n66), .B2(
        n65), .ZN(n67) );
  IOA21D1BWP30P140LVT U83 ( .A1(n216), .A2(i_data_bus[237]), .B(n67), .ZN(n68)
         );
  AOI21D1BWP30P140LVT U84 ( .A1(n7), .A2(i_data_bus[13]), .B(n68), .ZN(n71) );
  AOI22D1BWP30P140LVT U85 ( .A1(n134), .A2(i_data_bus[77]), .B1(n6), .B2(
        i_data_bus[45]), .ZN(n70) );
  AOI22D1BWP30P140LVT U86 ( .A1(n2), .A2(i_data_bus[109]), .B1(n3), .B2(
        i_data_bus[141]), .ZN(n69) );
  ND3D1BWP30P140LVT U87 ( .A1(n71), .A2(n70), .A3(n69), .ZN(N382) );
  AOI22D1BWP30P140LVT U88 ( .A1(n152), .A2(i_data_bus[221]), .B1(n1), .B2(
        i_data_bus[189]), .ZN(n72) );
  IOA21D1BWP30P140LVT U89 ( .A1(n216), .A2(i_data_bus[253]), .B(n72), .ZN(n73)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n7), .A2(i_data_bus[29]), .B(n73), .ZN(n76) );
  AOI22D1BWP30P140LVT U91 ( .A1(n155), .A2(i_data_bus[93]), .B1(n6), .B2(
        i_data_bus[61]), .ZN(n75) );
  AOI22D1BWP30P140LVT U92 ( .A1(n2), .A2(i_data_bus[125]), .B1(n3), .B2(
        i_data_bus[157]), .ZN(n74) );
  ND3D1BWP30P140LVT U93 ( .A1(n76), .A2(n75), .A3(n74), .ZN(N398) );
  AOI22D1BWP30P140LVT U94 ( .A1(n152), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n77) );
  IOA21D1BWP30P140LVT U95 ( .A1(n216), .A2(i_data_bus[242]), .B(n77), .ZN(n78)
         );
  AOI21D1BWP30P140LVT U96 ( .A1(n7), .A2(i_data_bus[18]), .B(n78), .ZN(n81) );
  AOI22D1BWP30P140LVT U97 ( .A1(n134), .A2(i_data_bus[82]), .B1(n6), .B2(
        i_data_bus[50]), .ZN(n80) );
  AOI22D1BWP30P140LVT U98 ( .A1(n2), .A2(i_data_bus[114]), .B1(n3), .B2(
        i_data_bus[146]), .ZN(n79) );
  ND3D1BWP30P140LVT U99 ( .A1(n81), .A2(n80), .A3(n79), .ZN(N387) );
  AOI22D1BWP30P140LVT U100 ( .A1(n152), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n82) );
  IOA21D1BWP30P140LVT U101 ( .A1(n216), .A2(i_data_bus[251]), .B(n82), .ZN(n83) );
  AOI21D1BWP30P140LVT U102 ( .A1(n7), .A2(i_data_bus[27]), .B(n83), .ZN(n86)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n155), .A2(i_data_bus[91]), .B1(n6), .B2(
        i_data_bus[59]), .ZN(n85) );
  AOI22D1BWP30P140LVT U104 ( .A1(n2), .A2(i_data_bus[123]), .B1(n3), .B2(
        i_data_bus[155]), .ZN(n84) );
  ND3D1BWP30P140LVT U105 ( .A1(n86), .A2(n85), .A3(n84), .ZN(N396) );
  AOI22D1BWP30P140LVT U106 ( .A1(n152), .A2(i_data_bus[208]), .B1(n1), .B2(
        i_data_bus[176]), .ZN(n87) );
  IOA21D1BWP30P140LVT U107 ( .A1(n216), .A2(i_data_bus[240]), .B(n87), .ZN(n88) );
  AOI21D1BWP30P140LVT U108 ( .A1(n7), .A2(i_data_bus[16]), .B(n88), .ZN(n91)
         );
  AOI22D1BWP30P140LVT U109 ( .A1(n134), .A2(i_data_bus[80]), .B1(n6), .B2(
        i_data_bus[48]), .ZN(n90) );
  AOI22D1BWP30P140LVT U110 ( .A1(n2), .A2(i_data_bus[112]), .B1(n3), .B2(
        i_data_bus[144]), .ZN(n89) );
  ND3D1BWP30P140LVT U111 ( .A1(n91), .A2(n90), .A3(n89), .ZN(N385) );
  AOI22D1BWP30P140LVT U112 ( .A1(n152), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n92) );
  IOA21D1BWP30P140LVT U113 ( .A1(n216), .A2(i_data_bus[249]), .B(n92), .ZN(n93) );
  AOI21D1BWP30P140LVT U114 ( .A1(n7), .A2(i_data_bus[25]), .B(n93), .ZN(n96)
         );
  AOI22D1BWP30P140LVT U115 ( .A1(n134), .A2(i_data_bus[89]), .B1(n6), .B2(
        i_data_bus[57]), .ZN(n95) );
  AOI22D1BWP30P140LVT U116 ( .A1(n2), .A2(i_data_bus[121]), .B1(n3), .B2(
        i_data_bus[153]), .ZN(n94) );
  ND3D1BWP30P140LVT U117 ( .A1(n96), .A2(n95), .A3(n94), .ZN(N394) );
  AOI22D1BWP30P140LVT U118 ( .A1(n152), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n97) );
  IOA21D1BWP30P140LVT U119 ( .A1(n216), .A2(i_data_bus[248]), .B(n97), .ZN(n98) );
  AOI21D1BWP30P140LVT U120 ( .A1(n7), .A2(i_data_bus[24]), .B(n98), .ZN(n101)
         );
  AOI22D1BWP30P140LVT U121 ( .A1(n134), .A2(i_data_bus[88]), .B1(n6), .B2(
        i_data_bus[56]), .ZN(n100) );
  AOI22D1BWP30P140LVT U122 ( .A1(n2), .A2(i_data_bus[120]), .B1(n3), .B2(
        i_data_bus[152]), .ZN(n99) );
  ND3D1BWP30P140LVT U123 ( .A1(n101), .A2(n100), .A3(n99), .ZN(N393) );
  AOI22D1BWP30P140LVT U124 ( .A1(n152), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n102) );
  IOA21D1BWP30P140LVT U125 ( .A1(n216), .A2(i_data_bus[243]), .B(n102), .ZN(
        n103) );
  AOI21D1BWP30P140LVT U126 ( .A1(n7), .A2(i_data_bus[19]), .B(n103), .ZN(n106)
         );
  AOI22D1BWP30P140LVT U127 ( .A1(n134), .A2(i_data_bus[83]), .B1(n6), .B2(
        i_data_bus[51]), .ZN(n105) );
  AOI22D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[115]), .B1(n3), .B2(
        i_data_bus[147]), .ZN(n104) );
  ND3D1BWP30P140LVT U129 ( .A1(n106), .A2(n105), .A3(n104), .ZN(N388) );
  AOI22D1BWP30P140LVT U130 ( .A1(n152), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n107) );
  IOA21D1BWP30P140LVT U131 ( .A1(n216), .A2(i_data_bus[246]), .B(n107), .ZN(
        n108) );
  AOI21D1BWP30P140LVT U132 ( .A1(n7), .A2(i_data_bus[22]), .B(n108), .ZN(n111)
         );
  AOI22D1BWP30P140LVT U133 ( .A1(n134), .A2(i_data_bus[86]), .B1(n6), .B2(
        i_data_bus[54]), .ZN(n110) );
  AOI22D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[118]), .B1(n3), .B2(
        i_data_bus[150]), .ZN(n109) );
  ND3D1BWP30P140LVT U135 ( .A1(n111), .A2(n110), .A3(n109), .ZN(N391) );
  AOI22D1BWP30P140LVT U136 ( .A1(n152), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n112) );
  IOA21D1BWP30P140LVT U137 ( .A1(n216), .A2(i_data_bus[245]), .B(n112), .ZN(
        n113) );
  AOI21D1BWP30P140LVT U138 ( .A1(n7), .A2(i_data_bus[21]), .B(n113), .ZN(n116)
         );
  AOI22D1BWP30P140LVT U139 ( .A1(n134), .A2(i_data_bus[85]), .B1(n6), .B2(
        i_data_bus[53]), .ZN(n115) );
  AOI22D1BWP30P140LVT U140 ( .A1(n2), .A2(i_data_bus[117]), .B1(n3), .B2(
        i_data_bus[149]), .ZN(n114) );
  ND3D1BWP30P140LVT U141 ( .A1(n116), .A2(n115), .A3(n114), .ZN(N390) );
  AOI22D1BWP30P140LVT U142 ( .A1(n214), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n117) );
  IOA21D1BWP30P140LVT U143 ( .A1(n216), .A2(i_data_bus[239]), .B(n117), .ZN(
        n118) );
  AOI21D1BWP30P140LVT U144 ( .A1(n7), .A2(i_data_bus[15]), .B(n118), .ZN(n121)
         );
  AOI22D1BWP30P140LVT U145 ( .A1(n134), .A2(i_data_bus[79]), .B1(n6), .B2(
        i_data_bus[47]), .ZN(n120) );
  AOI22D1BWP30P140LVT U146 ( .A1(n2), .A2(i_data_bus[111]), .B1(n3), .B2(
        i_data_bus[143]), .ZN(n119) );
  ND3D1BWP30P140LVT U147 ( .A1(n121), .A2(n120), .A3(n119), .ZN(N384) );
  AOI22D1BWP30P140LVT U148 ( .A1(n152), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n122) );
  IOA21D1BWP30P140LVT U149 ( .A1(n216), .A2(i_data_bus[244]), .B(n122), .ZN(
        n123) );
  AOI21D1BWP30P140LVT U150 ( .A1(n7), .A2(i_data_bus[20]), .B(n123), .ZN(n126)
         );
  AOI22D1BWP30P140LVT U151 ( .A1(n134), .A2(i_data_bus[84]), .B1(n6), .B2(
        i_data_bus[52]), .ZN(n125) );
  AOI22D1BWP30P140LVT U152 ( .A1(n2), .A2(i_data_bus[116]), .B1(n3), .B2(
        i_data_bus[148]), .ZN(n124) );
  ND3D1BWP30P140LVT U153 ( .A1(n126), .A2(n125), .A3(n124), .ZN(N389) );
  AOI22D1BWP30P140LVT U154 ( .A1(n152), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n127) );
  IOA21D1BWP30P140LVT U155 ( .A1(n216), .A2(i_data_bus[241]), .B(n127), .ZN(
        n128) );
  AOI21D1BWP30P140LVT U156 ( .A1(n7), .A2(i_data_bus[17]), .B(n128), .ZN(n131)
         );
  AOI22D1BWP30P140LVT U157 ( .A1(n134), .A2(i_data_bus[81]), .B1(n6), .B2(
        i_data_bus[49]), .ZN(n130) );
  AOI22D1BWP30P140LVT U158 ( .A1(n2), .A2(i_data_bus[113]), .B1(n3), .B2(
        i_data_bus[145]), .ZN(n129) );
  ND3D1BWP30P140LVT U159 ( .A1(n131), .A2(n130), .A3(n129), .ZN(N386) );
  AOI22D1BWP30P140LVT U160 ( .A1(n214), .A2(i_data_bus[206]), .B1(n1), .B2(
        i_data_bus[174]), .ZN(n132) );
  IOA21D1BWP30P140LVT U161 ( .A1(n216), .A2(i_data_bus[238]), .B(n132), .ZN(
        n133) );
  AOI22D1BWP30P140LVT U162 ( .A1(n134), .A2(i_data_bus[78]), .B1(n6), .B2(
        i_data_bus[46]), .ZN(n136) );
  AOI22D1BWP30P140LVT U163 ( .A1(n2), .A2(i_data_bus[110]), .B1(n3), .B2(
        i_data_bus[142]), .ZN(n135) );
  ND3D1BWP30P140LVT U164 ( .A1(n137), .A2(n136), .A3(n135), .ZN(N383) );
  AOI22D1BWP30P140LVT U165 ( .A1(n152), .A2(i_data_bus[223]), .B1(n1), .B2(
        i_data_bus[191]), .ZN(n138) );
  IOA21D1BWP30P140LVT U166 ( .A1(n216), .A2(i_data_bus[255]), .B(n138), .ZN(
        n139) );
  AOI21D1BWP30P140LVT U167 ( .A1(n7), .A2(i_data_bus[31]), .B(n139), .ZN(n146)
         );
  AOI22D1BWP30P140LVT U168 ( .A1(n155), .A2(i_data_bus[95]), .B1(n6), .B2(
        i_data_bus[63]), .ZN(n145) );
  INVD1BWP30P140LVT U169 ( .I(i_data_bus[127]), .ZN(n142) );
  INVD1BWP30P140LVT U170 ( .I(i_data_bus[159]), .ZN(n140) );
  OA22D1BWP30P140LVT U171 ( .A1(n143), .A2(n142), .B1(n141), .B2(n140), .Z(
        n144) );
  ND3D1BWP30P140LVT U172 ( .A1(n146), .A2(n145), .A3(n144), .ZN(N400) );
  AOI22D1BWP30P140LVT U173 ( .A1(n152), .A2(i_data_bus[222]), .B1(n1), .B2(
        i_data_bus[190]), .ZN(n147) );
  IOA21D1BWP30P140LVT U174 ( .A1(n216), .A2(i_data_bus[254]), .B(n147), .ZN(
        n148) );
  AOI21D1BWP30P140LVT U175 ( .A1(n7), .A2(i_data_bus[30]), .B(n148), .ZN(n151)
         );
  AOI22D1BWP30P140LVT U176 ( .A1(n155), .A2(i_data_bus[94]), .B1(n6), .B2(
        i_data_bus[62]), .ZN(n150) );
  AOI22D1BWP30P140LVT U177 ( .A1(n2), .A2(i_data_bus[126]), .B1(n3), .B2(
        i_data_bus[158]), .ZN(n149) );
  ND3D1BWP30P140LVT U178 ( .A1(n151), .A2(n150), .A3(n149), .ZN(N399) );
  AOI22D1BWP30P140LVT U179 ( .A1(n152), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n153) );
  IOA21D1BWP30P140LVT U180 ( .A1(n216), .A2(i_data_bus[252]), .B(n153), .ZN(
        n154) );
  AOI21D1BWP30P140LVT U181 ( .A1(n7), .A2(i_data_bus[28]), .B(n154), .ZN(n158)
         );
  AOI22D1BWP30P140LVT U182 ( .A1(n155), .A2(i_data_bus[92]), .B1(n6), .B2(
        i_data_bus[60]), .ZN(n157) );
  AOI22D1BWP30P140LVT U183 ( .A1(n2), .A2(i_data_bus[124]), .B1(n3), .B2(
        i_data_bus[156]), .ZN(n156) );
  ND3D1BWP30P140LVT U184 ( .A1(n158), .A2(n157), .A3(n156), .ZN(N397) );
  AOI22D1BWP30P140LVT U185 ( .A1(n214), .A2(i_data_bus[193]), .B1(n1), .B2(
        i_data_bus[161]), .ZN(n159) );
  IOA21D1BWP30P140LVT U186 ( .A1(n216), .A2(i_data_bus[225]), .B(n159), .ZN(
        n160) );
  AOI21D1BWP30P140LVT U187 ( .A1(n7), .A2(i_data_bus[1]), .B(n160), .ZN(n163)
         );
  AOI22D1BWP30P140LVT U188 ( .A1(n218), .A2(i_data_bus[65]), .B1(n6), .B2(
        i_data_bus[33]), .ZN(n162) );
  AOI22D1BWP30P140LVT U189 ( .A1(n2), .A2(i_data_bus[97]), .B1(n3), .B2(
        i_data_bus[129]), .ZN(n161) );
  ND3D1BWP30P140LVT U190 ( .A1(n163), .A2(n162), .A3(n161), .ZN(N370) );
  AOI22D1BWP30P140LVT U191 ( .A1(n214), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n164) );
  IOA21D1BWP30P140LVT U192 ( .A1(n216), .A2(i_data_bus[228]), .B(n164), .ZN(
        n165) );
  AOI21D1BWP30P140LVT U193 ( .A1(n7), .A2(i_data_bus[4]), .B(n165), .ZN(n168)
         );
  AOI22D1BWP30P140LVT U194 ( .A1(n218), .A2(i_data_bus[68]), .B1(n6), .B2(
        i_data_bus[36]), .ZN(n167) );
  AOI22D1BWP30P140LVT U195 ( .A1(n2), .A2(i_data_bus[100]), .B1(n3), .B2(
        i_data_bus[132]), .ZN(n166) );
  ND3D1BWP30P140LVT U196 ( .A1(n168), .A2(n167), .A3(n166), .ZN(N373) );
  AOI22D1BWP30P140LVT U197 ( .A1(n214), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n169) );
  IOA21D1BWP30P140LVT U198 ( .A1(n216), .A2(i_data_bus[235]), .B(n169), .ZN(
        n170) );
  AOI21D1BWP30P140LVT U199 ( .A1(n7), .A2(i_data_bus[11]), .B(n170), .ZN(n173)
         );
  AOI22D1BWP30P140LVT U200 ( .A1(n218), .A2(i_data_bus[75]), .B1(n6), .B2(
        i_data_bus[43]), .ZN(n172) );
  AOI22D1BWP30P140LVT U201 ( .A1(n2), .A2(i_data_bus[107]), .B1(n3), .B2(
        i_data_bus[139]), .ZN(n171) );
  ND3D1BWP30P140LVT U202 ( .A1(n173), .A2(n172), .A3(n171), .ZN(N380) );
  AOI22D1BWP30P140LVT U203 ( .A1(n214), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n174) );
  IOA21D1BWP30P140LVT U204 ( .A1(n216), .A2(i_data_bus[233]), .B(n174), .ZN(
        n175) );
  AOI21D1BWP30P140LVT U205 ( .A1(n7), .A2(i_data_bus[9]), .B(n175), .ZN(n178)
         );
  AOI22D1BWP30P140LVT U206 ( .A1(n218), .A2(i_data_bus[73]), .B1(n6), .B2(
        i_data_bus[41]), .ZN(n177) );
  AOI22D1BWP30P140LVT U207 ( .A1(n2), .A2(i_data_bus[105]), .B1(n3), .B2(
        i_data_bus[137]), .ZN(n176) );
  ND3D1BWP30P140LVT U208 ( .A1(n178), .A2(n177), .A3(n176), .ZN(N378) );
  AOI22D1BWP30P140LVT U209 ( .A1(n214), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n179) );
  IOA21D1BWP30P140LVT U210 ( .A1(n216), .A2(i_data_bus[236]), .B(n179), .ZN(
        n180) );
  AOI21D1BWP30P140LVT U211 ( .A1(n7), .A2(i_data_bus[12]), .B(n180), .ZN(n183)
         );
  AOI22D1BWP30P140LVT U212 ( .A1(n218), .A2(i_data_bus[76]), .B1(n6), .B2(
        i_data_bus[44]), .ZN(n182) );
  AOI22D1BWP30P140LVT U213 ( .A1(n2), .A2(i_data_bus[108]), .B1(n3), .B2(
        i_data_bus[140]), .ZN(n181) );
  ND3D1BWP30P140LVT U214 ( .A1(n183), .A2(n182), .A3(n181), .ZN(N381) );
  AOI22D1BWP30P140LVT U215 ( .A1(n214), .A2(i_data_bus[199]), .B1(n1), .B2(
        i_data_bus[167]), .ZN(n184) );
  IOA21D1BWP30P140LVT U216 ( .A1(n216), .A2(i_data_bus[231]), .B(n184), .ZN(
        n185) );
  AOI21D1BWP30P140LVT U217 ( .A1(n7), .A2(i_data_bus[7]), .B(n185), .ZN(n188)
         );
  AOI22D1BWP30P140LVT U218 ( .A1(n218), .A2(i_data_bus[71]), .B1(n6), .B2(
        i_data_bus[39]), .ZN(n187) );
  AOI22D1BWP30P140LVT U219 ( .A1(n2), .A2(i_data_bus[103]), .B1(n3), .B2(
        i_data_bus[135]), .ZN(n186) );
  ND3D1BWP30P140LVT U220 ( .A1(n188), .A2(n187), .A3(n186), .ZN(N376) );
  AOI22D1BWP30P140LVT U221 ( .A1(n214), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n189) );
  IOA21D1BWP30P140LVT U222 ( .A1(n216), .A2(i_data_bus[234]), .B(n189), .ZN(
        n190) );
  AOI21D1BWP30P140LVT U223 ( .A1(n7), .A2(i_data_bus[10]), .B(n190), .ZN(n193)
         );
  AOI22D1BWP30P140LVT U224 ( .A1(n218), .A2(i_data_bus[74]), .B1(n6), .B2(
        i_data_bus[42]), .ZN(n192) );
  AOI22D1BWP30P140LVT U225 ( .A1(n2), .A2(i_data_bus[106]), .B1(n3), .B2(
        i_data_bus[138]), .ZN(n191) );
  ND3D1BWP30P140LVT U226 ( .A1(n193), .A2(n192), .A3(n191), .ZN(N379) );
  AOI22D1BWP30P140LVT U227 ( .A1(n214), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n194) );
  IOA21D1BWP30P140LVT U228 ( .A1(n216), .A2(i_data_bus[230]), .B(n194), .ZN(
        n195) );
  AOI21D1BWP30P140LVT U229 ( .A1(n7), .A2(i_data_bus[6]), .B(n195), .ZN(n198)
         );
  AOI22D1BWP30P140LVT U230 ( .A1(n218), .A2(i_data_bus[70]), .B1(n6), .B2(
        i_data_bus[38]), .ZN(n197) );
  AOI22D1BWP30P140LVT U231 ( .A1(n2), .A2(i_data_bus[102]), .B1(n3), .B2(
        i_data_bus[134]), .ZN(n196) );
  ND3D1BWP30P140LVT U232 ( .A1(n198), .A2(n197), .A3(n196), .ZN(N375) );
  AOI22D1BWP30P140LVT U233 ( .A1(n214), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n199) );
  IOA21D1BWP30P140LVT U234 ( .A1(n216), .A2(i_data_bus[229]), .B(n199), .ZN(
        n200) );
  AOI21D1BWP30P140LVT U235 ( .A1(n7), .A2(i_data_bus[5]), .B(n200), .ZN(n203)
         );
  AOI22D1BWP30P140LVT U236 ( .A1(n218), .A2(i_data_bus[69]), .B1(n6), .B2(
        i_data_bus[37]), .ZN(n202) );
  AOI22D1BWP30P140LVT U237 ( .A1(n2), .A2(i_data_bus[101]), .B1(n3), .B2(
        i_data_bus[133]), .ZN(n201) );
  ND3D1BWP30P140LVT U238 ( .A1(n203), .A2(n202), .A3(n201), .ZN(N374) );
  AOI22D1BWP30P140LVT U239 ( .A1(n214), .A2(i_data_bus[195]), .B1(n1), .B2(
        i_data_bus[163]), .ZN(n204) );
  IOA21D1BWP30P140LVT U240 ( .A1(n216), .A2(i_data_bus[227]), .B(n204), .ZN(
        n205) );
  AOI21D1BWP30P140LVT U241 ( .A1(n7), .A2(i_data_bus[3]), .B(n205), .ZN(n208)
         );
  AOI22D1BWP30P140LVT U242 ( .A1(n218), .A2(i_data_bus[67]), .B1(n6), .B2(
        i_data_bus[35]), .ZN(n207) );
  AOI22D1BWP30P140LVT U243 ( .A1(n2), .A2(i_data_bus[99]), .B1(n3), .B2(
        i_data_bus[131]), .ZN(n206) );
  ND3D1BWP30P140LVT U244 ( .A1(n208), .A2(n207), .A3(n206), .ZN(N372) );
  AOI22D1BWP30P140LVT U245 ( .A1(n214), .A2(i_data_bus[194]), .B1(n1), .B2(
        i_data_bus[162]), .ZN(n209) );
  IOA21D1BWP30P140LVT U246 ( .A1(n216), .A2(i_data_bus[226]), .B(n209), .ZN(
        n210) );
  AOI21D1BWP30P140LVT U247 ( .A1(n7), .A2(i_data_bus[2]), .B(n210), .ZN(n213)
         );
  AOI22D1BWP30P140LVT U248 ( .A1(n218), .A2(i_data_bus[66]), .B1(n6), .B2(
        i_data_bus[34]), .ZN(n212) );
  AOI22D1BWP30P140LVT U249 ( .A1(n2), .A2(i_data_bus[98]), .B1(n3), .B2(
        i_data_bus[130]), .ZN(n211) );
  ND3D1BWP30P140LVT U250 ( .A1(n213), .A2(n212), .A3(n211), .ZN(N371) );
  AOI22D1BWP30P140LVT U251 ( .A1(n214), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n215) );
  IOA21D1BWP30P140LVT U252 ( .A1(n216), .A2(i_data_bus[232]), .B(n215), .ZN(
        n217) );
  AOI21D1BWP30P140LVT U253 ( .A1(n7), .A2(i_data_bus[8]), .B(n217), .ZN(n221)
         );
  AOI22D1BWP30P140LVT U254 ( .A1(n218), .A2(i_data_bus[72]), .B1(n6), .B2(
        i_data_bus[40]), .ZN(n220) );
  AOI22D1BWP30P140LVT U255 ( .A1(n2), .A2(i_data_bus[104]), .B1(n3), .B2(
        i_data_bus[136]), .ZN(n219) );
  ND3D1BWP30P140LVT U256 ( .A1(n221), .A2(n220), .A3(n219), .ZN(N377) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_2 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD6BWP30P140LVT U3 ( .I(n51), .ZN(n1) );
  NR2D1BWP30P140LVT U4 ( .A1(n30), .A2(i_cmd[1]), .ZN(n5) );
  CKND2D3BWP30P140LVT U5 ( .A1(n11), .A2(n10), .ZN(n17) );
  NR2OPTPAD1BWP30P140LVT U6 ( .A1(n9), .A2(rst), .ZN(n11) );
  INR2D2BWP30P140LVT U7 ( .A1(i_en), .B1(n32), .ZN(n10) );
  CKND2D2BWP30P140LVT U8 ( .A1(n8), .A2(n7), .ZN(n9) );
  INVD1BWP30P140LVT U9 ( .I(n45), .ZN(n228) );
  CKND2D3BWP30P140LVT U10 ( .A1(n4), .A2(n3), .ZN(n24) );
  ND3D2BWP30P140LVT U11 ( .A1(n38), .A2(i_cmd[0]), .A3(n6), .ZN(n45) );
  INR2D2BWP30P140LVT U12 ( .A1(n15), .B1(n17), .ZN(n43) );
  INVD2BWP30P140LVT U13 ( .I(n39), .ZN(n51) );
  INVD1BWP30P140LVT U14 ( .I(i_cmd[1]), .ZN(n27) );
  INVD1BWP30P140LVT U15 ( .I(n32), .ZN(n33) );
  INR2D1BWP30P140LVT U16 ( .A1(n38), .B1(n37), .ZN(n39) );
  OAI211D1BWP30P140LVT U17 ( .A1(n22), .A2(n21), .B(n20), .C(n19), .ZN(n23) );
  ND2D1BWP30P140LVT U18 ( .A1(n223), .A2(i_data_bus[175]), .ZN(n19) );
  INVD1BWP30P140LVT U19 ( .I(i_cmd[3]), .ZN(n26) );
  NR2D1BWP30P140LVT U20 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n25) );
  ND2OPTIBD1BWP30P140LVT U21 ( .A1(n109), .A2(n108), .ZN(n110) );
  ND2D1BWP30P140LVT U22 ( .A1(n176), .A2(i_data_bus[169]), .ZN(n109) );
  AOI22D1BWP30P140LVT U23 ( .A1(n114), .A2(i_data_bus[201]), .B1(n226), .B2(
        i_data_bus[233]), .ZN(n108) );
  INVD1BWP30P140LVT U24 ( .I(n50), .ZN(n136) );
  AOI22D1BWP30P140LVT U25 ( .A1(n224), .A2(i_data_bus[210]), .B1(n223), .B2(
        i_data_bus[178]), .ZN(n198) );
  AOI21D1BWP30P140LVT U26 ( .A1(n228), .A2(i_data_bus[14]), .B(n116), .ZN(n119) );
  ND3D1BWP30P140LVT U27 ( .A1(n42), .A2(n41), .A3(n40), .ZN(N384) );
  AOI21D1BWP30P140LVT U28 ( .A1(n228), .A2(i_data_bus[15]), .B(n23), .ZN(n42)
         );
  AOI21D1BWP30P140LVT U29 ( .A1(n228), .A2(i_data_bus[16]), .B(n209), .ZN(n212) );
  AOI21D1BWP30P140LVT U30 ( .A1(n228), .A2(i_data_bus[17]), .B(n204), .ZN(n207) );
  INVD1BWP30P140LVT U31 ( .I(n29), .ZN(n55) );
  INVD1BWP30P140LVT U32 ( .I(n36), .ZN(n56) );
  NR2D3BWP30P140LVT U33 ( .A1(n17), .A2(n13), .ZN(n226) );
  AN3D1BWP30P140LVT U34 ( .A1(n31), .A2(i_cmd[1]), .A3(i_valid[1]), .Z(n2) );
  OR2D4BWP30P140LVT U35 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n30) );
  NR3OPTPAD2BWP30P140LVT U36 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .A3(i_cmd[6]), 
        .ZN(n4) );
  INR2D1BWP30P140LVT U37 ( .A1(i_en), .B1(rst), .ZN(n3) );
  INR2D2BWP30P140LVT U38 ( .A1(n5), .B1(n24), .ZN(n38) );
  INR2D1BWP30P140LVT U39 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n6) );
  NR2OPTPAD2BWP30P140LVT U40 ( .A1(i_cmd[3]), .A2(i_cmd[4]), .ZN(n8) );
  INVD2BWP30P140LVT U41 ( .I(i_cmd[0]), .ZN(n7) );
  OR2D4BWP30P140LVT U42 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .Z(n32) );
  ND2D1BWP30P140LVT U43 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n12) );
  OR3D1BWP30P140LVT U44 ( .A1(n12), .A2(i_cmd[5]), .A3(i_cmd[6]), .Z(n13) );
  INVD1BWP30P140LVT U45 ( .I(n226), .ZN(n22) );
  INVD1BWP30P140LVT U46 ( .I(i_data_bus[239]), .ZN(n21) );
  ND2D1BWP30P140LVT U47 ( .A1(i_valid[6]), .A2(i_cmd[6]), .ZN(n14) );
  NR3D0P7BWP30P140LVT U48 ( .A1(n14), .A2(i_cmd[5]), .A3(i_cmd[7]), .ZN(n15)
         );
  BUFFD2BWP30P140LVT U49 ( .I(n43), .Z(n114) );
  ND2D1BWP30P140LVT U50 ( .A1(n114), .A2(i_data_bus[207]), .ZN(n20) );
  INVD1BWP30P140LVT U51 ( .I(i_cmd[5]), .ZN(n16) );
  INR4D1BWP30P140LVT U52 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n16), .ZN(n18) );
  INR2D2BWP30P140LVT U53 ( .A1(n18), .B1(n17), .ZN(n60) );
  BUFFD4BWP30P140LVT U54 ( .I(n60), .Z(n223) );
  INR2D2BWP30P140LVT U55 ( .A1(n25), .B1(n24), .ZN(n35) );
  ND4D1BWP30P140LVT U56 ( .A1(n27), .A2(n26), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n28) );
  INR2D1BWP30P140LVT U57 ( .A1(n35), .B1(n28), .ZN(n29) );
  INVD2BWP30P140LVT U58 ( .I(n55), .ZN(n230) );
  INVD1BWP30P140LVT U59 ( .I(n30), .ZN(n31) );
  ND2OPTIBD2BWP30P140LVT U60 ( .A1(n2), .A2(n35), .ZN(n50) );
  INVD2BWP30P140LVT U61 ( .I(n50), .ZN(n229) );
  AOI22D1BWP30P140LVT U62 ( .A1(n230), .A2(i_data_bus[79]), .B1(n229), .B2(
        i_data_bus[47]), .ZN(n41) );
  ND3D1BWP30P140LVT U63 ( .A1(n33), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n34)
         );
  INR2D1BWP30P140LVT U64 ( .A1(n35), .B1(n34), .ZN(n36) );
  INVD2BWP30P140LVT U65 ( .I(n56), .ZN(n231) );
  IND3D1BWP30P140LVT U66 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n37) );
  AOI22D1BWP30P140LVT U67 ( .A1(n231), .A2(i_data_bus[111]), .B1(n1), .B2(
        i_data_bus[143]), .ZN(n40) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[224]), .ZN(n49) );
  INVD2BWP30P140LVT U69 ( .I(n43), .ZN(n175) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[192]), .ZN(n44) );
  MAOI22D1BWP30P140LVT U71 ( .A1(n223), .A2(i_data_bus[160]), .B1(n175), .B2(
        n44), .ZN(n48) );
  INR2D1BWP30P140LVT U72 ( .A1(i_data_bus[0]), .B1(n45), .ZN(n46) );
  INVD1BWP30P140LVT U73 ( .I(n46), .ZN(n47) );
  OA211D1BWP30P140LVT U74 ( .A1(n22), .A2(n49), .B(n48), .C(n47), .Z(n54) );
  INVD2BWP30P140LVT U75 ( .I(n55), .ZN(n137) );
  AOI22D1BWP30P140LVT U76 ( .A1(n137), .A2(i_data_bus[64]), .B1(n229), .B2(
        i_data_bus[32]), .ZN(n53) );
  INVD2BWP30P140LVT U77 ( .I(n56), .ZN(n138) );
  AOI22D1BWP30P140LVT U78 ( .A1(n138), .A2(i_data_bus[96]), .B1(n1), .B2(
        i_data_bus[128]), .ZN(n52) );
  ND3D1BWP30P140LVT U79 ( .A1(n54), .A2(n53), .A3(n52), .ZN(N369) );
  INVD1BWP30P140LVT U80 ( .I(n45), .ZN(n179) );
  BUFFD4BWP30P140LVT U81 ( .I(n60), .Z(n176) );
  NR4D0BWP30P140LVT U82 ( .A1(n179), .A2(n226), .A3(n114), .A4(n176), .ZN(n59)
         );
  NR2D1BWP30P140LVT U83 ( .A1(n137), .A2(n229), .ZN(n58) );
  NR2D1BWP30P140LVT U84 ( .A1(n231), .A2(n1), .ZN(n57) );
  ND3D1BWP30P140LVT U85 ( .A1(n59), .A2(n58), .A3(n57), .ZN(N402) );
  INVD1BWP30P140LVT U86 ( .I(n60), .ZN(n62) );
  INVD1BWP30P140LVT U87 ( .I(i_data_bus[173]), .ZN(n61) );
  MAOI22D1BWP30P140LVT U88 ( .A1(n114), .A2(i_data_bus[205]), .B1(n62), .B2(
        n61), .ZN(n63) );
  IOA21D1BWP30P140LVT U89 ( .A1(n226), .A2(i_data_bus[237]), .B(n63), .ZN(n64)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n228), .A2(i_data_bus[13]), .B(n64), .ZN(n67)
         );
  AOI22D1BWP30P140LVT U91 ( .A1(n230), .A2(i_data_bus[77]), .B1(n229), .B2(
        i_data_bus[45]), .ZN(n66) );
  AOI22D1BWP30P140LVT U92 ( .A1(n231), .A2(i_data_bus[109]), .B1(n1), .B2(
        i_data_bus[141]), .ZN(n65) );
  ND3D1BWP30P140LVT U93 ( .A1(n67), .A2(n66), .A3(n65), .ZN(N382) );
  INVD2BWP30P140LVT U94 ( .I(n45), .ZN(n135) );
  AOI22D1BWP30P140LVT U95 ( .A1(n114), .A2(i_data_bus[198]), .B1(n176), .B2(
        i_data_bus[166]), .ZN(n68) );
  IOA21D1BWP30P140LVT U96 ( .A1(n226), .A2(i_data_bus[230]), .B(n68), .ZN(n69)
         );
  AOI21D1BWP30P140LVT U97 ( .A1(n135), .A2(i_data_bus[6]), .B(n69), .ZN(n72)
         );
  AOI22D1BWP30P140LVT U98 ( .A1(n137), .A2(i_data_bus[70]), .B1(n136), .B2(
        i_data_bus[38]), .ZN(n71) );
  AOI22D1BWP30P140LVT U99 ( .A1(n138), .A2(i_data_bus[102]), .B1(n1), .B2(
        i_data_bus[134]), .ZN(n70) );
  ND3D1BWP30P140LVT U100 ( .A1(n72), .A2(n71), .A3(n70), .ZN(N375) );
  AOI22D1BWP30P140LVT U101 ( .A1(n114), .A2(i_data_bus[200]), .B1(n176), .B2(
        i_data_bus[168]), .ZN(n73) );
  IOA21D1BWP30P140LVT U102 ( .A1(n226), .A2(i_data_bus[232]), .B(n73), .ZN(n74) );
  AOI21D1BWP30P140LVT U103 ( .A1(n135), .A2(i_data_bus[8]), .B(n74), .ZN(n77)
         );
  AOI22D1BWP30P140LVT U104 ( .A1(n137), .A2(i_data_bus[72]), .B1(n136), .B2(
        i_data_bus[40]), .ZN(n76) );
  AOI22D1BWP30P140LVT U105 ( .A1(n138), .A2(i_data_bus[104]), .B1(n1), .B2(
        i_data_bus[136]), .ZN(n75) );
  ND3D1BWP30P140LVT U106 ( .A1(n77), .A2(n76), .A3(n75), .ZN(N377) );
  AOI22D1BWP30P140LVT U107 ( .A1(n114), .A2(i_data_bus[202]), .B1(n176), .B2(
        i_data_bus[170]), .ZN(n78) );
  IOA21D1BWP30P140LVT U108 ( .A1(n226), .A2(i_data_bus[234]), .B(n78), .ZN(n79) );
  AOI21D1BWP30P140LVT U109 ( .A1(n135), .A2(i_data_bus[10]), .B(n79), .ZN(n82)
         );
  AOI22D1BWP30P140LVT U110 ( .A1(n137), .A2(i_data_bus[74]), .B1(n136), .B2(
        i_data_bus[42]), .ZN(n81) );
  AOI22D1BWP30P140LVT U111 ( .A1(n138), .A2(i_data_bus[106]), .B1(n1), .B2(
        i_data_bus[138]), .ZN(n80) );
  ND3D1BWP30P140LVT U112 ( .A1(n82), .A2(n81), .A3(n80), .ZN(N379) );
  AOI22D1BWP30P140LVT U113 ( .A1(n114), .A2(i_data_bus[196]), .B1(n176), .B2(
        i_data_bus[164]), .ZN(n83) );
  IOA21D1BWP30P140LVT U114 ( .A1(n226), .A2(i_data_bus[228]), .B(n83), .ZN(n84) );
  AOI21D1BWP30P140LVT U115 ( .A1(n135), .A2(i_data_bus[4]), .B(n84), .ZN(n87)
         );
  AOI22D1BWP30P140LVT U116 ( .A1(n137), .A2(i_data_bus[68]), .B1(n136), .B2(
        i_data_bus[36]), .ZN(n86) );
  AOI22D1BWP30P140LVT U117 ( .A1(n138), .A2(i_data_bus[100]), .B1(n1), .B2(
        i_data_bus[132]), .ZN(n85) );
  ND3D1BWP30P140LVT U118 ( .A1(n87), .A2(n86), .A3(n85), .ZN(N373) );
  AOI22D1BWP30P140LVT U119 ( .A1(n114), .A2(i_data_bus[199]), .B1(n176), .B2(
        i_data_bus[167]), .ZN(n88) );
  IOA21D1BWP30P140LVT U120 ( .A1(n226), .A2(i_data_bus[231]), .B(n88), .ZN(n89) );
  AOI21D1BWP30P140LVT U121 ( .A1(n135), .A2(i_data_bus[7]), .B(n89), .ZN(n92)
         );
  AOI22D1BWP30P140LVT U122 ( .A1(n137), .A2(i_data_bus[71]), .B1(n136), .B2(
        i_data_bus[39]), .ZN(n91) );
  AOI22D1BWP30P140LVT U123 ( .A1(n138), .A2(i_data_bus[103]), .B1(n1), .B2(
        i_data_bus[135]), .ZN(n90) );
  ND3D1BWP30P140LVT U124 ( .A1(n92), .A2(n91), .A3(n90), .ZN(N376) );
  AOI22D1BWP30P140LVT U125 ( .A1(n114), .A2(i_data_bus[204]), .B1(n176), .B2(
        i_data_bus[172]), .ZN(n93) );
  IOA21D1BWP30P140LVT U126 ( .A1(n226), .A2(i_data_bus[236]), .B(n93), .ZN(n94) );
  AOI21D1BWP30P140LVT U127 ( .A1(n135), .A2(i_data_bus[12]), .B(n94), .ZN(n97)
         );
  AOI22D1BWP30P140LVT U128 ( .A1(n137), .A2(i_data_bus[76]), .B1(n136), .B2(
        i_data_bus[44]), .ZN(n96) );
  AOI22D1BWP30P140LVT U129 ( .A1(n138), .A2(i_data_bus[108]), .B1(n1), .B2(
        i_data_bus[140]), .ZN(n95) );
  ND3D1BWP30P140LVT U130 ( .A1(n97), .A2(n96), .A3(n95), .ZN(N381) );
  AOI22D1BWP30P140LVT U131 ( .A1(n114), .A2(i_data_bus[203]), .B1(n176), .B2(
        i_data_bus[171]), .ZN(n98) );
  IOA21D1BWP30P140LVT U132 ( .A1(n226), .A2(i_data_bus[235]), .B(n98), .ZN(n99) );
  AOI21D1BWP30P140LVT U133 ( .A1(n135), .A2(i_data_bus[11]), .B(n99), .ZN(n102) );
  AOI22D1BWP30P140LVT U134 ( .A1(n137), .A2(i_data_bus[75]), .B1(n136), .B2(
        i_data_bus[43]), .ZN(n101) );
  AOI22D1BWP30P140LVT U135 ( .A1(n138), .A2(i_data_bus[107]), .B1(n1), .B2(
        i_data_bus[139]), .ZN(n100) );
  ND3D1BWP30P140LVT U136 ( .A1(n102), .A2(n101), .A3(n100), .ZN(N380) );
  AOI22D1BWP30P140LVT U137 ( .A1(n114), .A2(i_data_bus[197]), .B1(n176), .B2(
        i_data_bus[165]), .ZN(n103) );
  IOA21D1BWP30P140LVT U138 ( .A1(n226), .A2(i_data_bus[229]), .B(n103), .ZN(
        n104) );
  AOI21D1BWP30P140LVT U139 ( .A1(n135), .A2(i_data_bus[5]), .B(n104), .ZN(n107) );
  AOI22D1BWP30P140LVT U140 ( .A1(n137), .A2(i_data_bus[69]), .B1(n136), .B2(
        i_data_bus[37]), .ZN(n106) );
  AOI22D1BWP30P140LVT U141 ( .A1(n138), .A2(i_data_bus[101]), .B1(n1), .B2(
        i_data_bus[133]), .ZN(n105) );
  ND3D1BWP30P140LVT U142 ( .A1(n107), .A2(n106), .A3(n105), .ZN(N374) );
  AOI21D1BWP30P140LVT U143 ( .A1(n135), .A2(i_data_bus[9]), .B(n110), .ZN(n113) );
  AOI22D1BWP30P140LVT U144 ( .A1(n137), .A2(i_data_bus[73]), .B1(n136), .B2(
        i_data_bus[41]), .ZN(n112) );
  AOI22D1BWP30P140LVT U145 ( .A1(n138), .A2(i_data_bus[105]), .B1(n1), .B2(
        i_data_bus[137]), .ZN(n111) );
  ND3D1BWP30P140LVT U146 ( .A1(n113), .A2(n112), .A3(n111), .ZN(N378) );
  AOI22D1BWP30P140LVT U147 ( .A1(n114), .A2(i_data_bus[206]), .B1(n176), .B2(
        i_data_bus[174]), .ZN(n115) );
  IOA21D1BWP30P140LVT U148 ( .A1(n226), .A2(i_data_bus[238]), .B(n115), .ZN(
        n116) );
  AOI22D1BWP30P140LVT U149 ( .A1(n230), .A2(i_data_bus[78]), .B1(n229), .B2(
        i_data_bus[46]), .ZN(n118) );
  AOI22D1BWP30P140LVT U150 ( .A1(n231), .A2(i_data_bus[110]), .B1(n1), .B2(
        i_data_bus[142]), .ZN(n117) );
  ND3D1BWP30P140LVT U151 ( .A1(n119), .A2(n118), .A3(n117), .ZN(N383) );
  INVD1BWP30P140LVT U152 ( .I(i_data_bus[193]), .ZN(n120) );
  MAOI22D1BWP30P140LVT U153 ( .A1(n176), .A2(i_data_bus[161]), .B1(n175), .B2(
        n120), .ZN(n121) );
  IOA21D1BWP30P140LVT U154 ( .A1(n226), .A2(i_data_bus[225]), .B(n121), .ZN(
        n122) );
  AOI21D1BWP30P140LVT U155 ( .A1(n135), .A2(i_data_bus[1]), .B(n122), .ZN(n125) );
  AOI22D1BWP30P140LVT U156 ( .A1(n137), .A2(i_data_bus[65]), .B1(n136), .B2(
        i_data_bus[33]), .ZN(n124) );
  AOI22D1BWP30P140LVT U157 ( .A1(n138), .A2(i_data_bus[97]), .B1(n1), .B2(
        i_data_bus[129]), .ZN(n123) );
  ND3D1BWP30P140LVT U158 ( .A1(n125), .A2(n124), .A3(n123), .ZN(N370) );
  INVD1BWP30P140LVT U159 ( .I(i_data_bus[194]), .ZN(n126) );
  MAOI22D1BWP30P140LVT U160 ( .A1(n176), .A2(i_data_bus[162]), .B1(n175), .B2(
        n126), .ZN(n127) );
  IOA21D1BWP30P140LVT U161 ( .A1(n226), .A2(i_data_bus[226]), .B(n127), .ZN(
        n128) );
  AOI21D1BWP30P140LVT U162 ( .A1(n135), .A2(i_data_bus[2]), .B(n128), .ZN(n131) );
  AOI22D1BWP30P140LVT U163 ( .A1(n137), .A2(i_data_bus[66]), .B1(n136), .B2(
        i_data_bus[34]), .ZN(n130) );
  AOI22D1BWP30P140LVT U164 ( .A1(n138), .A2(i_data_bus[98]), .B1(n1), .B2(
        i_data_bus[130]), .ZN(n129) );
  ND3D1BWP30P140LVT U165 ( .A1(n131), .A2(n130), .A3(n129), .ZN(N371) );
  INVD1BWP30P140LVT U166 ( .I(i_data_bus[195]), .ZN(n132) );
  MAOI22D1BWP30P140LVT U167 ( .A1(n176), .A2(i_data_bus[163]), .B1(n175), .B2(
        n132), .ZN(n133) );
  IOA21D1BWP30P140LVT U168 ( .A1(n226), .A2(i_data_bus[227]), .B(n133), .ZN(
        n134) );
  AOI21D1BWP30P140LVT U169 ( .A1(n135), .A2(i_data_bus[3]), .B(n134), .ZN(n141) );
  AOI22D1BWP30P140LVT U170 ( .A1(n137), .A2(i_data_bus[67]), .B1(n136), .B2(
        i_data_bus[35]), .ZN(n140) );
  AOI22D1BWP30P140LVT U171 ( .A1(n138), .A2(i_data_bus[99]), .B1(n1), .B2(
        i_data_bus[131]), .ZN(n139) );
  ND3D1BWP30P140LVT U172 ( .A1(n141), .A2(n140), .A3(n139), .ZN(N372) );
  INVD2BWP30P140LVT U173 ( .I(n175), .ZN(n224) );
  AOI22D1BWP30P140LVT U174 ( .A1(n224), .A2(i_data_bus[218]), .B1(n223), .B2(
        i_data_bus[186]), .ZN(n142) );
  IOA21D1BWP30P140LVT U175 ( .A1(n226), .A2(i_data_bus[250]), .B(n142), .ZN(
        n143) );
  AOI21D1BWP30P140LVT U176 ( .A1(n179), .A2(i_data_bus[26]), .B(n143), .ZN(
        n146) );
  AOI22D1BWP30P140LVT U177 ( .A1(n137), .A2(i_data_bus[90]), .B1(n229), .B2(
        i_data_bus[58]), .ZN(n145) );
  AOI22D1BWP30P140LVT U178 ( .A1(n138), .A2(i_data_bus[122]), .B1(n1), .B2(
        i_data_bus[154]), .ZN(n144) );
  ND3D1BWP30P140LVT U179 ( .A1(n146), .A2(n145), .A3(n144), .ZN(N395) );
  INVD1BWP30P140LVT U180 ( .I(i_data_bus[223]), .ZN(n147) );
  MAOI22D1BWP30P140LVT U181 ( .A1(n176), .A2(i_data_bus[191]), .B1(n175), .B2(
        n147), .ZN(n148) );
  IOA21D1BWP30P140LVT U182 ( .A1(n226), .A2(i_data_bus[255]), .B(n148), .ZN(
        n149) );
  AOI21D1BWP30P140LVT U183 ( .A1(n179), .A2(i_data_bus[31]), .B(n149), .ZN(
        n152) );
  AOI22D1BWP30P140LVT U184 ( .A1(n137), .A2(i_data_bus[95]), .B1(n229), .B2(
        i_data_bus[63]), .ZN(n151) );
  AOI22D1BWP30P140LVT U185 ( .A1(n138), .A2(i_data_bus[127]), .B1(n1), .B2(
        i_data_bus[159]), .ZN(n150) );
  ND3D1BWP30P140LVT U186 ( .A1(n152), .A2(n151), .A3(n150), .ZN(N400) );
  INVD1BWP30P140LVT U187 ( .I(i_data_bus[222]), .ZN(n153) );
  MAOI22D1BWP30P140LVT U188 ( .A1(n176), .A2(i_data_bus[190]), .B1(n175), .B2(
        n153), .ZN(n154) );
  IOA21D1BWP30P140LVT U189 ( .A1(n226), .A2(i_data_bus[254]), .B(n154), .ZN(
        n155) );
  AOI21D1BWP30P140LVT U190 ( .A1(n179), .A2(i_data_bus[30]), .B(n155), .ZN(
        n158) );
  AOI22D1BWP30P140LVT U191 ( .A1(n137), .A2(i_data_bus[94]), .B1(n229), .B2(
        i_data_bus[62]), .ZN(n157) );
  AOI22D1BWP30P140LVT U192 ( .A1(n138), .A2(i_data_bus[126]), .B1(n1), .B2(
        i_data_bus[158]), .ZN(n156) );
  ND3D1BWP30P140LVT U193 ( .A1(n158), .A2(n157), .A3(n156), .ZN(N399) );
  AOI22D1BWP30P140LVT U194 ( .A1(n224), .A2(i_data_bus[217]), .B1(n223), .B2(
        i_data_bus[185]), .ZN(n159) );
  IOA21D1BWP30P140LVT U195 ( .A1(n226), .A2(i_data_bus[249]), .B(n159), .ZN(
        n160) );
  AOI21D1BWP30P140LVT U196 ( .A1(n179), .A2(i_data_bus[25]), .B(n160), .ZN(
        n163) );
  AOI22D1BWP30P140LVT U197 ( .A1(n230), .A2(i_data_bus[89]), .B1(n229), .B2(
        i_data_bus[57]), .ZN(n162) );
  AOI22D1BWP30P140LVT U198 ( .A1(n231), .A2(i_data_bus[121]), .B1(n1), .B2(
        i_data_bus[153]), .ZN(n161) );
  ND3D1BWP30P140LVT U199 ( .A1(n163), .A2(n162), .A3(n161), .ZN(N394) );
  AOI22D1BWP30P140LVT U200 ( .A1(n224), .A2(i_data_bus[220]), .B1(n223), .B2(
        i_data_bus[188]), .ZN(n164) );
  IOA21D1BWP30P140LVT U201 ( .A1(n226), .A2(i_data_bus[252]), .B(n164), .ZN(
        n165) );
  AOI21D1BWP30P140LVT U202 ( .A1(n179), .A2(i_data_bus[28]), .B(n165), .ZN(
        n168) );
  AOI22D1BWP30P140LVT U203 ( .A1(n230), .A2(i_data_bus[92]), .B1(n229), .B2(
        i_data_bus[60]), .ZN(n167) );
  AOI22D1BWP30P140LVT U204 ( .A1(n138), .A2(i_data_bus[124]), .B1(n1), .B2(
        i_data_bus[156]), .ZN(n166) );
  ND3D1BWP30P140LVT U205 ( .A1(n168), .A2(n167), .A3(n166), .ZN(N397) );
  AOI22D1BWP30P140LVT U206 ( .A1(n224), .A2(i_data_bus[219]), .B1(n223), .B2(
        i_data_bus[187]), .ZN(n169) );
  IOA21D1BWP30P140LVT U207 ( .A1(n226), .A2(i_data_bus[251]), .B(n169), .ZN(
        n170) );
  AOI21D1BWP30P140LVT U208 ( .A1(n179), .A2(i_data_bus[27]), .B(n170), .ZN(
        n173) );
  AOI22D1BWP30P140LVT U209 ( .A1(n137), .A2(i_data_bus[91]), .B1(n229), .B2(
        i_data_bus[59]), .ZN(n172) );
  AOI22D1BWP30P140LVT U210 ( .A1(n231), .A2(i_data_bus[123]), .B1(n1), .B2(
        i_data_bus[155]), .ZN(n171) );
  ND3D1BWP30P140LVT U211 ( .A1(n173), .A2(n172), .A3(n171), .ZN(N396) );
  INVD1BWP30P140LVT U212 ( .I(i_data_bus[221]), .ZN(n174) );
  MAOI22D1BWP30P140LVT U213 ( .A1(n176), .A2(i_data_bus[189]), .B1(n175), .B2(
        n174), .ZN(n177) );
  IOA21D1BWP30P140LVT U214 ( .A1(n226), .A2(i_data_bus[253]), .B(n177), .ZN(
        n178) );
  AOI21D1BWP30P140LVT U215 ( .A1(n179), .A2(i_data_bus[29]), .B(n178), .ZN(
        n182) );
  AOI22D1BWP30P140LVT U216 ( .A1(n230), .A2(i_data_bus[93]), .B1(n229), .B2(
        i_data_bus[61]), .ZN(n181) );
  AOI22D1BWP30P140LVT U217 ( .A1(n138), .A2(i_data_bus[125]), .B1(n1), .B2(
        i_data_bus[157]), .ZN(n180) );
  ND3D1BWP30P140LVT U218 ( .A1(n182), .A2(n181), .A3(n180), .ZN(N398) );
  AOI22D1BWP30P140LVT U219 ( .A1(n224), .A2(i_data_bus[214]), .B1(n223), .B2(
        i_data_bus[182]), .ZN(n183) );
  IOA21D1BWP30P140LVT U220 ( .A1(n226), .A2(i_data_bus[246]), .B(n183), .ZN(
        n184) );
  AOI21D1BWP30P140LVT U221 ( .A1(n228), .A2(i_data_bus[22]), .B(n184), .ZN(
        n187) );
  AOI22D1BWP30P140LVT U222 ( .A1(n230), .A2(i_data_bus[86]), .B1(n229), .B2(
        i_data_bus[54]), .ZN(n186) );
  AOI22D1BWP30P140LVT U223 ( .A1(n231), .A2(i_data_bus[118]), .B1(n1), .B2(
        i_data_bus[150]), .ZN(n185) );
  ND3D1BWP30P140LVT U224 ( .A1(n187), .A2(n186), .A3(n185), .ZN(N391) );
  AOI22D1BWP30P140LVT U225 ( .A1(n224), .A2(i_data_bus[213]), .B1(n223), .B2(
        i_data_bus[181]), .ZN(n188) );
  IOA21D1BWP30P140LVT U226 ( .A1(n226), .A2(i_data_bus[245]), .B(n188), .ZN(
        n189) );
  AOI21D1BWP30P140LVT U227 ( .A1(n228), .A2(i_data_bus[21]), .B(n189), .ZN(
        n192) );
  AOI22D1BWP30P140LVT U228 ( .A1(n230), .A2(i_data_bus[85]), .B1(n229), .B2(
        i_data_bus[53]), .ZN(n191) );
  AOI22D1BWP30P140LVT U229 ( .A1(n231), .A2(i_data_bus[117]), .B1(n1), .B2(
        i_data_bus[149]), .ZN(n190) );
  ND3D1BWP30P140LVT U230 ( .A1(n192), .A2(n191), .A3(n190), .ZN(N390) );
  AOI22D1BWP30P140LVT U231 ( .A1(n224), .A2(i_data_bus[212]), .B1(n223), .B2(
        i_data_bus[180]), .ZN(n193) );
  IOA21D1BWP30P140LVT U232 ( .A1(n226), .A2(i_data_bus[244]), .B(n193), .ZN(
        n194) );
  AOI21D1BWP30P140LVT U233 ( .A1(n228), .A2(i_data_bus[20]), .B(n194), .ZN(
        n197) );
  AOI22D1BWP30P140LVT U234 ( .A1(n230), .A2(i_data_bus[84]), .B1(n229), .B2(
        i_data_bus[52]), .ZN(n196) );
  AOI22D1BWP30P140LVT U235 ( .A1(n231), .A2(i_data_bus[116]), .B1(n1), .B2(
        i_data_bus[148]), .ZN(n195) );
  ND3D1BWP30P140LVT U236 ( .A1(n197), .A2(n196), .A3(n195), .ZN(N389) );
  IOA21D1BWP30P140LVT U237 ( .A1(n226), .A2(i_data_bus[242]), .B(n198), .ZN(
        n199) );
  AOI21D1BWP30P140LVT U238 ( .A1(n228), .A2(i_data_bus[18]), .B(n199), .ZN(
        n202) );
  AOI22D1BWP30P140LVT U239 ( .A1(n230), .A2(i_data_bus[82]), .B1(n229), .B2(
        i_data_bus[50]), .ZN(n201) );
  AOI22D1BWP30P140LVT U240 ( .A1(n231), .A2(i_data_bus[114]), .B1(n1), .B2(
        i_data_bus[146]), .ZN(n200) );
  ND3D1BWP30P140LVT U241 ( .A1(n202), .A2(n201), .A3(n200), .ZN(N387) );
  AOI22D1BWP30P140LVT U242 ( .A1(n224), .A2(i_data_bus[209]), .B1(n223), .B2(
        i_data_bus[177]), .ZN(n203) );
  IOA21D1BWP30P140LVT U243 ( .A1(n226), .A2(i_data_bus[241]), .B(n203), .ZN(
        n204) );
  AOI22D1BWP30P140LVT U244 ( .A1(n230), .A2(i_data_bus[81]), .B1(n229), .B2(
        i_data_bus[49]), .ZN(n206) );
  AOI22D1BWP30P140LVT U245 ( .A1(n231), .A2(i_data_bus[113]), .B1(n1), .B2(
        i_data_bus[145]), .ZN(n205) );
  ND3D1BWP30P140LVT U246 ( .A1(n207), .A2(n206), .A3(n205), .ZN(N386) );
  AOI22D1BWP30P140LVT U247 ( .A1(n224), .A2(i_data_bus[208]), .B1(n223), .B2(
        i_data_bus[176]), .ZN(n208) );
  IOA21D1BWP30P140LVT U248 ( .A1(n226), .A2(i_data_bus[240]), .B(n208), .ZN(
        n209) );
  AOI22D1BWP30P140LVT U249 ( .A1(n230), .A2(i_data_bus[80]), .B1(n229), .B2(
        i_data_bus[48]), .ZN(n211) );
  AOI22D1BWP30P140LVT U250 ( .A1(n231), .A2(i_data_bus[112]), .B1(n1), .B2(
        i_data_bus[144]), .ZN(n210) );
  ND3D1BWP30P140LVT U251 ( .A1(n212), .A2(n211), .A3(n210), .ZN(N385) );
  AOI22D1BWP30P140LVT U252 ( .A1(n224), .A2(i_data_bus[211]), .B1(n223), .B2(
        i_data_bus[179]), .ZN(n213) );
  IOA21D1BWP30P140LVT U253 ( .A1(n226), .A2(i_data_bus[243]), .B(n213), .ZN(
        n214) );
  AOI21D1BWP30P140LVT U254 ( .A1(n228), .A2(i_data_bus[19]), .B(n214), .ZN(
        n217) );
  AOI22D1BWP30P140LVT U255 ( .A1(n230), .A2(i_data_bus[83]), .B1(n229), .B2(
        i_data_bus[51]), .ZN(n216) );
  AOI22D1BWP30P140LVT U256 ( .A1(n231), .A2(i_data_bus[115]), .B1(n1), .B2(
        i_data_bus[147]), .ZN(n215) );
  ND3D1BWP30P140LVT U257 ( .A1(n217), .A2(n216), .A3(n215), .ZN(N388) );
  AOI22D1BWP30P140LVT U258 ( .A1(n224), .A2(i_data_bus[216]), .B1(n223), .B2(
        i_data_bus[184]), .ZN(n218) );
  IOA21D1BWP30P140LVT U259 ( .A1(n226), .A2(i_data_bus[248]), .B(n218), .ZN(
        n219) );
  AOI21D1BWP30P140LVT U260 ( .A1(n228), .A2(i_data_bus[24]), .B(n219), .ZN(
        n222) );
  AOI22D1BWP30P140LVT U261 ( .A1(n230), .A2(i_data_bus[88]), .B1(n229), .B2(
        i_data_bus[56]), .ZN(n221) );
  AOI22D1BWP30P140LVT U262 ( .A1(n231), .A2(i_data_bus[120]), .B1(n1), .B2(
        i_data_bus[152]), .ZN(n220) );
  ND3D1BWP30P140LVT U263 ( .A1(n222), .A2(n221), .A3(n220), .ZN(N393) );
  AOI22D1BWP30P140LVT U264 ( .A1(n224), .A2(i_data_bus[215]), .B1(n223), .B2(
        i_data_bus[183]), .ZN(n225) );
  IOA21D1BWP30P140LVT U265 ( .A1(n226), .A2(i_data_bus[247]), .B(n225), .ZN(
        n227) );
  AOI21D1BWP30P140LVT U266 ( .A1(n228), .A2(i_data_bus[23]), .B(n227), .ZN(
        n234) );
  AOI22D1BWP30P140LVT U267 ( .A1(n230), .A2(i_data_bus[87]), .B1(n229), .B2(
        i_data_bus[55]), .ZN(n233) );
  AOI22D1BWP30P140LVT U268 ( .A1(n231), .A2(i_data_bus[119]), .B1(n1), .B2(
        i_data_bus[151]), .ZN(n232) );
  ND3D1BWP30P140LVT U269 ( .A1(n234), .A2(n233), .A3(n232), .ZN(N392) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_3 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD2BWP30P140LVT U3 ( .I(n221), .ZN(n229) );
  NR2D1BWP30P140LVT U4 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n25) );
  INR4D2BWP30P140LVT U5 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n20), .ZN(n22) );
  CKND2D3BWP30P140LVT U6 ( .A1(n16), .A2(n3), .ZN(n21) );
  INR2D1BWP30P140LVT U7 ( .A1(n4), .B1(i_cmd[6]), .ZN(n5) );
  CKND2D2BWP30P140LVT U8 ( .A1(n13), .A2(n12), .ZN(n14) );
  INVD1BWP30P140LVT U9 ( .I(i_cmd[0]), .ZN(n12) );
  ND2OPTIBD1BWP30P140LVT U10 ( .A1(n18), .A2(n5), .ZN(n24) );
  INVD4BWP30P140LVT U11 ( .I(n106), .ZN(n1) );
  INVD4BWP30P140LVT U12 ( .I(n199), .ZN(n2) );
  INR2D4BWP30P140LVT U13 ( .A1(n22), .B1(n21), .ZN(n23) );
  INR2D2BWP30P140LVT U14 ( .A1(n25), .B1(n24), .ZN(n33) );
  INR2D2BWP30P140LVT U15 ( .A1(n15), .B1(n14), .ZN(n16) );
  ND2D1BWP30P140LVT U16 ( .A1(i_valid[1]), .A2(i_cmd[1]), .ZN(n29) );
  NR2D3BWP30P140LVT U17 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .ZN(n18) );
  INVD2BWP30P140LVT U18 ( .I(n47), .ZN(n128) );
  INR2D1BWP30P140LVT U19 ( .A1(i_en), .B1(rst), .ZN(n4) );
  NR2D3BWP30P140LVT U20 ( .A1(i_cmd[3]), .A2(i_cmd[4]), .ZN(n13) );
  ND3D1BWP30P140LVT U21 ( .A1(n18), .A2(i_valid[6]), .A3(i_cmd[6]), .ZN(n19)
         );
  ND2OPTIBD1BWP30P140LVT U22 ( .A1(n37), .A2(n36), .ZN(n47) );
  INVD1BWP30P140LVT U23 ( .I(n34), .ZN(n100) );
  INR2D1BWP30P140LVT U24 ( .A1(n33), .B1(n28), .ZN(n127) );
  INVD1BWP30P140LVT U25 ( .I(i_cmd[3]), .ZN(n26) );
  INVD1BWP30P140LVT U26 ( .I(n100), .ZN(n129) );
  OAI21D1BWP30P140LVT U27 ( .A1(n106), .A2(n105), .B(n104), .ZN(n107) );
  INVD1BWP30P140LVT U28 ( .I(i_data_bus[174]), .ZN(n105) );
  ND2D1BWP30P140LVT U29 ( .A1(n226), .A2(i_data_bus[238]), .ZN(n104) );
  INR2D1BWP30P140LVT U30 ( .A1(i_data_bus[206]), .B1(n199), .ZN(n108) );
  INVD1BWP30P140LVT U31 ( .I(n127), .ZN(n221) );
  INVD1BWP30P140LVT U32 ( .I(n100), .ZN(n231) );
  INVD2BWP30P140LVT U33 ( .I(n47), .ZN(n230) );
  INVD1BWP30P140LVT U34 ( .I(n100), .ZN(n169) );
  INVD2BWP30P140LVT U35 ( .I(n221), .ZN(n168) );
  INVD1BWP30P140LVT U36 ( .I(i_en), .ZN(n11) );
  NR2D1BWP30P140LVT U37 ( .A1(n6), .A2(n24), .ZN(n37) );
  NR2D1BWP30P140LVT U38 ( .A1(n11), .A2(rst), .ZN(n15) );
  OR2D1BWP30P140LVT U39 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n30) );
  INVD1BWP30P140LVT U40 ( .I(n226), .ZN(n46) );
  ND2OPTIBD1BWP30P140LVT U41 ( .A1(n33), .A2(n31), .ZN(n219) );
  NR2D1BWP30P140LVT U42 ( .A1(n30), .A2(n29), .ZN(n31) );
  AOI21D1BWP30P140LVT U43 ( .A1(n217), .A2(i_data_bus[3]), .B(n126), .ZN(n132)
         );
  AOI211D1BWP30P140LVT U44 ( .A1(n217), .A2(i_data_bus[14]), .B(n108), .C(n107), .ZN(n111) );
  AOI21D1BWP30P140LVT U45 ( .A1(n217), .A2(i_data_bus[29]), .B(n157), .ZN(n160) );
  ND2OPTIBD1BWP30P140LVT U46 ( .A1(n37), .A2(n9), .ZN(n61) );
  NR2D1BWP30P140LVT U47 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n3) );
  OR2D1BWP30P140LVT U48 ( .A1(n30), .A2(i_cmd[1]), .Z(n6) );
  INR2D1BWP30P140LVT U49 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n7) );
  INVD1BWP30P140LVT U50 ( .I(n7), .ZN(n8) );
  NR2D1BWP30P140LVT U51 ( .A1(n8), .A2(n12), .ZN(n9) );
  ND2D1BWP30P140LVT U52 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n10) );
  NR3D0P7BWP30P140LVT U53 ( .A1(n10), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n17)
         );
  INR2D4BWP30P140LVT U54 ( .A1(n17), .B1(n21), .ZN(n226) );
  OR2D4BWP30P140LVT U55 ( .A1(n21), .A2(n19), .Z(n199) );
  INVD1BWP30P140LVT U56 ( .I(i_cmd[5]), .ZN(n20) );
  INVD3BWP30P140LVT U57 ( .I(n23), .ZN(n106) );
  NR4D0BWP30P140LVT U58 ( .A1(n217), .A2(n226), .A3(n2), .A4(n1), .ZN(n40) );
  INVD1BWP30P140LVT U59 ( .I(i_cmd[1]), .ZN(n27) );
  ND4D1BWP30P140LVT U60 ( .A1(n27), .A2(n26), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n28) );
  INVD2BWP30P140LVT U61 ( .I(n219), .ZN(n228) );
  NR2D1BWP30P140LVT U62 ( .A1(n168), .A2(n228), .ZN(n39) );
  ND3D1BWP30P140LVT U63 ( .A1(n3), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n32) );
  INR2D1BWP30P140LVT U64 ( .A1(n33), .B1(n32), .ZN(n34) );
  IND3D1BWP30P140LVT U65 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n35) );
  INVD1BWP30P140LVT U66 ( .I(n35), .ZN(n36) );
  NR2D1BWP30P140LVT U67 ( .A1(n169), .A2(n230), .ZN(n38) );
  ND3D1BWP30P140LVT U68 ( .A1(n40), .A2(n39), .A3(n38), .ZN(N402) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[224]), .ZN(n45) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[192]), .ZN(n41) );
  MAOI22D1BWP30P140LVT U71 ( .A1(n1), .A2(i_data_bus[160]), .B1(n199), .B2(n41), .ZN(n44) );
  INR2D1BWP30P140LVT U72 ( .A1(i_data_bus[0]), .B1(n61), .ZN(n42) );
  INVD1BWP30P140LVT U73 ( .I(n42), .ZN(n43) );
  OA211D1BWP30P140LVT U74 ( .A1(n46), .A2(n45), .B(n44), .C(n43), .Z(n50) );
  AOI22D1BWP30P140LVT U75 ( .A1(n168), .A2(i_data_bus[64]), .B1(n228), .B2(
        i_data_bus[32]), .ZN(n49) );
  AOI22D1BWP30P140LVT U76 ( .A1(n129), .A2(i_data_bus[96]), .B1(n128), .B2(
        i_data_bus[128]), .ZN(n48) );
  ND3D1BWP30P140LVT U77 ( .A1(n50), .A2(n49), .A3(n48), .ZN(N369) );
  AOI22D1BWP30P140LVT U78 ( .A1(n2), .A2(i_data_bus[199]), .B1(n1), .B2(
        i_data_bus[167]), .ZN(n51) );
  IOA21D1BWP30P140LVT U79 ( .A1(n226), .A2(i_data_bus[231]), .B(n51), .ZN(n52)
         );
  AOI21D1BWP30P140LVT U80 ( .A1(n217), .A2(i_data_bus[7]), .B(n52), .ZN(n55)
         );
  AOI22D1BWP30P140LVT U81 ( .A1(n168), .A2(i_data_bus[71]), .B1(n228), .B2(
        i_data_bus[39]), .ZN(n54) );
  AOI22D1BWP30P140LVT U82 ( .A1(n129), .A2(i_data_bus[103]), .B1(n128), .B2(
        i_data_bus[135]), .ZN(n53) );
  ND3D1BWP30P140LVT U83 ( .A1(n55), .A2(n54), .A3(n53), .ZN(N376) );
  AOI22D1BWP30P140LVT U84 ( .A1(n2), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n56) );
  IOA21D1BWP30P140LVT U85 ( .A1(n226), .A2(i_data_bus[233]), .B(n56), .ZN(n57)
         );
  AOI21D1BWP30P140LVT U86 ( .A1(n217), .A2(i_data_bus[9]), .B(n57), .ZN(n60)
         );
  AOI22D1BWP30P140LVT U87 ( .A1(n168), .A2(i_data_bus[73]), .B1(n228), .B2(
        i_data_bus[41]), .ZN(n59) );
  AOI22D1BWP30P140LVT U88 ( .A1(n129), .A2(i_data_bus[105]), .B1(n128), .B2(
        i_data_bus[137]), .ZN(n58) );
  ND3D1BWP30P140LVT U89 ( .A1(n60), .A2(n59), .A3(n58), .ZN(N378) );
  INVD2BWP30P140LVT U90 ( .I(n61), .ZN(n217) );
  AOI22D1BWP30P140LVT U91 ( .A1(n2), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n62) );
  IOA21D1BWP30P140LVT U92 ( .A1(n226), .A2(i_data_bus[232]), .B(n62), .ZN(n63)
         );
  AOI21D1BWP30P140LVT U93 ( .A1(n217), .A2(i_data_bus[8]), .B(n63), .ZN(n66)
         );
  AOI22D1BWP30P140LVT U94 ( .A1(n168), .A2(i_data_bus[72]), .B1(n228), .B2(
        i_data_bus[40]), .ZN(n65) );
  AOI22D1BWP30P140LVT U95 ( .A1(n129), .A2(i_data_bus[104]), .B1(n128), .B2(
        i_data_bus[136]), .ZN(n64) );
  ND3D1BWP30P140LVT U96 ( .A1(n66), .A2(n65), .A3(n64), .ZN(N377) );
  AOI22D1BWP30P140LVT U97 ( .A1(n2), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n67) );
  IOA21D1BWP30P140LVT U98 ( .A1(n226), .A2(i_data_bus[230]), .B(n67), .ZN(n68)
         );
  AOI21D1BWP30P140LVT U99 ( .A1(n217), .A2(i_data_bus[6]), .B(n68), .ZN(n71)
         );
  AOI22D1BWP30P140LVT U100 ( .A1(n168), .A2(i_data_bus[70]), .B1(n228), .B2(
        i_data_bus[38]), .ZN(n70) );
  AOI22D1BWP30P140LVT U101 ( .A1(n129), .A2(i_data_bus[102]), .B1(n128), .B2(
        i_data_bus[134]), .ZN(n69) );
  ND3D1BWP30P140LVT U102 ( .A1(n71), .A2(n70), .A3(n69), .ZN(N375) );
  AOI22D1BWP30P140LVT U103 ( .A1(n2), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n72) );
  IOA21D1BWP30P140LVT U104 ( .A1(n226), .A2(i_data_bus[229]), .B(n72), .ZN(n73) );
  AOI21D1BWP30P140LVT U105 ( .A1(n217), .A2(i_data_bus[5]), .B(n73), .ZN(n76)
         );
  AOI22D1BWP30P140LVT U106 ( .A1(n168), .A2(i_data_bus[69]), .B1(n228), .B2(
        i_data_bus[37]), .ZN(n75) );
  AOI22D1BWP30P140LVT U107 ( .A1(n129), .A2(i_data_bus[101]), .B1(n128), .B2(
        i_data_bus[133]), .ZN(n74) );
  ND3D1BWP30P140LVT U108 ( .A1(n76), .A2(n75), .A3(n74), .ZN(N374) );
  AOI22D1BWP30P140LVT U109 ( .A1(n2), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n77) );
  IOA21D1BWP30P140LVT U110 ( .A1(n226), .A2(i_data_bus[228]), .B(n77), .ZN(n78) );
  AOI21D1BWP30P140LVT U111 ( .A1(n217), .A2(i_data_bus[4]), .B(n78), .ZN(n81)
         );
  AOI22D1BWP30P140LVT U112 ( .A1(n168), .A2(i_data_bus[68]), .B1(n228), .B2(
        i_data_bus[36]), .ZN(n80) );
  AOI22D1BWP30P140LVT U113 ( .A1(n129), .A2(i_data_bus[100]), .B1(n128), .B2(
        i_data_bus[132]), .ZN(n79) );
  ND3D1BWP30P140LVT U114 ( .A1(n81), .A2(n80), .A3(n79), .ZN(N373) );
  AOI22D1BWP30P140LVT U115 ( .A1(n2), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n82) );
  IOA21D1BWP30P140LVT U116 ( .A1(n226), .A2(i_data_bus[236]), .B(n82), .ZN(n83) );
  AOI21D1BWP30P140LVT U117 ( .A1(n217), .A2(i_data_bus[12]), .B(n83), .ZN(n86)
         );
  AOI22D1BWP30P140LVT U118 ( .A1(n229), .A2(i_data_bus[76]), .B1(n228), .B2(
        i_data_bus[44]), .ZN(n85) );
  AOI22D1BWP30P140LVT U119 ( .A1(n129), .A2(i_data_bus[108]), .B1(n128), .B2(
        i_data_bus[140]), .ZN(n84) );
  ND3D1BWP30P140LVT U120 ( .A1(n86), .A2(n85), .A3(n84), .ZN(N381) );
  AOI22D1BWP30P140LVT U121 ( .A1(n2), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n87) );
  IOA21D1BWP30P140LVT U122 ( .A1(n226), .A2(i_data_bus[234]), .B(n87), .ZN(n88) );
  AOI21D1BWP30P140LVT U123 ( .A1(n217), .A2(i_data_bus[10]), .B(n88), .ZN(n91)
         );
  AOI22D1BWP30P140LVT U124 ( .A1(n168), .A2(i_data_bus[74]), .B1(n228), .B2(
        i_data_bus[42]), .ZN(n90) );
  AOI22D1BWP30P140LVT U125 ( .A1(n129), .A2(i_data_bus[106]), .B1(n128), .B2(
        i_data_bus[138]), .ZN(n89) );
  ND3D1BWP30P140LVT U126 ( .A1(n91), .A2(n90), .A3(n89), .ZN(N379) );
  AOI22D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n92) );
  IOA21D1BWP30P140LVT U128 ( .A1(n226), .A2(i_data_bus[235]), .B(n92), .ZN(n93) );
  AOI21D1BWP30P140LVT U129 ( .A1(n217), .A2(i_data_bus[11]), .B(n93), .ZN(n96)
         );
  AOI22D1BWP30P140LVT U130 ( .A1(n229), .A2(i_data_bus[75]), .B1(n228), .B2(
        i_data_bus[43]), .ZN(n95) );
  AOI22D1BWP30P140LVT U131 ( .A1(n129), .A2(i_data_bus[107]), .B1(n128), .B2(
        i_data_bus[139]), .ZN(n94) );
  ND3D1BWP30P140LVT U132 ( .A1(n96), .A2(n95), .A3(n94), .ZN(N380) );
  INVD1BWP30P140LVT U133 ( .I(i_data_bus[173]), .ZN(n97) );
  MAOI22D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[205]), .B1(n106), .B2(
        n97), .ZN(n98) );
  IOA21D1BWP30P140LVT U135 ( .A1(n226), .A2(i_data_bus[237]), .B(n98), .ZN(n99) );
  AOI21D1BWP30P140LVT U136 ( .A1(n217), .A2(i_data_bus[13]), .B(n99), .ZN(n103) );
  AOI22D1BWP30P140LVT U137 ( .A1(n229), .A2(i_data_bus[77]), .B1(n228), .B2(
        i_data_bus[45]), .ZN(n102) );
  AOI22D1BWP30P140LVT U138 ( .A1(n231), .A2(i_data_bus[109]), .B1(n230), .B2(
        i_data_bus[141]), .ZN(n101) );
  ND3D1BWP30P140LVT U139 ( .A1(n103), .A2(n102), .A3(n101), .ZN(N382) );
  AOI22D1BWP30P140LVT U140 ( .A1(n229), .A2(i_data_bus[78]), .B1(n228), .B2(
        i_data_bus[46]), .ZN(n110) );
  AOI22D1BWP30P140LVT U141 ( .A1(n231), .A2(i_data_bus[110]), .B1(n230), .B2(
        i_data_bus[142]), .ZN(n109) );
  ND3D1BWP30P140LVT U142 ( .A1(n111), .A2(n110), .A3(n109), .ZN(N383) );
  INVD1BWP30P140LVT U143 ( .I(i_data_bus[193]), .ZN(n112) );
  MAOI22D1BWP30P140LVT U144 ( .A1(n1), .A2(i_data_bus[161]), .B1(n199), .B2(
        n112), .ZN(n113) );
  IOA21D1BWP30P140LVT U145 ( .A1(n226), .A2(i_data_bus[225]), .B(n113), .ZN(
        n114) );
  AOI21D1BWP30P140LVT U146 ( .A1(n217), .A2(i_data_bus[1]), .B(n114), .ZN(n117) );
  AOI22D1BWP30P140LVT U147 ( .A1(n168), .A2(i_data_bus[65]), .B1(n228), .B2(
        i_data_bus[33]), .ZN(n116) );
  AOI22D1BWP30P140LVT U148 ( .A1(n129), .A2(i_data_bus[97]), .B1(n128), .B2(
        i_data_bus[129]), .ZN(n115) );
  ND3D1BWP30P140LVT U149 ( .A1(n117), .A2(n116), .A3(n115), .ZN(N370) );
  INVD1BWP30P140LVT U150 ( .I(i_data_bus[194]), .ZN(n118) );
  MAOI22D1BWP30P140LVT U151 ( .A1(n1), .A2(i_data_bus[162]), .B1(n199), .B2(
        n118), .ZN(n119) );
  IOA21D1BWP30P140LVT U152 ( .A1(n226), .A2(i_data_bus[226]), .B(n119), .ZN(
        n120) );
  AOI21D1BWP30P140LVT U153 ( .A1(n217), .A2(i_data_bus[2]), .B(n120), .ZN(n123) );
  AOI22D1BWP30P140LVT U154 ( .A1(n229), .A2(i_data_bus[66]), .B1(n228), .B2(
        i_data_bus[34]), .ZN(n122) );
  AOI22D1BWP30P140LVT U155 ( .A1(n129), .A2(i_data_bus[98]), .B1(n128), .B2(
        i_data_bus[130]), .ZN(n121) );
  ND3D1BWP30P140LVT U156 ( .A1(n123), .A2(n122), .A3(n121), .ZN(N371) );
  INVD1BWP30P140LVT U157 ( .I(i_data_bus[195]), .ZN(n124) );
  MAOI22D1BWP30P140LVT U158 ( .A1(n1), .A2(i_data_bus[163]), .B1(n199), .B2(
        n124), .ZN(n125) );
  IOA21D1BWP30P140LVT U159 ( .A1(n226), .A2(i_data_bus[227]), .B(n125), .ZN(
        n126) );
  AOI22D1BWP30P140LVT U160 ( .A1(n127), .A2(i_data_bus[67]), .B1(n228), .B2(
        i_data_bus[35]), .ZN(n131) );
  AOI22D1BWP30P140LVT U161 ( .A1(n129), .A2(i_data_bus[99]), .B1(n128), .B2(
        i_data_bus[131]), .ZN(n130) );
  ND3D1BWP30P140LVT U162 ( .A1(n132), .A2(n131), .A3(n130), .ZN(N372) );
  AOI22D1BWP30P140LVT U163 ( .A1(n2), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n133) );
  IOA21D1BWP30P140LVT U164 ( .A1(n226), .A2(i_data_bus[249]), .B(n133), .ZN(
        n134) );
  AOI21D1BWP30P140LVT U165 ( .A1(n217), .A2(i_data_bus[25]), .B(n134), .ZN(
        n137) );
  AOI22D1BWP30P140LVT U166 ( .A1(n229), .A2(i_data_bus[89]), .B1(n228), .B2(
        i_data_bus[57]), .ZN(n136) );
  AOI22D1BWP30P140LVT U167 ( .A1(n231), .A2(i_data_bus[121]), .B1(n230), .B2(
        i_data_bus[153]), .ZN(n135) );
  ND3D1BWP30P140LVT U168 ( .A1(n137), .A2(n136), .A3(n135), .ZN(N394) );
  AOI22D1BWP30P140LVT U169 ( .A1(n2), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n138) );
  IOA21D1BWP30P140LVT U170 ( .A1(n226), .A2(i_data_bus[251]), .B(n138), .ZN(
        n139) );
  AOI21D1BWP30P140LVT U171 ( .A1(n217), .A2(i_data_bus[27]), .B(n139), .ZN(
        n142) );
  AOI22D1BWP30P140LVT U172 ( .A1(n168), .A2(i_data_bus[91]), .B1(n228), .B2(
        i_data_bus[59]), .ZN(n141) );
  AOI22D1BWP30P140LVT U173 ( .A1(n169), .A2(i_data_bus[123]), .B1(n230), .B2(
        i_data_bus[155]), .ZN(n140) );
  ND3D1BWP30P140LVT U174 ( .A1(n142), .A2(n141), .A3(n140), .ZN(N396) );
  INVD1BWP30P140LVT U175 ( .I(i_data_bus[223]), .ZN(n143) );
  MAOI22D1BWP30P140LVT U176 ( .A1(n1), .A2(i_data_bus[191]), .B1(n199), .B2(
        n143), .ZN(n144) );
  IOA21D1BWP30P140LVT U177 ( .A1(n226), .A2(i_data_bus[255]), .B(n144), .ZN(
        n145) );
  AOI21D1BWP30P140LVT U178 ( .A1(n217), .A2(i_data_bus[31]), .B(n145), .ZN(
        n148) );
  AOI22D1BWP30P140LVT U179 ( .A1(n168), .A2(i_data_bus[95]), .B1(n228), .B2(
        i_data_bus[63]), .ZN(n147) );
  AOI22D1BWP30P140LVT U180 ( .A1(n169), .A2(i_data_bus[127]), .B1(n230), .B2(
        i_data_bus[159]), .ZN(n146) );
  ND3D1BWP30P140LVT U181 ( .A1(n148), .A2(n147), .A3(n146), .ZN(N400) );
  INVD1BWP30P140LVT U182 ( .I(i_data_bus[222]), .ZN(n149) );
  MAOI22D1BWP30P140LVT U183 ( .A1(n1), .A2(i_data_bus[190]), .B1(n199), .B2(
        n149), .ZN(n150) );
  IOA21D1BWP30P140LVT U184 ( .A1(n226), .A2(i_data_bus[254]), .B(n150), .ZN(
        n151) );
  AOI21D1BWP30P140LVT U185 ( .A1(n217), .A2(i_data_bus[30]), .B(n151), .ZN(
        n154) );
  AOI22D1BWP30P140LVT U186 ( .A1(n168), .A2(i_data_bus[94]), .B1(n228), .B2(
        i_data_bus[62]), .ZN(n153) );
  AOI22D1BWP30P140LVT U187 ( .A1(n169), .A2(i_data_bus[126]), .B1(n230), .B2(
        i_data_bus[158]), .ZN(n152) );
  ND3D1BWP30P140LVT U188 ( .A1(n154), .A2(n153), .A3(n152), .ZN(N399) );
  INVD1BWP30P140LVT U189 ( .I(i_data_bus[221]), .ZN(n155) );
  MAOI22D1BWP30P140LVT U190 ( .A1(n1), .A2(i_data_bus[189]), .B1(n199), .B2(
        n155), .ZN(n156) );
  IOA21D1BWP30P140LVT U191 ( .A1(n226), .A2(i_data_bus[253]), .B(n156), .ZN(
        n157) );
  AOI22D1BWP30P140LVT U192 ( .A1(n168), .A2(i_data_bus[93]), .B1(n228), .B2(
        i_data_bus[61]), .ZN(n159) );
  AOI22D1BWP30P140LVT U193 ( .A1(n169), .A2(i_data_bus[125]), .B1(n230), .B2(
        i_data_bus[157]), .ZN(n158) );
  ND3D1BWP30P140LVT U194 ( .A1(n160), .A2(n159), .A3(n158), .ZN(N398) );
  AOI22D1BWP30P140LVT U195 ( .A1(n2), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n161) );
  IOA21D1BWP30P140LVT U196 ( .A1(n226), .A2(i_data_bus[250]), .B(n161), .ZN(
        n162) );
  AOI21D1BWP30P140LVT U197 ( .A1(n217), .A2(i_data_bus[26]), .B(n162), .ZN(
        n165) );
  AOI22D1BWP30P140LVT U198 ( .A1(n168), .A2(i_data_bus[90]), .B1(n228), .B2(
        i_data_bus[58]), .ZN(n164) );
  AOI22D1BWP30P140LVT U199 ( .A1(n169), .A2(i_data_bus[122]), .B1(n230), .B2(
        i_data_bus[154]), .ZN(n163) );
  ND3D1BWP30P140LVT U200 ( .A1(n165), .A2(n164), .A3(n163), .ZN(N395) );
  AOI22D1BWP30P140LVT U201 ( .A1(n2), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n166) );
  IOA21D1BWP30P140LVT U202 ( .A1(n226), .A2(i_data_bus[252]), .B(n166), .ZN(
        n167) );
  AOI21D1BWP30P140LVT U203 ( .A1(n217), .A2(i_data_bus[28]), .B(n167), .ZN(
        n172) );
  AOI22D1BWP30P140LVT U204 ( .A1(n168), .A2(i_data_bus[92]), .B1(n228), .B2(
        i_data_bus[60]), .ZN(n171) );
  AOI22D1BWP30P140LVT U205 ( .A1(n169), .A2(i_data_bus[124]), .B1(n230), .B2(
        i_data_bus[156]), .ZN(n170) );
  ND3D1BWP30P140LVT U206 ( .A1(n172), .A2(n171), .A3(n170), .ZN(N397) );
  AOI22D1BWP30P140LVT U207 ( .A1(n2), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n173) );
  IOA21D1BWP30P140LVT U208 ( .A1(n226), .A2(i_data_bus[244]), .B(n173), .ZN(
        n174) );
  AOI21D1BWP30P140LVT U209 ( .A1(n217), .A2(i_data_bus[20]), .B(n174), .ZN(
        n177) );
  AOI22D1BWP30P140LVT U210 ( .A1(n229), .A2(i_data_bus[84]), .B1(n228), .B2(
        i_data_bus[52]), .ZN(n176) );
  AOI22D1BWP30P140LVT U211 ( .A1(n231), .A2(i_data_bus[116]), .B1(n230), .B2(
        i_data_bus[148]), .ZN(n175) );
  ND3D1BWP30P140LVT U212 ( .A1(n177), .A2(n176), .A3(n175), .ZN(N389) );
  AOI22D1BWP30P140LVT U213 ( .A1(n2), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n178) );
  IOA21D1BWP30P140LVT U214 ( .A1(n226), .A2(i_data_bus[246]), .B(n178), .ZN(
        n179) );
  AOI21D1BWP30P140LVT U215 ( .A1(n217), .A2(i_data_bus[22]), .B(n179), .ZN(
        n182) );
  AOI22D1BWP30P140LVT U216 ( .A1(n229), .A2(i_data_bus[86]), .B1(n228), .B2(
        i_data_bus[54]), .ZN(n181) );
  AOI22D1BWP30P140LVT U217 ( .A1(n231), .A2(i_data_bus[118]), .B1(n230), .B2(
        i_data_bus[150]), .ZN(n180) );
  ND3D1BWP30P140LVT U218 ( .A1(n182), .A2(n181), .A3(n180), .ZN(N391) );
  AOI22D1BWP30P140LVT U219 ( .A1(n2), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n183) );
  IOA21D1BWP30P140LVT U220 ( .A1(n226), .A2(i_data_bus[243]), .B(n183), .ZN(
        n184) );
  AOI21D1BWP30P140LVT U221 ( .A1(n217), .A2(i_data_bus[19]), .B(n184), .ZN(
        n187) );
  AOI22D1BWP30P140LVT U222 ( .A1(n229), .A2(i_data_bus[83]), .B1(n228), .B2(
        i_data_bus[51]), .ZN(n186) );
  AOI22D1BWP30P140LVT U223 ( .A1(n231), .A2(i_data_bus[115]), .B1(n230), .B2(
        i_data_bus[147]), .ZN(n185) );
  ND3D1BWP30P140LVT U224 ( .A1(n187), .A2(n186), .A3(n185), .ZN(N388) );
  AOI22D1BWP30P140LVT U225 ( .A1(n2), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n188) );
  IOA21D1BWP30P140LVT U226 ( .A1(n226), .A2(i_data_bus[242]), .B(n188), .ZN(
        n189) );
  AOI21D1BWP30P140LVT U227 ( .A1(n217), .A2(i_data_bus[18]), .B(n189), .ZN(
        n192) );
  AOI22D1BWP30P140LVT U228 ( .A1(n229), .A2(i_data_bus[82]), .B1(n228), .B2(
        i_data_bus[50]), .ZN(n191) );
  AOI22D1BWP30P140LVT U229 ( .A1(n231), .A2(i_data_bus[114]), .B1(n230), .B2(
        i_data_bus[146]), .ZN(n190) );
  ND3D1BWP30P140LVT U230 ( .A1(n192), .A2(n191), .A3(n190), .ZN(N387) );
  AOI22D1BWP30P140LVT U231 ( .A1(n2), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n193) );
  IOA21D1BWP30P140LVT U232 ( .A1(n226), .A2(i_data_bus[245]), .B(n193), .ZN(
        n194) );
  AOI21D1BWP30P140LVT U233 ( .A1(n217), .A2(i_data_bus[21]), .B(n194), .ZN(
        n197) );
  AOI22D1BWP30P140LVT U234 ( .A1(n229), .A2(i_data_bus[85]), .B1(n228), .B2(
        i_data_bus[53]), .ZN(n196) );
  AOI22D1BWP30P140LVT U235 ( .A1(n231), .A2(i_data_bus[117]), .B1(n230), .B2(
        i_data_bus[149]), .ZN(n195) );
  ND3D1BWP30P140LVT U236 ( .A1(n197), .A2(n196), .A3(n195), .ZN(N390) );
  INVD1BWP30P140LVT U237 ( .I(i_data_bus[208]), .ZN(n198) );
  MAOI22D1BWP30P140LVT U238 ( .A1(n1), .A2(i_data_bus[176]), .B1(n199), .B2(
        n198), .ZN(n200) );
  IOA21D1BWP30P140LVT U239 ( .A1(n226), .A2(i_data_bus[240]), .B(n200), .ZN(
        n201) );
  AOI21D1BWP30P140LVT U240 ( .A1(n217), .A2(i_data_bus[16]), .B(n201), .ZN(
        n204) );
  AOI22D1BWP30P140LVT U241 ( .A1(n229), .A2(i_data_bus[80]), .B1(n228), .B2(
        i_data_bus[48]), .ZN(n203) );
  AOI22D1BWP30P140LVT U242 ( .A1(n231), .A2(i_data_bus[112]), .B1(n230), .B2(
        i_data_bus[144]), .ZN(n202) );
  ND3D1BWP30P140LVT U243 ( .A1(n204), .A2(n203), .A3(n202), .ZN(N385) );
  AOI22D1BWP30P140LVT U244 ( .A1(n2), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n205) );
  IOA21D1BWP30P140LVT U245 ( .A1(n226), .A2(i_data_bus[241]), .B(n205), .ZN(
        n206) );
  AOI21D1BWP30P140LVT U246 ( .A1(n217), .A2(i_data_bus[17]), .B(n206), .ZN(
        n209) );
  AOI22D1BWP30P140LVT U247 ( .A1(n229), .A2(i_data_bus[81]), .B1(n228), .B2(
        i_data_bus[49]), .ZN(n208) );
  AOI22D1BWP30P140LVT U248 ( .A1(n231), .A2(i_data_bus[113]), .B1(n230), .B2(
        i_data_bus[145]), .ZN(n207) );
  ND3D1BWP30P140LVT U249 ( .A1(n209), .A2(n208), .A3(n207), .ZN(N386) );
  AOI22D1BWP30P140LVT U250 ( .A1(n2), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n210) );
  IOA21D1BWP30P140LVT U251 ( .A1(n226), .A2(i_data_bus[247]), .B(n210), .ZN(
        n211) );
  AOI21D1BWP30P140LVT U252 ( .A1(n217), .A2(i_data_bus[23]), .B(n211), .ZN(
        n214) );
  AOI22D1BWP30P140LVT U253 ( .A1(n229), .A2(i_data_bus[87]), .B1(n228), .B2(
        i_data_bus[55]), .ZN(n213) );
  AOI22D1BWP30P140LVT U254 ( .A1(n231), .A2(i_data_bus[119]), .B1(n230), .B2(
        i_data_bus[151]), .ZN(n212) );
  ND3D1BWP30P140LVT U255 ( .A1(n214), .A2(n213), .A3(n212), .ZN(N392) );
  AOI22D1BWP30P140LVT U256 ( .A1(n2), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n215) );
  IOA21D1BWP30P140LVT U257 ( .A1(n226), .A2(i_data_bus[239]), .B(n215), .ZN(
        n216) );
  AOI21D1BWP30P140LVT U258 ( .A1(n217), .A2(i_data_bus[15]), .B(n216), .ZN(
        n224) );
  INVD1BWP30P140LVT U259 ( .I(i_data_bus[79]), .ZN(n220) );
  INVD1BWP30P140LVT U260 ( .I(i_data_bus[47]), .ZN(n218) );
  OA22D1BWP30P140LVT U261 ( .A1(n221), .A2(n220), .B1(n219), .B2(n218), .Z(
        n223) );
  AOI22D1BWP30P140LVT U262 ( .A1(n231), .A2(i_data_bus[111]), .B1(n230), .B2(
        i_data_bus[143]), .ZN(n222) );
  ND3D1BWP30P140LVT U263 ( .A1(n224), .A2(n223), .A3(n222), .ZN(N384) );
  AOI22D1BWP30P140LVT U264 ( .A1(n2), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n225) );
  IOA21D1BWP30P140LVT U265 ( .A1(n226), .A2(i_data_bus[248]), .B(n225), .ZN(
        n227) );
  AOI21D1BWP30P140LVT U266 ( .A1(n217), .A2(i_data_bus[24]), .B(n227), .ZN(
        n234) );
  AOI22D1BWP30P140LVT U267 ( .A1(n229), .A2(i_data_bus[88]), .B1(n228), .B2(
        i_data_bus[56]), .ZN(n233) );
  AOI22D1BWP30P140LVT U268 ( .A1(n231), .A2(i_data_bus[120]), .B1(n230), .B2(
        i_data_bus[152]), .ZN(n232) );
  ND3D1BWP30P140LVT U269 ( .A1(n234), .A2(n233), .A3(n232), .ZN(N393) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_4 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n46), .ZN(n231) );
  INVD2BWP30P140LVT U4 ( .I(n228), .ZN(n221) );
  INVD4BWP30P140LVT U5 ( .I(n65), .ZN(n4) );
  INVD4BWP30P140LVT U6 ( .I(n6), .ZN(n20) );
  BUFFD2BWP30P140LVT U7 ( .I(n51), .Z(n65) );
  INVD6BWP30P140LVT U8 ( .I(n113), .ZN(n3) );
  INVD2BWP30P140LVT U9 ( .I(n27), .ZN(n113) );
  NR2D1BWP30P140LVT U10 ( .A1(n11), .A2(n28), .ZN(n45) );
  NR2D1BWP30P140LVT U11 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n29) );
  INR4D1BWP30P140LVT U12 ( .A1(i_valid[6]), .B1(i_cmd[5]), .B2(i_cmd[7]), .B3(
        n21), .ZN(n22) );
  INR4D1BWP30P140LVT U13 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n24), .ZN(n26) );
  ND2OPTIBD1BWP30P140LVT U14 ( .A1(n45), .A2(n44), .ZN(n46) );
  INVD1BWP30P140LVT U15 ( .I(n36), .ZN(n228) );
  INVD2BWP30P140LVT U16 ( .I(n230), .ZN(n1) );
  INVD4BWP30P140LVT U17 ( .I(n188), .ZN(n2) );
  ND2OPTIBD2BWP30P140LVT U18 ( .A1(n10), .A2(n9), .ZN(n28) );
  INR2D1BWP30P140LVT U19 ( .A1(i_en), .B1(rst), .ZN(n8) );
  INR2D1BWP30P140LVT U20 ( .A1(n41), .B1(n35), .ZN(n36) );
  ND2D1BWP30P140LVT U21 ( .A1(n17), .A2(n16), .ZN(n18) );
  IND3D1BWP30P140LVT U22 ( .A1(n12), .B1(i_cmd[0]), .B2(n45), .ZN(n51) );
  INR2D2BWP30P140LVT U23 ( .A1(n29), .B1(n28), .ZN(n41) );
  OR2D1BWP30P140LVT U24 ( .A1(n33), .A2(i_cmd[1]), .Z(n11) );
  INVD2BWP30P140LVT U25 ( .I(n228), .ZN(n134) );
  AOI21D1BWP30P140LVT U26 ( .A1(n4), .A2(i_data_bus[14]), .B(n107), .ZN(n111)
         );
  AOI21D1BWP30P140LVT U27 ( .A1(n4), .A2(i_data_bus[18]), .B(n200), .ZN(n203)
         );
  OR2D2BWP30P140LVT U28 ( .A1(n5), .A2(n25), .Z(n6) );
  INVD1BWP30P140LVT U29 ( .I(n19), .ZN(n5) );
  INVD1BWP30P140LVT U30 ( .I(n32), .ZN(n230) );
  INVD1BWP30P140LVT U31 ( .I(n42), .ZN(n108) );
  INR2D1BWP30P140LVT U32 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n7) );
  INVD1BWP30P140LVT U33 ( .I(n7), .ZN(n12) );
  OR2D1BWP30P140LVT U34 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n33) );
  NR2OPTPAD1BWP30P140LVT U35 ( .A1(i_cmd[7]), .A2(i_cmd[6]), .ZN(n10) );
  INR2D2BWP30P140LVT U36 ( .A1(n8), .B1(i_cmd[5]), .ZN(n9) );
  ND2D1BWP30P140LVT U37 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n13) );
  NR3D0P7BWP30P140LVT U38 ( .A1(n13), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n19)
         );
  INVD1BWP30P140LVT U39 ( .I(i_cmd[2]), .ZN(n14) );
  INVD2BWP30P140LVT U40 ( .I(i_cmd[1]), .ZN(n30) );
  ND2OPTIBD2BWP30P140LVT U41 ( .A1(n14), .A2(n30), .ZN(n37) );
  NR2D1BWP30P140LVT U42 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n17) );
  INR2D1BWP30P140LVT U43 ( .A1(i_en), .B1(rst), .ZN(n15) );
  INR2D1BWP30P140LVT U44 ( .A1(n15), .B1(i_cmd[3]), .ZN(n16) );
  OR2D4BWP30P140LVT U45 ( .A1(n37), .A2(n18), .Z(n25) );
  INVD1BWP30P140LVT U46 ( .I(i_cmd[6]), .ZN(n21) );
  INR2D2BWP30P140LVT U47 ( .A1(n22), .B1(n25), .ZN(n23) );
  INVD3BWP30P140LVT U48 ( .I(n23), .ZN(n188) );
  INVD1BWP30P140LVT U49 ( .I(i_cmd[5]), .ZN(n24) );
  INR2D2BWP30P140LVT U50 ( .A1(n26), .B1(n25), .ZN(n27) );
  NR4D0BWP30P140LVT U51 ( .A1(n4), .A2(n20), .A3(n2), .A4(n3), .ZN(n49) );
  INVD1BWP30P140LVT U52 ( .I(i_cmd[3]), .ZN(n38) );
  ND4D1BWP30P140LVT U53 ( .A1(n30), .A2(n38), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n31) );
  INR2D1BWP30P140LVT U54 ( .A1(n41), .B1(n31), .ZN(n32) );
  INVD1BWP30P140LVT U55 ( .I(n33), .ZN(n34) );
  ND3D1BWP30P140LVT U56 ( .A1(n34), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n35)
         );
  NR2D1BWP30P140LVT U57 ( .A1(n1), .A2(n221), .ZN(n48) );
  INVD1BWP30P140LVT U58 ( .I(n37), .ZN(n39) );
  ND3D1BWP30P140LVT U59 ( .A1(n39), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n40)
         );
  INR2D1BWP30P140LVT U60 ( .A1(n41), .B1(n40), .ZN(n42) );
  IND3D1BWP30P140LVT U61 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n43) );
  INVD1BWP30P140LVT U62 ( .I(n43), .ZN(n44) );
  NR2D1BWP30P140LVT U63 ( .A1(n42), .A2(n231), .ZN(n47) );
  ND3D1BWP30P140LVT U64 ( .A1(n49), .A2(n48), .A3(n47), .ZN(N402) );
  INVD1BWP30P140LVT U65 ( .I(n20), .ZN(n56) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[224]), .ZN(n55) );
  INVD1BWP30P140LVT U67 ( .I(i_data_bus[192]), .ZN(n50) );
  MAOI22D1BWP30P140LVT U68 ( .A1(n3), .A2(i_data_bus[160]), .B1(n188), .B2(n50), .ZN(n54) );
  INR2D1BWP30P140LVT U69 ( .A1(i_data_bus[0]), .B1(n51), .ZN(n52) );
  INVD1BWP30P140LVT U70 ( .I(n52), .ZN(n53) );
  OA211D1BWP30P140LVT U71 ( .A1(n56), .A2(n55), .B(n54), .C(n53), .Z(n59) );
  AOI22D1BWP30P140LVT U72 ( .A1(n1), .A2(i_data_bus[64]), .B1(n134), .B2(
        i_data_bus[32]), .ZN(n58) );
  INVD2BWP30P140LVT U73 ( .I(n108), .ZN(n135) );
  AOI22D1BWP30P140LVT U74 ( .A1(n135), .A2(i_data_bus[96]), .B1(n231), .B2(
        i_data_bus[128]), .ZN(n57) );
  ND3D1BWP30P140LVT U75 ( .A1(n59), .A2(n58), .A3(n57), .ZN(N369) );
  AOI22D1BWP30P140LVT U76 ( .A1(n2), .A2(i_data_bus[204]), .B1(n3), .B2(
        i_data_bus[172]), .ZN(n60) );
  IOA21D1BWP30P140LVT U77 ( .A1(n20), .A2(i_data_bus[236]), .B(n60), .ZN(n61)
         );
  AOI21D1BWP30P140LVT U78 ( .A1(n4), .A2(i_data_bus[12]), .B(n61), .ZN(n64) );
  AOI22D1BWP30P140LVT U79 ( .A1(n1), .A2(i_data_bus[76]), .B1(n134), .B2(
        i_data_bus[44]), .ZN(n63) );
  AOI22D1BWP30P140LVT U80 ( .A1(n135), .A2(i_data_bus[108]), .B1(n231), .B2(
        i_data_bus[140]), .ZN(n62) );
  ND3D1BWP30P140LVT U81 ( .A1(n64), .A2(n63), .A3(n62), .ZN(N381) );
  AOI22D1BWP30P140LVT U82 ( .A1(n2), .A2(i_data_bus[203]), .B1(n3), .B2(
        i_data_bus[171]), .ZN(n66) );
  IOA21D1BWP30P140LVT U83 ( .A1(n20), .A2(i_data_bus[235]), .B(n66), .ZN(n67)
         );
  AOI21D1BWP30P140LVT U84 ( .A1(n4), .A2(i_data_bus[11]), .B(n67), .ZN(n70) );
  AOI22D1BWP30P140LVT U85 ( .A1(n1), .A2(i_data_bus[75]), .B1(n134), .B2(
        i_data_bus[43]), .ZN(n69) );
  AOI22D1BWP30P140LVT U86 ( .A1(n135), .A2(i_data_bus[107]), .B1(n231), .B2(
        i_data_bus[139]), .ZN(n68) );
  ND3D1BWP30P140LVT U87 ( .A1(n70), .A2(n69), .A3(n68), .ZN(N380) );
  AOI22D1BWP30P140LVT U88 ( .A1(n2), .A2(i_data_bus[202]), .B1(n3), .B2(
        i_data_bus[170]), .ZN(n71) );
  IOA21D1BWP30P140LVT U89 ( .A1(n20), .A2(i_data_bus[234]), .B(n71), .ZN(n72)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n4), .A2(i_data_bus[10]), .B(n72), .ZN(n75) );
  AOI22D1BWP30P140LVT U91 ( .A1(n1), .A2(i_data_bus[74]), .B1(n134), .B2(
        i_data_bus[42]), .ZN(n74) );
  AOI22D1BWP30P140LVT U92 ( .A1(n135), .A2(i_data_bus[106]), .B1(n231), .B2(
        i_data_bus[138]), .ZN(n73) );
  ND3D1BWP30P140LVT U93 ( .A1(n75), .A2(n74), .A3(n73), .ZN(N379) );
  AOI22D1BWP30P140LVT U94 ( .A1(n2), .A2(i_data_bus[201]), .B1(n3), .B2(
        i_data_bus[169]), .ZN(n76) );
  IOA21D1BWP30P140LVT U95 ( .A1(n20), .A2(i_data_bus[233]), .B(n76), .ZN(n77)
         );
  AOI21D1BWP30P140LVT U96 ( .A1(n4), .A2(i_data_bus[9]), .B(n77), .ZN(n80) );
  AOI22D1BWP30P140LVT U97 ( .A1(n1), .A2(i_data_bus[73]), .B1(n134), .B2(
        i_data_bus[41]), .ZN(n79) );
  AOI22D1BWP30P140LVT U98 ( .A1(n135), .A2(i_data_bus[105]), .B1(n231), .B2(
        i_data_bus[137]), .ZN(n78) );
  ND3D1BWP30P140LVT U99 ( .A1(n80), .A2(n79), .A3(n78), .ZN(N378) );
  AOI22D1BWP30P140LVT U100 ( .A1(n2), .A2(i_data_bus[200]), .B1(n3), .B2(
        i_data_bus[168]), .ZN(n81) );
  IOA21D1BWP30P140LVT U101 ( .A1(n20), .A2(i_data_bus[232]), .B(n81), .ZN(n82)
         );
  AOI21D1BWP30P140LVT U102 ( .A1(n4), .A2(i_data_bus[8]), .B(n82), .ZN(n85) );
  AOI22D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[72]), .B1(n134), .B2(
        i_data_bus[40]), .ZN(n84) );
  AOI22D1BWP30P140LVT U104 ( .A1(n135), .A2(i_data_bus[104]), .B1(n231), .B2(
        i_data_bus[136]), .ZN(n83) );
  ND3D1BWP30P140LVT U105 ( .A1(n85), .A2(n84), .A3(n83), .ZN(N377) );
  AOI22D1BWP30P140LVT U106 ( .A1(n2), .A2(i_data_bus[199]), .B1(n3), .B2(
        i_data_bus[167]), .ZN(n86) );
  IOA21D1BWP30P140LVT U107 ( .A1(n20), .A2(i_data_bus[231]), .B(n86), .ZN(n87)
         );
  AOI21D1BWP30P140LVT U108 ( .A1(n4), .A2(i_data_bus[7]), .B(n87), .ZN(n90) );
  AOI22D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[71]), .B1(n134), .B2(
        i_data_bus[39]), .ZN(n89) );
  AOI22D1BWP30P140LVT U110 ( .A1(n135), .A2(i_data_bus[103]), .B1(n231), .B2(
        i_data_bus[135]), .ZN(n88) );
  ND3D1BWP30P140LVT U111 ( .A1(n90), .A2(n89), .A3(n88), .ZN(N376) );
  AOI22D1BWP30P140LVT U112 ( .A1(n2), .A2(i_data_bus[198]), .B1(n3), .B2(
        i_data_bus[166]), .ZN(n91) );
  IOA21D1BWP30P140LVT U113 ( .A1(n20), .A2(i_data_bus[230]), .B(n91), .ZN(n92)
         );
  AOI21D1BWP30P140LVT U114 ( .A1(n4), .A2(i_data_bus[6]), .B(n92), .ZN(n95) );
  AOI22D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[70]), .B1(n134), .B2(
        i_data_bus[38]), .ZN(n94) );
  AOI22D1BWP30P140LVT U116 ( .A1(n135), .A2(i_data_bus[102]), .B1(n231), .B2(
        i_data_bus[134]), .ZN(n93) );
  ND3D1BWP30P140LVT U117 ( .A1(n95), .A2(n94), .A3(n93), .ZN(N375) );
  AOI22D1BWP30P140LVT U118 ( .A1(n2), .A2(i_data_bus[197]), .B1(n3), .B2(
        i_data_bus[165]), .ZN(n96) );
  IOA21D1BWP30P140LVT U119 ( .A1(n20), .A2(i_data_bus[229]), .B(n96), .ZN(n97)
         );
  AOI21D1BWP30P140LVT U120 ( .A1(n4), .A2(i_data_bus[5]), .B(n97), .ZN(n100)
         );
  AOI22D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[69]), .B1(n134), .B2(
        i_data_bus[37]), .ZN(n99) );
  AOI22D1BWP30P140LVT U122 ( .A1(n135), .A2(i_data_bus[101]), .B1(n231), .B2(
        i_data_bus[133]), .ZN(n98) );
  ND3D1BWP30P140LVT U123 ( .A1(n100), .A2(n99), .A3(n98), .ZN(N374) );
  AOI22D1BWP30P140LVT U124 ( .A1(n2), .A2(i_data_bus[196]), .B1(n3), .B2(
        i_data_bus[164]), .ZN(n101) );
  IOA21D1BWP30P140LVT U125 ( .A1(n20), .A2(i_data_bus[228]), .B(n101), .ZN(
        n102) );
  AOI21D1BWP30P140LVT U126 ( .A1(n4), .A2(i_data_bus[4]), .B(n102), .ZN(n105)
         );
  AOI22D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[68]), .B1(n134), .B2(
        i_data_bus[36]), .ZN(n104) );
  AOI22D1BWP30P140LVT U128 ( .A1(n135), .A2(i_data_bus[100]), .B1(n231), .B2(
        i_data_bus[132]), .ZN(n103) );
  ND3D1BWP30P140LVT U129 ( .A1(n105), .A2(n104), .A3(n103), .ZN(N373) );
  AOI22D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[206]), .B1(n3), .B2(
        i_data_bus[174]), .ZN(n106) );
  IOA21D1BWP30P140LVT U131 ( .A1(n20), .A2(i_data_bus[238]), .B(n106), .ZN(
        n107) );
  AOI22D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[78]), .B1(n221), .B2(
        i_data_bus[46]), .ZN(n110) );
  INVD2BWP30P140LVT U133 ( .I(n108), .ZN(n232) );
  AOI22D1BWP30P140LVT U134 ( .A1(n232), .A2(i_data_bus[110]), .B1(n231), .B2(
        i_data_bus[142]), .ZN(n109) );
  ND3D1BWP30P140LVT U135 ( .A1(n111), .A2(n110), .A3(n109), .ZN(N383) );
  INVD1BWP30P140LVT U136 ( .I(i_data_bus[173]), .ZN(n112) );
  MAOI22D1BWP30P140LVT U137 ( .A1(n2), .A2(i_data_bus[205]), .B1(n113), .B2(
        n112), .ZN(n114) );
  IOA21D1BWP30P140LVT U138 ( .A1(n20), .A2(i_data_bus[237]), .B(n114), .ZN(
        n115) );
  AOI21D1BWP30P140LVT U139 ( .A1(n4), .A2(i_data_bus[13]), .B(n115), .ZN(n118)
         );
  AOI22D1BWP30P140LVT U140 ( .A1(n1), .A2(i_data_bus[77]), .B1(n221), .B2(
        i_data_bus[45]), .ZN(n117) );
  AOI22D1BWP30P140LVT U141 ( .A1(n232), .A2(i_data_bus[109]), .B1(n231), .B2(
        i_data_bus[141]), .ZN(n116) );
  ND3D1BWP30P140LVT U142 ( .A1(n118), .A2(n117), .A3(n116), .ZN(N382) );
  INVD1BWP30P140LVT U143 ( .I(i_data_bus[193]), .ZN(n119) );
  MAOI22D1BWP30P140LVT U144 ( .A1(n3), .A2(i_data_bus[161]), .B1(n188), .B2(
        n119), .ZN(n120) );
  IOA21D1BWP30P140LVT U145 ( .A1(n20), .A2(i_data_bus[225]), .B(n120), .ZN(
        n121) );
  AOI21D1BWP30P140LVT U146 ( .A1(n4), .A2(i_data_bus[1]), .B(n121), .ZN(n124)
         );
  AOI22D1BWP30P140LVT U147 ( .A1(n1), .A2(i_data_bus[65]), .B1(n134), .B2(
        i_data_bus[33]), .ZN(n123) );
  AOI22D1BWP30P140LVT U148 ( .A1(n135), .A2(i_data_bus[97]), .B1(n231), .B2(
        i_data_bus[129]), .ZN(n122) );
  ND3D1BWP30P140LVT U149 ( .A1(n124), .A2(n123), .A3(n122), .ZN(N370) );
  INVD1BWP30P140LVT U150 ( .I(i_data_bus[194]), .ZN(n125) );
  MAOI22D1BWP30P140LVT U151 ( .A1(n3), .A2(i_data_bus[162]), .B1(n188), .B2(
        n125), .ZN(n126) );
  IOA21D1BWP30P140LVT U152 ( .A1(n20), .A2(i_data_bus[226]), .B(n126), .ZN(
        n127) );
  AOI21D1BWP30P140LVT U153 ( .A1(n4), .A2(i_data_bus[2]), .B(n127), .ZN(n130)
         );
  AOI22D1BWP30P140LVT U154 ( .A1(n1), .A2(i_data_bus[66]), .B1(n134), .B2(
        i_data_bus[34]), .ZN(n129) );
  AOI22D1BWP30P140LVT U155 ( .A1(n135), .A2(i_data_bus[98]), .B1(n231), .B2(
        i_data_bus[130]), .ZN(n128) );
  ND3D1BWP30P140LVT U156 ( .A1(n130), .A2(n129), .A3(n128), .ZN(N371) );
  INVD1BWP30P140LVT U157 ( .I(i_data_bus[195]), .ZN(n131) );
  MAOI22D1BWP30P140LVT U158 ( .A1(n3), .A2(i_data_bus[163]), .B1(n188), .B2(
        n131), .ZN(n132) );
  IOA21D1BWP30P140LVT U159 ( .A1(n20), .A2(i_data_bus[227]), .B(n132), .ZN(
        n133) );
  AOI21D1BWP30P140LVT U160 ( .A1(n4), .A2(i_data_bus[3]), .B(n133), .ZN(n138)
         );
  AOI22D1BWP30P140LVT U161 ( .A1(n1), .A2(i_data_bus[67]), .B1(n134), .B2(
        i_data_bus[35]), .ZN(n137) );
  AOI22D1BWP30P140LVT U162 ( .A1(n135), .A2(i_data_bus[99]), .B1(n231), .B2(
        i_data_bus[131]), .ZN(n136) );
  ND3D1BWP30P140LVT U163 ( .A1(n138), .A2(n137), .A3(n136), .ZN(N372) );
  INVD1BWP30P140LVT U164 ( .I(i_data_bus[223]), .ZN(n139) );
  MAOI22D1BWP30P140LVT U165 ( .A1(n3), .A2(i_data_bus[191]), .B1(n188), .B2(
        n139), .ZN(n140) );
  IOA21D1BWP30P140LVT U166 ( .A1(n20), .A2(i_data_bus[255]), .B(n140), .ZN(
        n141) );
  AOI21D1BWP30P140LVT U167 ( .A1(n4), .A2(i_data_bus[31]), .B(n141), .ZN(n144)
         );
  AOI22D1BWP30P140LVT U168 ( .A1(n1), .A2(i_data_bus[95]), .B1(n221), .B2(
        i_data_bus[63]), .ZN(n143) );
  AOI22D1BWP30P140LVT U169 ( .A1(n135), .A2(i_data_bus[127]), .B1(n231), .B2(
        i_data_bus[159]), .ZN(n142) );
  ND3D1BWP30P140LVT U170 ( .A1(n144), .A2(n143), .A3(n142), .ZN(N400) );
  AOI22D1BWP30P140LVT U171 ( .A1(n2), .A2(i_data_bus[217]), .B1(n3), .B2(
        i_data_bus[185]), .ZN(n145) );
  IOA21D1BWP30P140LVT U172 ( .A1(n20), .A2(i_data_bus[249]), .B(n145), .ZN(
        n146) );
  AOI21D1BWP30P140LVT U173 ( .A1(n4), .A2(i_data_bus[25]), .B(n146), .ZN(n149)
         );
  AOI22D1BWP30P140LVT U174 ( .A1(n1), .A2(i_data_bus[89]), .B1(n221), .B2(
        i_data_bus[57]), .ZN(n148) );
  AOI22D1BWP30P140LVT U175 ( .A1(n232), .A2(i_data_bus[121]), .B1(n231), .B2(
        i_data_bus[153]), .ZN(n147) );
  ND3D1BWP30P140LVT U176 ( .A1(n149), .A2(n148), .A3(n147), .ZN(N394) );
  AOI22D1BWP30P140LVT U177 ( .A1(n2), .A2(i_data_bus[219]), .B1(n3), .B2(
        i_data_bus[187]), .ZN(n150) );
  IOA21D1BWP30P140LVT U178 ( .A1(n20), .A2(i_data_bus[251]), .B(n150), .ZN(
        n151) );
  AOI21D1BWP30P140LVT U179 ( .A1(n4), .A2(i_data_bus[27]), .B(n151), .ZN(n154)
         );
  AOI22D1BWP30P140LVT U180 ( .A1(n1), .A2(i_data_bus[91]), .B1(n221), .B2(
        i_data_bus[59]), .ZN(n153) );
  AOI22D1BWP30P140LVT U181 ( .A1(n232), .A2(i_data_bus[123]), .B1(n231), .B2(
        i_data_bus[155]), .ZN(n152) );
  ND3D1BWP30P140LVT U182 ( .A1(n154), .A2(n153), .A3(n152), .ZN(N396) );
  AOI22D1BWP30P140LVT U183 ( .A1(n2), .A2(i_data_bus[220]), .B1(n3), .B2(
        i_data_bus[188]), .ZN(n155) );
  IOA21D1BWP30P140LVT U184 ( .A1(n20), .A2(i_data_bus[252]), .B(n155), .ZN(
        n156) );
  AOI21D1BWP30P140LVT U185 ( .A1(n4), .A2(i_data_bus[28]), .B(n156), .ZN(n159)
         );
  AOI22D1BWP30P140LVT U186 ( .A1(n1), .A2(i_data_bus[92]), .B1(n221), .B2(
        i_data_bus[60]), .ZN(n158) );
  AOI22D1BWP30P140LVT U187 ( .A1(n135), .A2(i_data_bus[124]), .B1(n231), .B2(
        i_data_bus[156]), .ZN(n157) );
  ND3D1BWP30P140LVT U188 ( .A1(n159), .A2(n158), .A3(n157), .ZN(N397) );
  INVD1BWP30P140LVT U189 ( .I(i_data_bus[221]), .ZN(n160) );
  MAOI22D1BWP30P140LVT U190 ( .A1(n3), .A2(i_data_bus[189]), .B1(n188), .B2(
        n160), .ZN(n161) );
  IOA21D1BWP30P140LVT U191 ( .A1(n20), .A2(i_data_bus[253]), .B(n161), .ZN(
        n162) );
  AOI21D1BWP30P140LVT U192 ( .A1(n4), .A2(i_data_bus[29]), .B(n162), .ZN(n165)
         );
  AOI22D1BWP30P140LVT U193 ( .A1(n1), .A2(i_data_bus[93]), .B1(n221), .B2(
        i_data_bus[61]), .ZN(n164) );
  AOI22D1BWP30P140LVT U194 ( .A1(n232), .A2(i_data_bus[125]), .B1(n231), .B2(
        i_data_bus[157]), .ZN(n163) );
  ND3D1BWP30P140LVT U195 ( .A1(n165), .A2(n164), .A3(n163), .ZN(N398) );
  INVD1BWP30P140LVT U196 ( .I(i_data_bus[222]), .ZN(n166) );
  MAOI22D1BWP30P140LVT U197 ( .A1(n3), .A2(i_data_bus[190]), .B1(n188), .B2(
        n166), .ZN(n167) );
  IOA21D1BWP30P140LVT U198 ( .A1(n20), .A2(i_data_bus[254]), .B(n167), .ZN(
        n168) );
  AOI21D1BWP30P140LVT U199 ( .A1(n4), .A2(i_data_bus[30]), .B(n168), .ZN(n171)
         );
  AOI22D1BWP30P140LVT U200 ( .A1(n1), .A2(i_data_bus[94]), .B1(n221), .B2(
        i_data_bus[62]), .ZN(n170) );
  AOI22D1BWP30P140LVT U201 ( .A1(n135), .A2(i_data_bus[126]), .B1(n231), .B2(
        i_data_bus[158]), .ZN(n169) );
  ND3D1BWP30P140LVT U202 ( .A1(n171), .A2(n170), .A3(n169), .ZN(N399) );
  AOI22D1BWP30P140LVT U203 ( .A1(n2), .A2(i_data_bus[218]), .B1(n3), .B2(
        i_data_bus[186]), .ZN(n172) );
  IOA21D1BWP30P140LVT U204 ( .A1(n20), .A2(i_data_bus[250]), .B(n172), .ZN(
        n173) );
  AOI21D1BWP30P140LVT U205 ( .A1(n4), .A2(i_data_bus[26]), .B(n173), .ZN(n176)
         );
  AOI22D1BWP30P140LVT U206 ( .A1(n1), .A2(i_data_bus[90]), .B1(n221), .B2(
        i_data_bus[58]), .ZN(n175) );
  AOI22D1BWP30P140LVT U207 ( .A1(n232), .A2(i_data_bus[122]), .B1(n231), .B2(
        i_data_bus[154]), .ZN(n174) );
  ND3D1BWP30P140LVT U208 ( .A1(n176), .A2(n175), .A3(n174), .ZN(N395) );
  AOI22D1BWP30P140LVT U209 ( .A1(n2), .A2(i_data_bus[216]), .B1(n3), .B2(
        i_data_bus[184]), .ZN(n177) );
  IOA21D1BWP30P140LVT U210 ( .A1(n20), .A2(i_data_bus[248]), .B(n177), .ZN(
        n178) );
  AOI21D1BWP30P140LVT U211 ( .A1(n4), .A2(i_data_bus[24]), .B(n178), .ZN(n181)
         );
  AOI22D1BWP30P140LVT U212 ( .A1(n1), .A2(i_data_bus[88]), .B1(n221), .B2(
        i_data_bus[56]), .ZN(n180) );
  AOI22D1BWP30P140LVT U213 ( .A1(n232), .A2(i_data_bus[120]), .B1(n231), .B2(
        i_data_bus[152]), .ZN(n179) );
  ND3D1BWP30P140LVT U214 ( .A1(n181), .A2(n180), .A3(n179), .ZN(N393) );
  AOI22D1BWP30P140LVT U215 ( .A1(n2), .A2(i_data_bus[209]), .B1(n3), .B2(
        i_data_bus[177]), .ZN(n182) );
  IOA21D1BWP30P140LVT U216 ( .A1(n20), .A2(i_data_bus[241]), .B(n182), .ZN(
        n183) );
  AOI21D1BWP30P140LVT U217 ( .A1(n4), .A2(i_data_bus[17]), .B(n183), .ZN(n186)
         );
  AOI22D1BWP30P140LVT U218 ( .A1(n1), .A2(i_data_bus[81]), .B1(n221), .B2(
        i_data_bus[49]), .ZN(n185) );
  AOI22D1BWP30P140LVT U219 ( .A1(n232), .A2(i_data_bus[113]), .B1(n231), .B2(
        i_data_bus[145]), .ZN(n184) );
  ND3D1BWP30P140LVT U220 ( .A1(n186), .A2(n185), .A3(n184), .ZN(N386) );
  INVD1BWP30P140LVT U221 ( .I(i_data_bus[208]), .ZN(n187) );
  MAOI22D1BWP30P140LVT U222 ( .A1(n3), .A2(i_data_bus[176]), .B1(n188), .B2(
        n187), .ZN(n189) );
  IOA21D1BWP30P140LVT U223 ( .A1(n20), .A2(i_data_bus[240]), .B(n189), .ZN(
        n190) );
  AOI21D1BWP30P140LVT U224 ( .A1(n4), .A2(i_data_bus[16]), .B(n190), .ZN(n193)
         );
  AOI22D1BWP30P140LVT U225 ( .A1(n1), .A2(i_data_bus[80]), .B1(n221), .B2(
        i_data_bus[48]), .ZN(n192) );
  AOI22D1BWP30P140LVT U226 ( .A1(n232), .A2(i_data_bus[112]), .B1(n231), .B2(
        i_data_bus[144]), .ZN(n191) );
  ND3D1BWP30P140LVT U227 ( .A1(n193), .A2(n192), .A3(n191), .ZN(N385) );
  AOI22D1BWP30P140LVT U228 ( .A1(n2), .A2(i_data_bus[212]), .B1(n3), .B2(
        i_data_bus[180]), .ZN(n194) );
  IOA21D1BWP30P140LVT U229 ( .A1(n20), .A2(i_data_bus[244]), .B(n194), .ZN(
        n195) );
  AOI21D1BWP30P140LVT U230 ( .A1(n4), .A2(i_data_bus[20]), .B(n195), .ZN(n198)
         );
  AOI22D1BWP30P140LVT U231 ( .A1(n1), .A2(i_data_bus[84]), .B1(n221), .B2(
        i_data_bus[52]), .ZN(n197) );
  AOI22D1BWP30P140LVT U232 ( .A1(n232), .A2(i_data_bus[116]), .B1(n231), .B2(
        i_data_bus[148]), .ZN(n196) );
  ND3D1BWP30P140LVT U233 ( .A1(n198), .A2(n197), .A3(n196), .ZN(N389) );
  AOI22D1BWP30P140LVT U234 ( .A1(n2), .A2(i_data_bus[210]), .B1(n3), .B2(
        i_data_bus[178]), .ZN(n199) );
  IOA21D1BWP30P140LVT U235 ( .A1(n20), .A2(i_data_bus[242]), .B(n199), .ZN(
        n200) );
  AOI22D1BWP30P140LVT U236 ( .A1(n1), .A2(i_data_bus[82]), .B1(n221), .B2(
        i_data_bus[50]), .ZN(n202) );
  AOI22D1BWP30P140LVT U237 ( .A1(n232), .A2(i_data_bus[114]), .B1(n231), .B2(
        i_data_bus[146]), .ZN(n201) );
  ND3D1BWP30P140LVT U238 ( .A1(n203), .A2(n202), .A3(n201), .ZN(N387) );
  AOI22D1BWP30P140LVT U239 ( .A1(n2), .A2(i_data_bus[211]), .B1(n3), .B2(
        i_data_bus[179]), .ZN(n204) );
  IOA21D1BWP30P140LVT U240 ( .A1(n20), .A2(i_data_bus[243]), .B(n204), .ZN(
        n205) );
  AOI21D1BWP30P140LVT U241 ( .A1(n4), .A2(i_data_bus[19]), .B(n205), .ZN(n208)
         );
  AOI22D1BWP30P140LVT U242 ( .A1(n1), .A2(i_data_bus[83]), .B1(n221), .B2(
        i_data_bus[51]), .ZN(n207) );
  AOI22D1BWP30P140LVT U243 ( .A1(n232), .A2(i_data_bus[115]), .B1(n231), .B2(
        i_data_bus[147]), .ZN(n206) );
  ND3D1BWP30P140LVT U244 ( .A1(n208), .A2(n207), .A3(n206), .ZN(N388) );
  AOI22D1BWP30P140LVT U245 ( .A1(n2), .A2(i_data_bus[214]), .B1(n3), .B2(
        i_data_bus[182]), .ZN(n209) );
  IOA21D1BWP30P140LVT U246 ( .A1(n20), .A2(i_data_bus[246]), .B(n209), .ZN(
        n210) );
  AOI21D1BWP30P140LVT U247 ( .A1(n4), .A2(i_data_bus[22]), .B(n210), .ZN(n213)
         );
  AOI22D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[86]), .B1(n221), .B2(
        i_data_bus[54]), .ZN(n212) );
  AOI22D1BWP30P140LVT U249 ( .A1(n232), .A2(i_data_bus[118]), .B1(n231), .B2(
        i_data_bus[150]), .ZN(n211) );
  ND3D1BWP30P140LVT U250 ( .A1(n213), .A2(n212), .A3(n211), .ZN(N391) );
  AOI22D1BWP30P140LVT U251 ( .A1(n2), .A2(i_data_bus[215]), .B1(n3), .B2(
        i_data_bus[183]), .ZN(n214) );
  IOA21D1BWP30P140LVT U252 ( .A1(n20), .A2(i_data_bus[247]), .B(n214), .ZN(
        n215) );
  AOI21D1BWP30P140LVT U253 ( .A1(n4), .A2(i_data_bus[23]), .B(n215), .ZN(n218)
         );
  AOI22D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[87]), .B1(n221), .B2(
        i_data_bus[55]), .ZN(n217) );
  AOI22D1BWP30P140LVT U255 ( .A1(n232), .A2(i_data_bus[119]), .B1(n231), .B2(
        i_data_bus[151]), .ZN(n216) );
  ND3D1BWP30P140LVT U256 ( .A1(n218), .A2(n217), .A3(n216), .ZN(N392) );
  AOI22D1BWP30P140LVT U257 ( .A1(n2), .A2(i_data_bus[213]), .B1(n3), .B2(
        i_data_bus[181]), .ZN(n219) );
  IOA21D1BWP30P140LVT U258 ( .A1(n20), .A2(i_data_bus[245]), .B(n219), .ZN(
        n220) );
  AOI21D1BWP30P140LVT U259 ( .A1(n4), .A2(i_data_bus[21]), .B(n220), .ZN(n224)
         );
  AOI22D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[85]), .B1(n221), .B2(
        i_data_bus[53]), .ZN(n223) );
  AOI22D1BWP30P140LVT U261 ( .A1(n232), .A2(i_data_bus[117]), .B1(n231), .B2(
        i_data_bus[149]), .ZN(n222) );
  ND3D1BWP30P140LVT U262 ( .A1(n224), .A2(n223), .A3(n222), .ZN(N390) );
  AOI22D1BWP30P140LVT U263 ( .A1(n2), .A2(i_data_bus[207]), .B1(n3), .B2(
        i_data_bus[175]), .ZN(n225) );
  IOA21D1BWP30P140LVT U264 ( .A1(n20), .A2(i_data_bus[239]), .B(n225), .ZN(
        n226) );
  AOI21D1BWP30P140LVT U265 ( .A1(n4), .A2(i_data_bus[15]), .B(n226), .ZN(n235)
         );
  INVD1BWP30P140LVT U266 ( .I(i_data_bus[79]), .ZN(n229) );
  INVD1BWP30P140LVT U267 ( .I(i_data_bus[47]), .ZN(n227) );
  OA22D1BWP30P140LVT U268 ( .A1(n230), .A2(n229), .B1(n228), .B2(n227), .Z(
        n234) );
  AOI22D1BWP30P140LVT U269 ( .A1(n232), .A2(i_data_bus[111]), .B1(n231), .B2(
        i_data_bus[143]), .ZN(n233) );
  ND3D1BWP30P140LVT U270 ( .A1(n235), .A2(n234), .A3(n233), .ZN(N384) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_5 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD2BWP30P140LVT U3 ( .I(n220), .ZN(n211) );
  INVD2BWP30P140LVT U4 ( .I(n56), .ZN(n231) );
  INVD6BWP30P140LVT U5 ( .I(n226), .ZN(n2) );
  INVD1BWP30P140LVT U6 ( .I(n38), .ZN(n39) );
  NR2OPTPAD1BWP30P140LVT U7 ( .A1(n11), .A2(n32), .ZN(n45) );
  CKND2D3BWP30P140LVT U8 ( .A1(n10), .A2(n9), .ZN(n32) );
  NR2D1BWP30P140LVT U9 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n33) );
  NR3OPTPAD2BWP30P140LVT U10 ( .A1(i_cmd[6]), .A2(i_cmd[5]), .A3(i_cmd[7]), 
        .ZN(n10) );
  MAOI22D1BWP30P140LVT U11 ( .A1(n2), .A2(i_data_bus[205]), .B1(n111), .B2(
        n110), .ZN(n112) );
  ND2OPTIBD1BWP30P140LVT U12 ( .A1(n46), .A2(n45), .ZN(n56) );
  ND2OPTIBD2BWP30P140LVT U13 ( .A1(n39), .A2(n43), .ZN(n218) );
  INVD8BWP30P140LVT U14 ( .I(n111), .ZN(n1) );
  INVD2BWP30P140LVT U15 ( .I(n51), .ZN(n3) );
  INR2D1BWP30P140LVT U16 ( .A1(n15), .B1(i_cmd[3]), .ZN(n16) );
  INVD3BWP30P140LVT U17 ( .I(n26), .ZN(n226) );
  INVD1BWP30P140LVT U18 ( .I(i_valid[5]), .ZN(n27) );
  ND2OPTIBD1BWP30P140LVT U19 ( .A1(n22), .A2(i_valid[6]), .ZN(n24) );
  NR2D1BWP30P140LVT U20 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .ZN(n22) );
  INVD1BWP30P140LVT U21 ( .I(n44), .ZN(n46) );
  INVD1BWP30P140LVT U22 ( .I(n5), .ZN(n51) );
  NR4D0BWP30P140LVT U23 ( .A1(n11), .A2(n32), .A3(n12), .A4(n4), .ZN(n5) );
  INVD1BWP30P140LVT U24 ( .I(i_cmd[0]), .ZN(n4) );
  INR2D1BWP30P140LVT U25 ( .A1(n43), .B1(n35), .ZN(n172) );
  INVD1BWP30P140LVT U26 ( .I(n172), .ZN(n220) );
  INVD2BWP30P140LVT U27 ( .I(n220), .ZN(n230) );
  INR2D1BWP30P140LVT U28 ( .A1(i_en), .B1(rst), .ZN(n9) );
  NR4D0BWP30P140LVT U29 ( .A1(n28), .A2(n27), .A3(i_cmd[6]), .A4(i_cmd[7]), 
        .ZN(n30) );
  INVD1BWP30P140LVT U30 ( .I(i_cmd[5]), .ZN(n28) );
  NR2D1BWP30P140LVT U31 ( .A1(n24), .A2(n23), .ZN(n25) );
  AOI21D1BWP30P140LVT U32 ( .A1(n3), .A2(i_data_bus[4]), .B(n76), .ZN(n79) );
  AOI21D1BWP30P140LVT U33 ( .A1(n3), .A2(i_data_bus[14]), .B(n106), .ZN(n109)
         );
  AOI22D1BWP30P140LVT U34 ( .A1(n7), .A2(i_data_bus[111]), .B1(n221), .B2(
        i_data_bus[143]), .ZN(n222) );
  AN3D1BWP30P140LVT U35 ( .A1(n42), .A2(i_cmd[3]), .A3(i_valid[3]), .Z(n6) );
  AN2D2BWP30P140LVT U36 ( .A1(n43), .A2(n6), .Z(n7) );
  INVD1BWP30P140LVT U37 ( .I(n20), .ZN(n21) );
  INR2D1BWP30P140LVT U38 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n8) );
  INVD1BWP30P140LVT U39 ( .I(n8), .ZN(n12) );
  OR2D1BWP30P140LVT U40 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n36) );
  OR2D1BWP30P140LVT U41 ( .A1(n36), .A2(i_cmd[1]), .Z(n11) );
  ND2D1BWP30P140LVT U42 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n13) );
  NR3D0P7BWP30P140LVT U43 ( .A1(n13), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n19)
         );
  INVD1BWP30P140LVT U44 ( .I(i_cmd[2]), .ZN(n14) );
  INVD2BWP30P140LVT U45 ( .I(i_cmd[1]), .ZN(n34) );
  ND2OPTIBD2BWP30P140LVT U46 ( .A1(n14), .A2(n34), .ZN(n40) );
  NR2OPTPAD1BWP30P140LVT U47 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n17) );
  INR2D1BWP30P140LVT U48 ( .A1(i_en), .B1(rst), .ZN(n15) );
  ND2OPTIBD1BWP30P140LVT U49 ( .A1(n17), .A2(n16), .ZN(n18) );
  OR2D2BWP30P140LVT U50 ( .A1(n40), .A2(n18), .Z(n29) );
  INR2D2BWP30P140LVT U51 ( .A1(n19), .B1(n29), .ZN(n20) );
  INVD1BWP30P140LVT U52 ( .I(i_cmd[6]), .ZN(n23) );
  INR2D1BWP30P140LVT U53 ( .A1(n25), .B1(n29), .ZN(n26) );
  INR2D1BWP30P140LVT U54 ( .A1(n30), .B1(n29), .ZN(n31) );
  INVD2BWP30P140LVT U55 ( .I(n31), .ZN(n111) );
  NR4D0BWP30P140LVT U56 ( .A1(n3), .A2(n20), .A3(n2), .A4(n1), .ZN(n49) );
  INR2D4BWP30P140LVT U57 ( .A1(n33), .B1(n32), .ZN(n43) );
  INVD1BWP30P140LVT U58 ( .I(i_cmd[3]), .ZN(n41) );
  ND4D1BWP30P140LVT U59 ( .A1(n34), .A2(n41), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n35) );
  INVD1BWP30P140LVT U60 ( .I(n36), .ZN(n37) );
  ND3D2BWP30P140LVT U61 ( .A1(n37), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n38)
         );
  INVD2BWP30P140LVT U62 ( .I(n218), .ZN(n229) );
  NR2D1BWP30P140LVT U63 ( .A1(n211), .A2(n229), .ZN(n48) );
  INVD1BWP30P140LVT U64 ( .I(n40), .ZN(n42) );
  IND3D1BWP30P140LVT U65 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n44) );
  NR2D1BWP30P140LVT U66 ( .A1(n7), .A2(n231), .ZN(n47) );
  ND3D1BWP30P140LVT U67 ( .A1(n49), .A2(n48), .A3(n47), .ZN(N402) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[224]), .ZN(n55) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[192]), .ZN(n50) );
  MAOI22D1BWP30P140LVT U70 ( .A1(n1), .A2(i_data_bus[160]), .B1(n226), .B2(n50), .ZN(n54) );
  INR2D1BWP30P140LVT U71 ( .A1(i_data_bus[0]), .B1(n51), .ZN(n52) );
  INVD1BWP30P140LVT U72 ( .I(n52), .ZN(n53) );
  OA211D1BWP30P140LVT U73 ( .A1(n21), .A2(n55), .B(n54), .C(n53), .Z(n59) );
  AOI22D1BWP30P140LVT U74 ( .A1(n211), .A2(i_data_bus[64]), .B1(n229), .B2(
        i_data_bus[32]), .ZN(n58) );
  INVD2BWP30P140LVT U75 ( .I(n56), .ZN(n221) );
  AOI22D1BWP30P140LVT U76 ( .A1(n7), .A2(i_data_bus[96]), .B1(n221), .B2(
        i_data_bus[128]), .ZN(n57) );
  ND3D1BWP30P140LVT U77 ( .A1(n59), .A2(n58), .A3(n57), .ZN(N369) );
  AOI22D1BWP30P140LVT U78 ( .A1(n2), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n60) );
  IOA21D1BWP30P140LVT U79 ( .A1(n20), .A2(i_data_bus[229]), .B(n60), .ZN(n61)
         );
  AOI21D1BWP30P140LVT U80 ( .A1(n3), .A2(i_data_bus[5]), .B(n61), .ZN(n64) );
  AOI22D1BWP30P140LVT U81 ( .A1(n211), .A2(i_data_bus[69]), .B1(n229), .B2(
        i_data_bus[37]), .ZN(n63) );
  AOI22D1BWP30P140LVT U82 ( .A1(n7), .A2(i_data_bus[101]), .B1(n231), .B2(
        i_data_bus[133]), .ZN(n62) );
  ND3D1BWP30P140LVT U83 ( .A1(n64), .A2(n63), .A3(n62), .ZN(N374) );
  AOI22D1BWP30P140LVT U84 ( .A1(n2), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n65) );
  IOA21D1BWP30P140LVT U85 ( .A1(n20), .A2(i_data_bus[230]), .B(n65), .ZN(n66)
         );
  AOI21D1BWP30P140LVT U86 ( .A1(n3), .A2(i_data_bus[6]), .B(n66), .ZN(n69) );
  AOI22D1BWP30P140LVT U87 ( .A1(n211), .A2(i_data_bus[70]), .B1(n229), .B2(
        i_data_bus[38]), .ZN(n68) );
  AOI22D1BWP30P140LVT U88 ( .A1(n7), .A2(i_data_bus[102]), .B1(n221), .B2(
        i_data_bus[134]), .ZN(n67) );
  ND3D1BWP30P140LVT U89 ( .A1(n69), .A2(n68), .A3(n67), .ZN(N375) );
  AOI22D1BWP30P140LVT U90 ( .A1(n2), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n70) );
  IOA21D1BWP30P140LVT U91 ( .A1(n20), .A2(i_data_bus[232]), .B(n70), .ZN(n71)
         );
  AOI21D1BWP30P140LVT U92 ( .A1(n3), .A2(i_data_bus[8]), .B(n71), .ZN(n74) );
  AOI22D1BWP30P140LVT U93 ( .A1(n211), .A2(i_data_bus[72]), .B1(n229), .B2(
        i_data_bus[40]), .ZN(n73) );
  AOI22D1BWP30P140LVT U94 ( .A1(n7), .A2(i_data_bus[104]), .B1(n231), .B2(
        i_data_bus[136]), .ZN(n72) );
  ND3D1BWP30P140LVT U95 ( .A1(n74), .A2(n73), .A3(n72), .ZN(N377) );
  AOI22D1BWP30P140LVT U96 ( .A1(n2), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n75) );
  IOA21D1BWP30P140LVT U97 ( .A1(n20), .A2(i_data_bus[228]), .B(n75), .ZN(n76)
         );
  AOI22D1BWP30P140LVT U98 ( .A1(n211), .A2(i_data_bus[68]), .B1(n229), .B2(
        i_data_bus[36]), .ZN(n78) );
  AOI22D1BWP30P140LVT U99 ( .A1(n7), .A2(i_data_bus[100]), .B1(n221), .B2(
        i_data_bus[132]), .ZN(n77) );
  ND3D1BWP30P140LVT U100 ( .A1(n79), .A2(n78), .A3(n77), .ZN(N373) );
  AOI22D1BWP30P140LVT U101 ( .A1(n2), .A2(i_data_bus[199]), .B1(n1), .B2(
        i_data_bus[167]), .ZN(n80) );
  IOA21D1BWP30P140LVT U102 ( .A1(n20), .A2(i_data_bus[231]), .B(n80), .ZN(n81)
         );
  AOI21D1BWP30P140LVT U103 ( .A1(n3), .A2(i_data_bus[7]), .B(n81), .ZN(n84) );
  AOI22D1BWP30P140LVT U104 ( .A1(n211), .A2(i_data_bus[71]), .B1(n229), .B2(
        i_data_bus[39]), .ZN(n83) );
  AOI22D1BWP30P140LVT U105 ( .A1(n7), .A2(i_data_bus[103]), .B1(n231), .B2(
        i_data_bus[135]), .ZN(n82) );
  ND3D1BWP30P140LVT U106 ( .A1(n84), .A2(n83), .A3(n82), .ZN(N376) );
  AOI22D1BWP30P140LVT U107 ( .A1(n2), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n85) );
  IOA21D1BWP30P140LVT U108 ( .A1(n20), .A2(i_data_bus[236]), .B(n85), .ZN(n86)
         );
  AOI21D1BWP30P140LVT U109 ( .A1(n3), .A2(i_data_bus[12]), .B(n86), .ZN(n89)
         );
  AOI22D1BWP30P140LVT U110 ( .A1(n211), .A2(i_data_bus[76]), .B1(n229), .B2(
        i_data_bus[44]), .ZN(n88) );
  AOI22D1BWP30P140LVT U111 ( .A1(n7), .A2(i_data_bus[108]), .B1(n221), .B2(
        i_data_bus[140]), .ZN(n87) );
  ND3D1BWP30P140LVT U112 ( .A1(n89), .A2(n88), .A3(n87), .ZN(N381) );
  AOI22D1BWP30P140LVT U113 ( .A1(n2), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n90) );
  IOA21D1BWP30P140LVT U114 ( .A1(n20), .A2(i_data_bus[233]), .B(n90), .ZN(n91)
         );
  AOI21D1BWP30P140LVT U115 ( .A1(n3), .A2(i_data_bus[9]), .B(n91), .ZN(n94) );
  AOI22D1BWP30P140LVT U116 ( .A1(n230), .A2(i_data_bus[73]), .B1(n229), .B2(
        i_data_bus[41]), .ZN(n93) );
  AOI22D1BWP30P140LVT U117 ( .A1(n7), .A2(i_data_bus[105]), .B1(n231), .B2(
        i_data_bus[137]), .ZN(n92) );
  ND3D1BWP30P140LVT U118 ( .A1(n94), .A2(n93), .A3(n92), .ZN(N378) );
  AOI22D1BWP30P140LVT U119 ( .A1(n2), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n95) );
  IOA21D1BWP30P140LVT U120 ( .A1(n20), .A2(i_data_bus[234]), .B(n95), .ZN(n96)
         );
  AOI21D1BWP30P140LVT U121 ( .A1(n3), .A2(i_data_bus[10]), .B(n96), .ZN(n99)
         );
  AOI22D1BWP30P140LVT U122 ( .A1(n211), .A2(i_data_bus[74]), .B1(n229), .B2(
        i_data_bus[42]), .ZN(n98) );
  AOI22D1BWP30P140LVT U123 ( .A1(n7), .A2(i_data_bus[106]), .B1(n221), .B2(
        i_data_bus[138]), .ZN(n97) );
  ND3D1BWP30P140LVT U124 ( .A1(n99), .A2(n98), .A3(n97), .ZN(N379) );
  AOI22D1BWP30P140LVT U125 ( .A1(n2), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n100) );
  IOA21D1BWP30P140LVT U126 ( .A1(n20), .A2(i_data_bus[235]), .B(n100), .ZN(
        n101) );
  AOI21D1BWP30P140LVT U127 ( .A1(n3), .A2(i_data_bus[11]), .B(n101), .ZN(n104)
         );
  AOI22D1BWP30P140LVT U128 ( .A1(n230), .A2(i_data_bus[75]), .B1(n229), .B2(
        i_data_bus[43]), .ZN(n103) );
  AOI22D1BWP30P140LVT U129 ( .A1(n7), .A2(i_data_bus[107]), .B1(n231), .B2(
        i_data_bus[139]), .ZN(n102) );
  ND3D1BWP30P140LVT U130 ( .A1(n104), .A2(n103), .A3(n102), .ZN(N380) );
  AOI22D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[206]), .B1(n1), .B2(
        i_data_bus[174]), .ZN(n105) );
  IOA21D1BWP30P140LVT U132 ( .A1(n20), .A2(i_data_bus[238]), .B(n105), .ZN(
        n106) );
  AOI22D1BWP30P140LVT U133 ( .A1(n230), .A2(i_data_bus[78]), .B1(n229), .B2(
        i_data_bus[46]), .ZN(n108) );
  AOI22D1BWP30P140LVT U134 ( .A1(n7), .A2(i_data_bus[110]), .B1(n221), .B2(
        i_data_bus[142]), .ZN(n107) );
  ND3D1BWP30P140LVT U135 ( .A1(n109), .A2(n108), .A3(n107), .ZN(N383) );
  INVD1BWP30P140LVT U136 ( .I(i_data_bus[173]), .ZN(n110) );
  IOA21D1BWP30P140LVT U137 ( .A1(n20), .A2(i_data_bus[237]), .B(n112), .ZN(
        n113) );
  AOI21D1BWP30P140LVT U138 ( .A1(n3), .A2(i_data_bus[13]), .B(n113), .ZN(n116)
         );
  AOI22D1BWP30P140LVT U139 ( .A1(n230), .A2(i_data_bus[77]), .B1(n229), .B2(
        i_data_bus[45]), .ZN(n115) );
  AOI22D1BWP30P140LVT U140 ( .A1(n7), .A2(i_data_bus[109]), .B1(n231), .B2(
        i_data_bus[141]), .ZN(n114) );
  ND3D1BWP30P140LVT U141 ( .A1(n116), .A2(n115), .A3(n114), .ZN(N382) );
  AOI22D1BWP30P140LVT U142 ( .A1(n2), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n117) );
  IOA21D1BWP30P140LVT U143 ( .A1(n20), .A2(i_data_bus[242]), .B(n117), .ZN(
        n118) );
  AOI21D1BWP30P140LVT U144 ( .A1(n3), .A2(i_data_bus[18]), .B(n118), .ZN(n121)
         );
  AOI22D1BWP30P140LVT U145 ( .A1(n230), .A2(i_data_bus[82]), .B1(n229), .B2(
        i_data_bus[50]), .ZN(n120) );
  AOI22D1BWP30P140LVT U146 ( .A1(n7), .A2(i_data_bus[114]), .B1(n221), .B2(
        i_data_bus[146]), .ZN(n119) );
  ND3D1BWP30P140LVT U147 ( .A1(n121), .A2(n120), .A3(n119), .ZN(N387) );
  AOI22D1BWP30P140LVT U148 ( .A1(n2), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n122) );
  IOA21D1BWP30P140LVT U149 ( .A1(n20), .A2(i_data_bus[241]), .B(n122), .ZN(
        n123) );
  AOI21D1BWP30P140LVT U150 ( .A1(n3), .A2(i_data_bus[17]), .B(n123), .ZN(n126)
         );
  AOI22D1BWP30P140LVT U151 ( .A1(n230), .A2(i_data_bus[81]), .B1(n229), .B2(
        i_data_bus[49]), .ZN(n125) );
  AOI22D1BWP30P140LVT U152 ( .A1(n7), .A2(i_data_bus[113]), .B1(n221), .B2(
        i_data_bus[145]), .ZN(n124) );
  ND3D1BWP30P140LVT U153 ( .A1(n126), .A2(n125), .A3(n124), .ZN(N386) );
  AOI22D1BWP30P140LVT U154 ( .A1(n2), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n127) );
  IOA21D1BWP30P140LVT U155 ( .A1(n20), .A2(i_data_bus[248]), .B(n127), .ZN(
        n128) );
  AOI21D1BWP30P140LVT U156 ( .A1(n3), .A2(i_data_bus[24]), .B(n128), .ZN(n131)
         );
  AOI22D1BWP30P140LVT U157 ( .A1(n230), .A2(i_data_bus[88]), .B1(n229), .B2(
        i_data_bus[56]), .ZN(n130) );
  AOI22D1BWP30P140LVT U158 ( .A1(n7), .A2(i_data_bus[120]), .B1(n231), .B2(
        i_data_bus[152]), .ZN(n129) );
  ND3D1BWP30P140LVT U159 ( .A1(n131), .A2(n130), .A3(n129), .ZN(N393) );
  AOI22D1BWP30P140LVT U160 ( .A1(n2), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n132) );
  IOA21D1BWP30P140LVT U161 ( .A1(n20), .A2(i_data_bus[247]), .B(n132), .ZN(
        n133) );
  AOI21D1BWP30P140LVT U162 ( .A1(n3), .A2(i_data_bus[23]), .B(n133), .ZN(n136)
         );
  AOI22D1BWP30P140LVT U163 ( .A1(n230), .A2(i_data_bus[87]), .B1(n229), .B2(
        i_data_bus[55]), .ZN(n135) );
  AOI22D1BWP30P140LVT U164 ( .A1(n7), .A2(i_data_bus[119]), .B1(n221), .B2(
        i_data_bus[151]), .ZN(n134) );
  ND3D1BWP30P140LVT U165 ( .A1(n136), .A2(n135), .A3(n134), .ZN(N392) );
  AOI22D1BWP30P140LVT U166 ( .A1(n2), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n137) );
  IOA21D1BWP30P140LVT U167 ( .A1(n20), .A2(i_data_bus[246]), .B(n137), .ZN(
        n138) );
  AOI21D1BWP30P140LVT U168 ( .A1(n3), .A2(i_data_bus[22]), .B(n138), .ZN(n141)
         );
  AOI22D1BWP30P140LVT U169 ( .A1(n230), .A2(i_data_bus[86]), .B1(n229), .B2(
        i_data_bus[54]), .ZN(n140) );
  AOI22D1BWP30P140LVT U170 ( .A1(n7), .A2(i_data_bus[118]), .B1(n231), .B2(
        i_data_bus[150]), .ZN(n139) );
  ND3D1BWP30P140LVT U171 ( .A1(n141), .A2(n140), .A3(n139), .ZN(N391) );
  AOI22D1BWP30P140LVT U172 ( .A1(n2), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n142) );
  IOA21D1BWP30P140LVT U173 ( .A1(n20), .A2(i_data_bus[245]), .B(n142), .ZN(
        n143) );
  AOI21D1BWP30P140LVT U174 ( .A1(n3), .A2(i_data_bus[21]), .B(n143), .ZN(n146)
         );
  AOI22D1BWP30P140LVT U175 ( .A1(n230), .A2(i_data_bus[85]), .B1(n229), .B2(
        i_data_bus[53]), .ZN(n145) );
  AOI22D1BWP30P140LVT U176 ( .A1(n7), .A2(i_data_bus[117]), .B1(n221), .B2(
        i_data_bus[149]), .ZN(n144) );
  ND3D1BWP30P140LVT U177 ( .A1(n146), .A2(n145), .A3(n144), .ZN(N390) );
  AOI22D1BWP30P140LVT U178 ( .A1(n2), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n147) );
  IOA21D1BWP30P140LVT U179 ( .A1(n20), .A2(i_data_bus[244]), .B(n147), .ZN(
        n148) );
  AOI21D1BWP30P140LVT U180 ( .A1(n3), .A2(i_data_bus[20]), .B(n148), .ZN(n151)
         );
  AOI22D1BWP30P140LVT U181 ( .A1(n230), .A2(i_data_bus[84]), .B1(n229), .B2(
        i_data_bus[52]), .ZN(n150) );
  AOI22D1BWP30P140LVT U182 ( .A1(n7), .A2(i_data_bus[116]), .B1(n231), .B2(
        i_data_bus[148]), .ZN(n149) );
  ND3D1BWP30P140LVT U183 ( .A1(n151), .A2(n150), .A3(n149), .ZN(N389) );
  AOI22D1BWP30P140LVT U184 ( .A1(n2), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n152) );
  IOA21D1BWP30P140LVT U185 ( .A1(n20), .A2(i_data_bus[243]), .B(n152), .ZN(
        n153) );
  AOI21D1BWP30P140LVT U186 ( .A1(n3), .A2(i_data_bus[19]), .B(n153), .ZN(n156)
         );
  AOI22D1BWP30P140LVT U187 ( .A1(n230), .A2(i_data_bus[83]), .B1(n229), .B2(
        i_data_bus[51]), .ZN(n155) );
  AOI22D1BWP30P140LVT U188 ( .A1(n7), .A2(i_data_bus[115]), .B1(n221), .B2(
        i_data_bus[147]), .ZN(n154) );
  ND3D1BWP30P140LVT U189 ( .A1(n156), .A2(n155), .A3(n154), .ZN(N388) );
  INVD1BWP30P140LVT U190 ( .I(i_data_bus[195]), .ZN(n157) );
  MAOI22D1BWP30P140LVT U191 ( .A1(n1), .A2(i_data_bus[163]), .B1(n226), .B2(
        n157), .ZN(n158) );
  IOA21D1BWP30P140LVT U192 ( .A1(n20), .A2(i_data_bus[227]), .B(n158), .ZN(
        n159) );
  AOI21D1BWP30P140LVT U193 ( .A1(n3), .A2(i_data_bus[3]), .B(n159), .ZN(n162)
         );
  AOI22D1BWP30P140LVT U194 ( .A1(n211), .A2(i_data_bus[67]), .B1(n229), .B2(
        i_data_bus[35]), .ZN(n161) );
  AOI22D1BWP30P140LVT U195 ( .A1(n7), .A2(i_data_bus[99]), .B1(n221), .B2(
        i_data_bus[131]), .ZN(n160) );
  ND3D1BWP30P140LVT U196 ( .A1(n162), .A2(n161), .A3(n160), .ZN(N372) );
  INVD1BWP30P140LVT U197 ( .I(i_data_bus[193]), .ZN(n163) );
  MAOI22D1BWP30P140LVT U198 ( .A1(n1), .A2(i_data_bus[161]), .B1(n226), .B2(
        n163), .ZN(n164) );
  IOA21D1BWP30P140LVT U199 ( .A1(n20), .A2(i_data_bus[225]), .B(n164), .ZN(
        n165) );
  AOI21D1BWP30P140LVT U200 ( .A1(n3), .A2(i_data_bus[1]), .B(n165), .ZN(n168)
         );
  AOI22D1BWP30P140LVT U201 ( .A1(n230), .A2(i_data_bus[65]), .B1(n229), .B2(
        i_data_bus[33]), .ZN(n167) );
  AOI22D1BWP30P140LVT U202 ( .A1(n7), .A2(i_data_bus[97]), .B1(n231), .B2(
        i_data_bus[129]), .ZN(n166) );
  ND3D1BWP30P140LVT U203 ( .A1(n168), .A2(n167), .A3(n166), .ZN(N370) );
  INVD1BWP30P140LVT U204 ( .I(i_data_bus[194]), .ZN(n169) );
  MAOI22D1BWP30P140LVT U205 ( .A1(n1), .A2(i_data_bus[162]), .B1(n226), .B2(
        n169), .ZN(n170) );
  IOA21D1BWP30P140LVT U206 ( .A1(n20), .A2(i_data_bus[226]), .B(n170), .ZN(
        n171) );
  AOI21D1BWP30P140LVT U207 ( .A1(n3), .A2(i_data_bus[2]), .B(n171), .ZN(n175)
         );
  AOI22D1BWP30P140LVT U208 ( .A1(n172), .A2(i_data_bus[66]), .B1(n229), .B2(
        i_data_bus[34]), .ZN(n174) );
  AOI22D1BWP30P140LVT U209 ( .A1(n7), .A2(i_data_bus[98]), .B1(n221), .B2(
        i_data_bus[130]), .ZN(n173) );
  ND3D1BWP30P140LVT U210 ( .A1(n175), .A2(n174), .A3(n173), .ZN(N371) );
  INVD1BWP30P140LVT U211 ( .I(i_data_bus[222]), .ZN(n176) );
  MAOI22D1BWP30P140LVT U212 ( .A1(n1), .A2(i_data_bus[190]), .B1(n226), .B2(
        n176), .ZN(n177) );
  IOA21D1BWP30P140LVT U213 ( .A1(n20), .A2(i_data_bus[254]), .B(n177), .ZN(
        n178) );
  AOI21D1BWP30P140LVT U214 ( .A1(n3), .A2(i_data_bus[30]), .B(n178), .ZN(n181)
         );
  AOI22D1BWP30P140LVT U215 ( .A1(n211), .A2(i_data_bus[94]), .B1(n229), .B2(
        i_data_bus[62]), .ZN(n180) );
  AOI22D1BWP30P140LVT U216 ( .A1(n7), .A2(i_data_bus[126]), .B1(n231), .B2(
        i_data_bus[158]), .ZN(n179) );
  ND3D1BWP30P140LVT U217 ( .A1(n181), .A2(n180), .A3(n179), .ZN(N399) );
  AOI22D1BWP30P140LVT U218 ( .A1(n2), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n182) );
  IOA21D1BWP30P140LVT U219 ( .A1(n20), .A2(i_data_bus[251]), .B(n182), .ZN(
        n183) );
  AOI21D1BWP30P140LVT U220 ( .A1(n3), .A2(i_data_bus[27]), .B(n183), .ZN(n186)
         );
  AOI22D1BWP30P140LVT U221 ( .A1(n211), .A2(i_data_bus[91]), .B1(n229), .B2(
        i_data_bus[59]), .ZN(n185) );
  AOI22D1BWP30P140LVT U222 ( .A1(n7), .A2(i_data_bus[123]), .B1(n221), .B2(
        i_data_bus[155]), .ZN(n184) );
  ND3D1BWP30P140LVT U223 ( .A1(n186), .A2(n185), .A3(n184), .ZN(N396) );
  AOI22D1BWP30P140LVT U224 ( .A1(n2), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n187) );
  IOA21D1BWP30P140LVT U225 ( .A1(n20), .A2(i_data_bus[249]), .B(n187), .ZN(
        n188) );
  AOI21D1BWP30P140LVT U226 ( .A1(n3), .A2(i_data_bus[25]), .B(n188), .ZN(n191)
         );
  AOI22D1BWP30P140LVT U227 ( .A1(n230), .A2(i_data_bus[89]), .B1(n229), .B2(
        i_data_bus[57]), .ZN(n190) );
  AOI22D1BWP30P140LVT U228 ( .A1(n7), .A2(i_data_bus[121]), .B1(n231), .B2(
        i_data_bus[153]), .ZN(n189) );
  ND3D1BWP30P140LVT U229 ( .A1(n191), .A2(n190), .A3(n189), .ZN(N394) );
  AOI22D1BWP30P140LVT U230 ( .A1(n2), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n192) );
  IOA21D1BWP30P140LVT U231 ( .A1(n20), .A2(i_data_bus[250]), .B(n192), .ZN(
        n193) );
  AOI21D1BWP30P140LVT U232 ( .A1(n3), .A2(i_data_bus[26]), .B(n193), .ZN(n196)
         );
  AOI22D1BWP30P140LVT U233 ( .A1(n211), .A2(i_data_bus[90]), .B1(n229), .B2(
        i_data_bus[58]), .ZN(n195) );
  AOI22D1BWP30P140LVT U234 ( .A1(n7), .A2(i_data_bus[122]), .B1(n221), .B2(
        i_data_bus[154]), .ZN(n194) );
  ND3D1BWP30P140LVT U235 ( .A1(n196), .A2(n195), .A3(n194), .ZN(N395) );
  AOI22D1BWP30P140LVT U236 ( .A1(n2), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n197) );
  IOA21D1BWP30P140LVT U237 ( .A1(n20), .A2(i_data_bus[252]), .B(n197), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U238 ( .A1(n3), .A2(i_data_bus[28]), .B(n198), .ZN(n201)
         );
  AOI22D1BWP30P140LVT U239 ( .A1(n211), .A2(i_data_bus[92]), .B1(n229), .B2(
        i_data_bus[60]), .ZN(n200) );
  AOI22D1BWP30P140LVT U240 ( .A1(n7), .A2(i_data_bus[124]), .B1(n231), .B2(
        i_data_bus[156]), .ZN(n199) );
  ND3D1BWP30P140LVT U241 ( .A1(n201), .A2(n200), .A3(n199), .ZN(N397) );
  INVD1BWP30P140LVT U242 ( .I(i_data_bus[221]), .ZN(n202) );
  MAOI22D1BWP30P140LVT U243 ( .A1(n1), .A2(i_data_bus[189]), .B1(n226), .B2(
        n202), .ZN(n203) );
  IOA21D1BWP30P140LVT U244 ( .A1(n20), .A2(i_data_bus[253]), .B(n203), .ZN(
        n204) );
  AOI21D1BWP30P140LVT U245 ( .A1(n3), .A2(i_data_bus[29]), .B(n204), .ZN(n207)
         );
  AOI22D1BWP30P140LVT U246 ( .A1(n211), .A2(i_data_bus[93]), .B1(n229), .B2(
        i_data_bus[61]), .ZN(n206) );
  AOI22D1BWP30P140LVT U247 ( .A1(n7), .A2(i_data_bus[125]), .B1(n221), .B2(
        i_data_bus[157]), .ZN(n205) );
  ND3D1BWP30P140LVT U248 ( .A1(n207), .A2(n206), .A3(n205), .ZN(N398) );
  INVD1BWP30P140LVT U249 ( .I(i_data_bus[223]), .ZN(n208) );
  MAOI22D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[191]), .B1(n226), .B2(
        n208), .ZN(n209) );
  IOA21D1BWP30P140LVT U251 ( .A1(n20), .A2(i_data_bus[255]), .B(n209), .ZN(
        n210) );
  AOI21D1BWP30P140LVT U252 ( .A1(n3), .A2(i_data_bus[31]), .B(n210), .ZN(n214)
         );
  AOI22D1BWP30P140LVT U253 ( .A1(n211), .A2(i_data_bus[95]), .B1(n229), .B2(
        i_data_bus[63]), .ZN(n213) );
  AOI22D1BWP30P140LVT U254 ( .A1(n7), .A2(i_data_bus[127]), .B1(n231), .B2(
        i_data_bus[159]), .ZN(n212) );
  ND3D1BWP30P140LVT U255 ( .A1(n214), .A2(n213), .A3(n212), .ZN(N400) );
  AOI22D1BWP30P140LVT U256 ( .A1(n2), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n215) );
  IOA21D1BWP30P140LVT U257 ( .A1(n20), .A2(i_data_bus[239]), .B(n215), .ZN(
        n216) );
  AOI21D1BWP30P140LVT U258 ( .A1(n3), .A2(i_data_bus[15]), .B(n216), .ZN(n224)
         );
  INVD1BWP30P140LVT U259 ( .I(i_data_bus[79]), .ZN(n219) );
  INVD1BWP30P140LVT U260 ( .I(i_data_bus[47]), .ZN(n217) );
  OA22D1BWP30P140LVT U261 ( .A1(n220), .A2(n219), .B1(n218), .B2(n217), .Z(
        n223) );
  ND3D1BWP30P140LVT U262 ( .A1(n224), .A2(n223), .A3(n222), .ZN(N384) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[208]), .ZN(n225) );
  MAOI22D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[176]), .B1(n226), .B2(
        n225), .ZN(n227) );
  IOA21D1BWP30P140LVT U265 ( .A1(n20), .A2(i_data_bus[240]), .B(n227), .ZN(
        n228) );
  AOI21D1BWP30P140LVT U266 ( .A1(n3), .A2(i_data_bus[16]), .B(n228), .ZN(n234)
         );
  AOI22D1BWP30P140LVT U267 ( .A1(n230), .A2(i_data_bus[80]), .B1(n229), .B2(
        i_data_bus[48]), .ZN(n233) );
  AOI22D1BWP30P140LVT U268 ( .A1(n7), .A2(i_data_bus[112]), .B1(n231), .B2(
        i_data_bus[144]), .ZN(n232) );
  ND3D1BWP30P140LVT U269 ( .A1(n234), .A2(n233), .A3(n232), .ZN(N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_6 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n52), .ZN(n4) );
  INR2D4BWP30P140LVT U4 ( .A1(n37), .B1(n32), .ZN(n227) );
  INVD6BWP30P140LVT U5 ( .I(n142), .ZN(n2) );
  INVD2BWP30P140LVT U6 ( .I(n25), .ZN(n142) );
  NR2D1BWP30P140LVT U7 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n27) );
  ND2OPTIBD1BWP30P140LVT U8 ( .A1(n41), .A2(n40), .ZN(n52) );
  OR4D1BWP30P140LVT U9 ( .A1(n9), .A2(n26), .A3(n10), .A4(n5), .Z(n1) );
  INVD2BWP30P140LVT U10 ( .I(n1), .ZN(n3) );
  INR4D1BWP30P140LVT U11 ( .A1(i_valid[6]), .B1(i_cmd[5]), .B2(i_cmd[7]), .B3(
        n19), .ZN(n20) );
  AOI21D1BWP30P140LVT U12 ( .A1(n3), .A2(i_data_bus[6]), .B(n62), .ZN(n65) );
  INVD1BWP30P140LVT U13 ( .I(n227), .ZN(n216) );
  ND2OPTIBD2BWP30P140LVT U14 ( .A1(n8), .A2(n7), .ZN(n26) );
  INR2D1BWP30P140LVT U15 ( .A1(i_en), .B1(rst), .ZN(n7) );
  NR3D1P5BWP30P140LVT U16 ( .A1(i_cmd[7]), .A2(i_cmd[6]), .A3(i_cmd[5]), .ZN(
        n8) );
  INVD1BWP30P140LVT U17 ( .I(n38), .ZN(n51) );
  INR2D1BWP30P140LVT U18 ( .A1(n37), .B1(n36), .ZN(n38) );
  NR3D0P7BWP30P140LVT U19 ( .A1(n22), .A2(i_cmd[6]), .A3(i_cmd[7]), .ZN(n24)
         );
  ND2D1BWP30P140LVT U20 ( .A1(i_valid[5]), .A2(i_cmd[5]), .ZN(n22) );
  NR2D1BWP30P140LVT U21 ( .A1(n9), .A2(n26), .ZN(n41) );
  INR2D2BWP30P140LVT U22 ( .A1(n27), .B1(n26), .ZN(n37) );
  INVD1BWP30P140LVT U23 ( .I(n1), .ZN(n201) );
  INVD2BWP30P140LVT U24 ( .I(n51), .ZN(n219) );
  ND2D1BWP30P140LVT U25 ( .A1(n15), .A2(n14), .ZN(n16) );
  INVD2BWP30P140LVT U26 ( .I(n51), .ZN(n228) );
  ND3D2BWP30P140LVT U27 ( .A1(n31), .A2(i_valid[1]), .A3(i_cmd[1]), .ZN(n32)
         );
  INVD1BWP30P140LVT U28 ( .I(n30), .ZN(n31) );
  NR2D1BWP30P140LVT U29 ( .A1(n219), .A2(n4), .ZN(n42) );
  AOI22D1BWP30P140LVT U30 ( .A1(n208), .A2(i_data_bus[94]), .B1(n227), .B2(
        i_data_bus[62]), .ZN(n191) );
  INVD1BWP30P140LVT U31 ( .I(i_cmd[0]), .ZN(n5) );
  INR2D4BWP30P140LVT U32 ( .A1(n17), .B1(n23), .ZN(n18) );
  INVD1BWP30P140LVT U33 ( .I(n208), .ZN(n218) );
  INR2D1BWP30P140LVT U34 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n6) );
  INVD1BWP30P140LVT U35 ( .I(n6), .ZN(n10) );
  OR2D1BWP30P140LVT U36 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n30) );
  OR2D1BWP30P140LVT U37 ( .A1(n30), .A2(i_cmd[1]), .Z(n9) );
  ND2D1BWP30P140LVT U38 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n11) );
  NR3D0P7BWP30P140LVT U39 ( .A1(n11), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n17)
         );
  INVD1BWP30P140LVT U40 ( .I(i_cmd[2]), .ZN(n12) );
  INVD1BWP30P140LVT U41 ( .I(i_cmd[1]), .ZN(n28) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n12), .A2(n28), .ZN(n33) );
  NR2D1BWP30P140LVT U43 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n15) );
  INR2D1BWP30P140LVT U44 ( .A1(i_en), .B1(rst), .ZN(n13) );
  INR2D1BWP30P140LVT U45 ( .A1(n13), .B1(i_cmd[3]), .ZN(n14) );
  OR2D4BWP30P140LVT U46 ( .A1(n33), .A2(n16), .Z(n23) );
  INVD1BWP30P140LVT U47 ( .I(i_cmd[6]), .ZN(n19) );
  INR2D2BWP30P140LVT U48 ( .A1(n20), .B1(n23), .ZN(n21) );
  INVD4BWP30P140LVT U49 ( .I(n21), .ZN(n224) );
  INVD2BWP30P140LVT U50 ( .I(n224), .ZN(n205) );
  INR2D2BWP30P140LVT U51 ( .A1(n24), .B1(n23), .ZN(n25) );
  NR4D0BWP30P140LVT U52 ( .A1(n201), .A2(n18), .A3(n205), .A4(n2), .ZN(n44) );
  INVD1BWP30P140LVT U53 ( .I(i_cmd[3]), .ZN(n34) );
  ND4D1BWP30P140LVT U54 ( .A1(n28), .A2(n34), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n29) );
  INR2D4BWP30P140LVT U55 ( .A1(n37), .B1(n29), .ZN(n208) );
  NR2D1BWP30P140LVT U56 ( .A1(n208), .A2(n227), .ZN(n43) );
  INVD1BWP30P140LVT U57 ( .I(n33), .ZN(n35) );
  ND3D1BWP30P140LVT U58 ( .A1(n35), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n36)
         );
  IND3D1BWP30P140LVT U59 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n39) );
  INVD1BWP30P140LVT U60 ( .I(n39), .ZN(n40) );
  ND3D1BWP30P140LVT U61 ( .A1(n44), .A2(n43), .A3(n42), .ZN(N402) );
  INVD1BWP30P140LVT U62 ( .I(n18), .ZN(n50) );
  INVD1BWP30P140LVT U63 ( .I(i_data_bus[224]), .ZN(n49) );
  INVD1BWP30P140LVT U64 ( .I(i_data_bus[192]), .ZN(n45) );
  MAOI22D1BWP30P140LVT U65 ( .A1(n2), .A2(i_data_bus[160]), .B1(n224), .B2(n45), .ZN(n48) );
  INR2D1BWP30P140LVT U66 ( .A1(i_data_bus[0]), .B1(n1), .ZN(n46) );
  INVD1BWP30P140LVT U67 ( .I(n46), .ZN(n47) );
  OA211D1BWP30P140LVT U68 ( .A1(n50), .A2(n49), .B(n48), .C(n47), .Z(n55) );
  AOI22D1BWP30P140LVT U69 ( .A1(n208), .A2(i_data_bus[64]), .B1(n227), .B2(
        i_data_bus[32]), .ZN(n54) );
  AOI22D1BWP30P140LVT U70 ( .A1(n228), .A2(i_data_bus[96]), .B1(n4), .B2(
        i_data_bus[128]), .ZN(n53) );
  ND3D1BWP30P140LVT U71 ( .A1(n55), .A2(n54), .A3(n53), .ZN(N369) );
  INVD2BWP30P140LVT U72 ( .I(n224), .ZN(n212) );
  AOI22D1BWP30P140LVT U73 ( .A1(n212), .A2(i_data_bus[196]), .B1(n2), .B2(
        i_data_bus[164]), .ZN(n56) );
  IOA21D1BWP30P140LVT U74 ( .A1(n18), .A2(i_data_bus[228]), .B(n56), .ZN(n57)
         );
  AOI21D1BWP30P140LVT U75 ( .A1(n201), .A2(i_data_bus[4]), .B(n57), .ZN(n60)
         );
  AOI22D1BWP30P140LVT U76 ( .A1(n208), .A2(i_data_bus[68]), .B1(n227), .B2(
        i_data_bus[36]), .ZN(n59) );
  AOI22D1BWP30P140LVT U77 ( .A1(n228), .A2(i_data_bus[100]), .B1(n4), .B2(
        i_data_bus[132]), .ZN(n58) );
  ND3D1BWP30P140LVT U78 ( .A1(n60), .A2(n59), .A3(n58), .ZN(N373) );
  AOI22D1BWP30P140LVT U79 ( .A1(n212), .A2(i_data_bus[198]), .B1(n2), .B2(
        i_data_bus[166]), .ZN(n61) );
  IOA21D1BWP30P140LVT U80 ( .A1(n18), .A2(i_data_bus[230]), .B(n61), .ZN(n62)
         );
  AOI22D1BWP30P140LVT U81 ( .A1(n208), .A2(i_data_bus[70]), .B1(n227), .B2(
        i_data_bus[38]), .ZN(n64) );
  AOI22D1BWP30P140LVT U82 ( .A1(n228), .A2(i_data_bus[102]), .B1(n4), .B2(
        i_data_bus[134]), .ZN(n63) );
  ND3D1BWP30P140LVT U83 ( .A1(n65), .A2(n64), .A3(n63), .ZN(N375) );
  AOI22D1BWP30P140LVT U84 ( .A1(n212), .A2(i_data_bus[197]), .B1(n2), .B2(
        i_data_bus[165]), .ZN(n66) );
  IOA21D1BWP30P140LVT U85 ( .A1(n18), .A2(i_data_bus[229]), .B(n66), .ZN(n67)
         );
  AOI21D1BWP30P140LVT U86 ( .A1(n3), .A2(i_data_bus[5]), .B(n67), .ZN(n70) );
  AOI22D1BWP30P140LVT U87 ( .A1(n208), .A2(i_data_bus[69]), .B1(n227), .B2(
        i_data_bus[37]), .ZN(n69) );
  AOI22D1BWP30P140LVT U88 ( .A1(n228), .A2(i_data_bus[101]), .B1(n4), .B2(
        i_data_bus[133]), .ZN(n68) );
  ND3D1BWP30P140LVT U89 ( .A1(n70), .A2(n69), .A3(n68), .ZN(N374) );
  AOI22D1BWP30P140LVT U90 ( .A1(n212), .A2(i_data_bus[204]), .B1(n2), .B2(
        i_data_bus[172]), .ZN(n71) );
  IOA21D1BWP30P140LVT U91 ( .A1(n18), .A2(i_data_bus[236]), .B(n71), .ZN(n72)
         );
  AOI21D1BWP30P140LVT U92 ( .A1(n201), .A2(i_data_bus[12]), .B(n72), .ZN(n75)
         );
  AOI22D1BWP30P140LVT U93 ( .A1(n208), .A2(i_data_bus[76]), .B1(n227), .B2(
        i_data_bus[44]), .ZN(n74) );
  AOI22D1BWP30P140LVT U94 ( .A1(n228), .A2(i_data_bus[108]), .B1(n4), .B2(
        i_data_bus[140]), .ZN(n73) );
  ND3D1BWP30P140LVT U95 ( .A1(n75), .A2(n74), .A3(n73), .ZN(N381) );
  AOI22D1BWP30P140LVT U96 ( .A1(n212), .A2(i_data_bus[203]), .B1(n2), .B2(
        i_data_bus[171]), .ZN(n76) );
  IOA21D1BWP30P140LVT U97 ( .A1(n18), .A2(i_data_bus[235]), .B(n76), .ZN(n77)
         );
  AOI21D1BWP30P140LVT U98 ( .A1(n3), .A2(i_data_bus[11]), .B(n77), .ZN(n80) );
  AOI22D1BWP30P140LVT U99 ( .A1(n208), .A2(i_data_bus[75]), .B1(n227), .B2(
        i_data_bus[43]), .ZN(n79) );
  AOI22D1BWP30P140LVT U100 ( .A1(n228), .A2(i_data_bus[107]), .B1(n4), .B2(
        i_data_bus[139]), .ZN(n78) );
  ND3D1BWP30P140LVT U101 ( .A1(n80), .A2(n79), .A3(n78), .ZN(N380) );
  AOI22D1BWP30P140LVT U102 ( .A1(n212), .A2(i_data_bus[202]), .B1(n2), .B2(
        i_data_bus[170]), .ZN(n81) );
  IOA21D1BWP30P140LVT U103 ( .A1(n18), .A2(i_data_bus[234]), .B(n81), .ZN(n82)
         );
  AOI21D1BWP30P140LVT U104 ( .A1(n3), .A2(i_data_bus[10]), .B(n82), .ZN(n85)
         );
  AOI22D1BWP30P140LVT U105 ( .A1(n208), .A2(i_data_bus[74]), .B1(n227), .B2(
        i_data_bus[42]), .ZN(n84) );
  AOI22D1BWP30P140LVT U106 ( .A1(n228), .A2(i_data_bus[106]), .B1(n4), .B2(
        i_data_bus[138]), .ZN(n83) );
  ND3D1BWP30P140LVT U107 ( .A1(n85), .A2(n84), .A3(n83), .ZN(N379) );
  AOI22D1BWP30P140LVT U108 ( .A1(n212), .A2(i_data_bus[199]), .B1(n2), .B2(
        i_data_bus[167]), .ZN(n86) );
  IOA21D1BWP30P140LVT U109 ( .A1(n18), .A2(i_data_bus[231]), .B(n86), .ZN(n87)
         );
  AOI21D1BWP30P140LVT U110 ( .A1(n201), .A2(i_data_bus[7]), .B(n87), .ZN(n90)
         );
  AOI22D1BWP30P140LVT U111 ( .A1(n208), .A2(i_data_bus[71]), .B1(n227), .B2(
        i_data_bus[39]), .ZN(n89) );
  AOI22D1BWP30P140LVT U112 ( .A1(n228), .A2(i_data_bus[103]), .B1(n4), .B2(
        i_data_bus[135]), .ZN(n88) );
  ND3D1BWP30P140LVT U113 ( .A1(n90), .A2(n89), .A3(n88), .ZN(N376) );
  AOI22D1BWP30P140LVT U114 ( .A1(n212), .A2(i_data_bus[200]), .B1(n2), .B2(
        i_data_bus[168]), .ZN(n91) );
  IOA21D1BWP30P140LVT U115 ( .A1(n18), .A2(i_data_bus[232]), .B(n91), .ZN(n92)
         );
  AOI21D1BWP30P140LVT U116 ( .A1(n3), .A2(i_data_bus[8]), .B(n92), .ZN(n95) );
  AOI22D1BWP30P140LVT U117 ( .A1(n208), .A2(i_data_bus[72]), .B1(n227), .B2(
        i_data_bus[40]), .ZN(n94) );
  AOI22D1BWP30P140LVT U118 ( .A1(n228), .A2(i_data_bus[104]), .B1(n4), .B2(
        i_data_bus[136]), .ZN(n93) );
  ND3D1BWP30P140LVT U119 ( .A1(n95), .A2(n94), .A3(n93), .ZN(N377) );
  AOI22D1BWP30P140LVT U120 ( .A1(n212), .A2(i_data_bus[201]), .B1(n2), .B2(
        i_data_bus[169]), .ZN(n96) );
  IOA21D1BWP30P140LVT U121 ( .A1(n18), .A2(i_data_bus[233]), .B(n96), .ZN(n97)
         );
  AOI21D1BWP30P140LVT U122 ( .A1(n3), .A2(i_data_bus[9]), .B(n97), .ZN(n100)
         );
  AOI22D1BWP30P140LVT U123 ( .A1(n208), .A2(i_data_bus[73]), .B1(n227), .B2(
        i_data_bus[41]), .ZN(n99) );
  AOI22D1BWP30P140LVT U124 ( .A1(n228), .A2(i_data_bus[105]), .B1(n4), .B2(
        i_data_bus[137]), .ZN(n98) );
  ND3D1BWP30P140LVT U125 ( .A1(n100), .A2(n99), .A3(n98), .ZN(N378) );
  AOI22D1BWP30P140LVT U126 ( .A1(n212), .A2(i_data_bus[206]), .B1(n2), .B2(
        i_data_bus[174]), .ZN(n101) );
  IOA21D1BWP30P140LVT U127 ( .A1(n18), .A2(i_data_bus[238]), .B(n101), .ZN(
        n102) );
  AOI21D1BWP30P140LVT U128 ( .A1(n201), .A2(i_data_bus[14]), .B(n102), .ZN(
        n105) );
  AOI22D1BWP30P140LVT U129 ( .A1(n208), .A2(i_data_bus[78]), .B1(n227), .B2(
        i_data_bus[46]), .ZN(n104) );
  AOI22D1BWP30P140LVT U130 ( .A1(n219), .A2(i_data_bus[110]), .B1(n4), .B2(
        i_data_bus[142]), .ZN(n103) );
  ND3D1BWP30P140LVT U131 ( .A1(n105), .A2(n104), .A3(n103), .ZN(N383) );
  AOI22D1BWP30P140LVT U132 ( .A1(n205), .A2(i_data_bus[213]), .B1(n2), .B2(
        i_data_bus[181]), .ZN(n106) );
  IOA21D1BWP30P140LVT U133 ( .A1(n18), .A2(i_data_bus[245]), .B(n106), .ZN(
        n107) );
  AOI21D1BWP30P140LVT U134 ( .A1(n3), .A2(i_data_bus[21]), .B(n107), .ZN(n110)
         );
  AOI22D1BWP30P140LVT U135 ( .A1(n208), .A2(i_data_bus[85]), .B1(n227), .B2(
        i_data_bus[53]), .ZN(n109) );
  AOI22D1BWP30P140LVT U136 ( .A1(n219), .A2(i_data_bus[117]), .B1(n4), .B2(
        i_data_bus[149]), .ZN(n108) );
  ND3D1BWP30P140LVT U137 ( .A1(n110), .A2(n109), .A3(n108), .ZN(N390) );
  AOI22D1BWP30P140LVT U138 ( .A1(n205), .A2(i_data_bus[214]), .B1(n2), .B2(
        i_data_bus[182]), .ZN(n111) );
  IOA21D1BWP30P140LVT U139 ( .A1(n18), .A2(i_data_bus[246]), .B(n111), .ZN(
        n112) );
  AOI21D1BWP30P140LVT U140 ( .A1(n3), .A2(i_data_bus[22]), .B(n112), .ZN(n115)
         );
  AOI22D1BWP30P140LVT U141 ( .A1(n208), .A2(i_data_bus[86]), .B1(n227), .B2(
        i_data_bus[54]), .ZN(n114) );
  AOI22D1BWP30P140LVT U142 ( .A1(n219), .A2(i_data_bus[118]), .B1(n4), .B2(
        i_data_bus[150]), .ZN(n113) );
  ND3D1BWP30P140LVT U143 ( .A1(n115), .A2(n114), .A3(n113), .ZN(N391) );
  AOI22D1BWP30P140LVT U144 ( .A1(n205), .A2(i_data_bus[215]), .B1(n2), .B2(
        i_data_bus[183]), .ZN(n116) );
  IOA21D1BWP30P140LVT U145 ( .A1(n18), .A2(i_data_bus[247]), .B(n116), .ZN(
        n117) );
  AOI21D1BWP30P140LVT U146 ( .A1(n201), .A2(i_data_bus[23]), .B(n117), .ZN(
        n120) );
  AOI22D1BWP30P140LVT U147 ( .A1(n208), .A2(i_data_bus[87]), .B1(n227), .B2(
        i_data_bus[55]), .ZN(n119) );
  AOI22D1BWP30P140LVT U148 ( .A1(n219), .A2(i_data_bus[119]), .B1(n4), .B2(
        i_data_bus[151]), .ZN(n118) );
  ND3D1BWP30P140LVT U149 ( .A1(n120), .A2(n119), .A3(n118), .ZN(N392) );
  AOI22D1BWP30P140LVT U150 ( .A1(n205), .A2(i_data_bus[216]), .B1(n2), .B2(
        i_data_bus[184]), .ZN(n121) );
  IOA21D1BWP30P140LVT U151 ( .A1(n18), .A2(i_data_bus[248]), .B(n121), .ZN(
        n122) );
  AOI21D1BWP30P140LVT U152 ( .A1(n3), .A2(i_data_bus[24]), .B(n122), .ZN(n125)
         );
  AOI22D1BWP30P140LVT U153 ( .A1(n208), .A2(i_data_bus[88]), .B1(n227), .B2(
        i_data_bus[56]), .ZN(n124) );
  AOI22D1BWP30P140LVT U154 ( .A1(n219), .A2(i_data_bus[120]), .B1(n4), .B2(
        i_data_bus[152]), .ZN(n123) );
  ND3D1BWP30P140LVT U155 ( .A1(n125), .A2(n124), .A3(n123), .ZN(N393) );
  AOI22D1BWP30P140LVT U156 ( .A1(n205), .A2(i_data_bus[210]), .B1(n2), .B2(
        i_data_bus[178]), .ZN(n126) );
  IOA21D1BWP30P140LVT U157 ( .A1(n18), .A2(i_data_bus[242]), .B(n126), .ZN(
        n127) );
  AOI21D1BWP30P140LVT U158 ( .A1(n3), .A2(i_data_bus[18]), .B(n127), .ZN(n130)
         );
  AOI22D1BWP30P140LVT U159 ( .A1(n208), .A2(i_data_bus[82]), .B1(n227), .B2(
        i_data_bus[50]), .ZN(n129) );
  AOI22D1BWP30P140LVT U160 ( .A1(n219), .A2(i_data_bus[114]), .B1(n4), .B2(
        i_data_bus[146]), .ZN(n128) );
  ND3D1BWP30P140LVT U161 ( .A1(n130), .A2(n129), .A3(n128), .ZN(N387) );
  AOI22D1BWP30P140LVT U162 ( .A1(n205), .A2(i_data_bus[211]), .B1(n2), .B2(
        i_data_bus[179]), .ZN(n131) );
  IOA21D1BWP30P140LVT U163 ( .A1(n18), .A2(i_data_bus[243]), .B(n131), .ZN(
        n132) );
  AOI21D1BWP30P140LVT U164 ( .A1(n201), .A2(i_data_bus[19]), .B(n132), .ZN(
        n135) );
  AOI22D1BWP30P140LVT U165 ( .A1(n208), .A2(i_data_bus[83]), .B1(n227), .B2(
        i_data_bus[51]), .ZN(n134) );
  AOI22D1BWP30P140LVT U166 ( .A1(n219), .A2(i_data_bus[115]), .B1(n4), .B2(
        i_data_bus[147]), .ZN(n133) );
  ND3D1BWP30P140LVT U167 ( .A1(n135), .A2(n134), .A3(n133), .ZN(N388) );
  AOI22D1BWP30P140LVT U168 ( .A1(n205), .A2(i_data_bus[209]), .B1(n2), .B2(
        i_data_bus[177]), .ZN(n136) );
  IOA21D1BWP30P140LVT U169 ( .A1(n18), .A2(i_data_bus[241]), .B(n136), .ZN(
        n137) );
  AOI21D1BWP30P140LVT U170 ( .A1(n3), .A2(i_data_bus[17]), .B(n137), .ZN(n140)
         );
  AOI22D1BWP30P140LVT U171 ( .A1(n208), .A2(i_data_bus[81]), .B1(n227), .B2(
        i_data_bus[49]), .ZN(n139) );
  AOI22D1BWP30P140LVT U172 ( .A1(n219), .A2(i_data_bus[113]), .B1(n4), .B2(
        i_data_bus[145]), .ZN(n138) );
  ND3D1BWP30P140LVT U173 ( .A1(n140), .A2(n139), .A3(n138), .ZN(N386) );
  INVD1BWP30P140LVT U174 ( .I(i_data_bus[173]), .ZN(n141) );
  MAOI22D1BWP30P140LVT U175 ( .A1(n212), .A2(i_data_bus[205]), .B1(n142), .B2(
        n141), .ZN(n143) );
  IOA21D1BWP30P140LVT U176 ( .A1(n18), .A2(i_data_bus[237]), .B(n143), .ZN(
        n144) );
  AOI21D1BWP30P140LVT U177 ( .A1(n3), .A2(i_data_bus[13]), .B(n144), .ZN(n147)
         );
  AOI22D1BWP30P140LVT U178 ( .A1(n208), .A2(i_data_bus[77]), .B1(n227), .B2(
        i_data_bus[45]), .ZN(n146) );
  AOI22D1BWP30P140LVT U179 ( .A1(n228), .A2(i_data_bus[109]), .B1(n4), .B2(
        i_data_bus[141]), .ZN(n145) );
  ND3D1BWP30P140LVT U180 ( .A1(n147), .A2(n146), .A3(n145), .ZN(N382) );
  AOI22D1BWP30P140LVT U181 ( .A1(n205), .A2(i_data_bus[212]), .B1(n2), .B2(
        i_data_bus[180]), .ZN(n148) );
  IOA21D1BWP30P140LVT U182 ( .A1(n18), .A2(i_data_bus[244]), .B(n148), .ZN(
        n149) );
  AOI21D1BWP30P140LVT U183 ( .A1(n201), .A2(i_data_bus[20]), .B(n149), .ZN(
        n152) );
  AOI22D1BWP30P140LVT U184 ( .A1(n208), .A2(i_data_bus[84]), .B1(n227), .B2(
        i_data_bus[52]), .ZN(n151) );
  AOI22D1BWP30P140LVT U185 ( .A1(n219), .A2(i_data_bus[116]), .B1(n4), .B2(
        i_data_bus[148]), .ZN(n150) );
  ND3D1BWP30P140LVT U186 ( .A1(n152), .A2(n151), .A3(n150), .ZN(N389) );
  INVD1BWP30P140LVT U187 ( .I(i_data_bus[193]), .ZN(n153) );
  MAOI22D1BWP30P140LVT U188 ( .A1(n2), .A2(i_data_bus[161]), .B1(n224), .B2(
        n153), .ZN(n154) );
  IOA21D1BWP30P140LVT U189 ( .A1(n18), .A2(i_data_bus[225]), .B(n154), .ZN(
        n155) );
  AOI21D1BWP30P140LVT U190 ( .A1(n201), .A2(i_data_bus[1]), .B(n155), .ZN(n158) );
  AOI22D1BWP30P140LVT U191 ( .A1(n208), .A2(i_data_bus[65]), .B1(n227), .B2(
        i_data_bus[33]), .ZN(n157) );
  AOI22D1BWP30P140LVT U192 ( .A1(n228), .A2(i_data_bus[97]), .B1(n4), .B2(
        i_data_bus[129]), .ZN(n156) );
  ND3D1BWP30P140LVT U193 ( .A1(n158), .A2(n157), .A3(n156), .ZN(N370) );
  INVD1BWP30P140LVT U194 ( .I(i_data_bus[194]), .ZN(n159) );
  MAOI22D1BWP30P140LVT U195 ( .A1(n2), .A2(i_data_bus[162]), .B1(n224), .B2(
        n159), .ZN(n160) );
  IOA21D1BWP30P140LVT U196 ( .A1(n18), .A2(i_data_bus[226]), .B(n160), .ZN(
        n161) );
  AOI21D1BWP30P140LVT U197 ( .A1(n3), .A2(i_data_bus[2]), .B(n161), .ZN(n164)
         );
  AOI22D1BWP30P140LVT U198 ( .A1(n208), .A2(i_data_bus[66]), .B1(n227), .B2(
        i_data_bus[34]), .ZN(n163) );
  AOI22D1BWP30P140LVT U199 ( .A1(n228), .A2(i_data_bus[98]), .B1(n4), .B2(
        i_data_bus[130]), .ZN(n162) );
  ND3D1BWP30P140LVT U200 ( .A1(n164), .A2(n163), .A3(n162), .ZN(N371) );
  INVD1BWP30P140LVT U201 ( .I(i_data_bus[195]), .ZN(n165) );
  MAOI22D1BWP30P140LVT U202 ( .A1(n2), .A2(i_data_bus[163]), .B1(n224), .B2(
        n165), .ZN(n166) );
  IOA21D1BWP30P140LVT U203 ( .A1(n18), .A2(i_data_bus[227]), .B(n166), .ZN(
        n167) );
  AOI21D1BWP30P140LVT U204 ( .A1(n3), .A2(i_data_bus[3]), .B(n167), .ZN(n170)
         );
  AOI22D1BWP30P140LVT U205 ( .A1(n208), .A2(i_data_bus[67]), .B1(n227), .B2(
        i_data_bus[35]), .ZN(n169) );
  AOI22D1BWP30P140LVT U206 ( .A1(n228), .A2(i_data_bus[99]), .B1(n4), .B2(
        i_data_bus[131]), .ZN(n168) );
  ND3D1BWP30P140LVT U207 ( .A1(n170), .A2(n169), .A3(n168), .ZN(N372) );
  AOI22D1BWP30P140LVT U208 ( .A1(n205), .A2(i_data_bus[218]), .B1(n2), .B2(
        i_data_bus[186]), .ZN(n171) );
  IOA21D1BWP30P140LVT U209 ( .A1(n18), .A2(i_data_bus[250]), .B(n171), .ZN(
        n172) );
  AOI21D1BWP30P140LVT U210 ( .A1(n3), .A2(i_data_bus[26]), .B(n172), .ZN(n175)
         );
  AOI22D1BWP30P140LVT U211 ( .A1(n208), .A2(i_data_bus[90]), .B1(n227), .B2(
        i_data_bus[58]), .ZN(n174) );
  AOI22D1BWP30P140LVT U212 ( .A1(n219), .A2(i_data_bus[122]), .B1(n4), .B2(
        i_data_bus[154]), .ZN(n173) );
  ND3D1BWP30P140LVT U213 ( .A1(n175), .A2(n174), .A3(n173), .ZN(N395) );
  AOI22D1BWP30P140LVT U214 ( .A1(n205), .A2(i_data_bus[219]), .B1(n2), .B2(
        i_data_bus[187]), .ZN(n176) );
  IOA21D1BWP30P140LVT U215 ( .A1(n18), .A2(i_data_bus[251]), .B(n176), .ZN(
        n177) );
  AOI21D1BWP30P140LVT U216 ( .A1(n3), .A2(i_data_bus[27]), .B(n177), .ZN(n180)
         );
  AOI22D1BWP30P140LVT U217 ( .A1(n208), .A2(i_data_bus[91]), .B1(n227), .B2(
        i_data_bus[59]), .ZN(n179) );
  AOI22D1BWP30P140LVT U218 ( .A1(n219), .A2(i_data_bus[123]), .B1(n4), .B2(
        i_data_bus[155]), .ZN(n178) );
  ND3D1BWP30P140LVT U219 ( .A1(n180), .A2(n179), .A3(n178), .ZN(N396) );
  INVD1BWP30P140LVT U220 ( .I(i_data_bus[221]), .ZN(n181) );
  MAOI22D1BWP30P140LVT U221 ( .A1(n2), .A2(i_data_bus[189]), .B1(n224), .B2(
        n181), .ZN(n182) );
  IOA21D1BWP30P140LVT U222 ( .A1(n18), .A2(i_data_bus[253]), .B(n182), .ZN(
        n183) );
  AOI21D1BWP30P140LVT U223 ( .A1(n201), .A2(i_data_bus[29]), .B(n183), .ZN(
        n186) );
  AOI22D1BWP30P140LVT U224 ( .A1(n208), .A2(i_data_bus[93]), .B1(n227), .B2(
        i_data_bus[61]), .ZN(n185) );
  AOI22D1BWP30P140LVT U225 ( .A1(n219), .A2(i_data_bus[125]), .B1(n4), .B2(
        i_data_bus[157]), .ZN(n184) );
  ND3D1BWP30P140LVT U226 ( .A1(n186), .A2(n185), .A3(n184), .ZN(N398) );
  INVD1BWP30P140LVT U227 ( .I(i_data_bus[222]), .ZN(n187) );
  MAOI22D1BWP30P140LVT U228 ( .A1(n2), .A2(i_data_bus[190]), .B1(n224), .B2(
        n187), .ZN(n188) );
  IOA21D1BWP30P140LVT U229 ( .A1(n18), .A2(i_data_bus[254]), .B(n188), .ZN(
        n189) );
  AOI21D1BWP30P140LVT U230 ( .A1(n3), .A2(i_data_bus[30]), .B(n189), .ZN(n192)
         );
  AOI22D1BWP30P140LVT U231 ( .A1(n219), .A2(i_data_bus[126]), .B1(n4), .B2(
        i_data_bus[158]), .ZN(n190) );
  ND3D1BWP30P140LVT U232 ( .A1(n192), .A2(n191), .A3(n190), .ZN(N399) );
  INVD1BWP30P140LVT U233 ( .I(i_data_bus[223]), .ZN(n193) );
  MAOI22D1BWP30P140LVT U234 ( .A1(n2), .A2(i_data_bus[191]), .B1(n224), .B2(
        n193), .ZN(n194) );
  IOA21D1BWP30P140LVT U235 ( .A1(n18), .A2(i_data_bus[255]), .B(n194), .ZN(
        n195) );
  AOI21D1BWP30P140LVT U236 ( .A1(n3), .A2(i_data_bus[31]), .B(n195), .ZN(n198)
         );
  AOI22D1BWP30P140LVT U237 ( .A1(n208), .A2(i_data_bus[95]), .B1(n227), .B2(
        i_data_bus[63]), .ZN(n197) );
  AOI22D1BWP30P140LVT U238 ( .A1(n219), .A2(i_data_bus[127]), .B1(n4), .B2(
        i_data_bus[159]), .ZN(n196) );
  ND3D1BWP30P140LVT U239 ( .A1(n198), .A2(n197), .A3(n196), .ZN(N400) );
  AOI22D1BWP30P140LVT U240 ( .A1(n205), .A2(i_data_bus[217]), .B1(n2), .B2(
        i_data_bus[185]), .ZN(n199) );
  IOA21D1BWP30P140LVT U241 ( .A1(n18), .A2(i_data_bus[249]), .B(n199), .ZN(
        n200) );
  AOI21D1BWP30P140LVT U242 ( .A1(n201), .A2(i_data_bus[25]), .B(n200), .ZN(
        n204) );
  AOI22D1BWP30P140LVT U243 ( .A1(n208), .A2(i_data_bus[89]), .B1(n227), .B2(
        i_data_bus[57]), .ZN(n203) );
  AOI22D1BWP30P140LVT U244 ( .A1(n228), .A2(i_data_bus[121]), .B1(n4), .B2(
        i_data_bus[153]), .ZN(n202) );
  ND3D1BWP30P140LVT U245 ( .A1(n204), .A2(n203), .A3(n202), .ZN(N394) );
  AOI22D1BWP30P140LVT U246 ( .A1(n205), .A2(i_data_bus[220]), .B1(n2), .B2(
        i_data_bus[188]), .ZN(n206) );
  IOA21D1BWP30P140LVT U247 ( .A1(n18), .A2(i_data_bus[252]), .B(n206), .ZN(
        n207) );
  AOI21D1BWP30P140LVT U248 ( .A1(n3), .A2(i_data_bus[28]), .B(n207), .ZN(n211)
         );
  AOI22D1BWP30P140LVT U249 ( .A1(n208), .A2(i_data_bus[92]), .B1(n227), .B2(
        i_data_bus[60]), .ZN(n210) );
  AOI22D1BWP30P140LVT U250 ( .A1(n219), .A2(i_data_bus[124]), .B1(n4), .B2(
        i_data_bus[156]), .ZN(n209) );
  ND3D1BWP30P140LVT U251 ( .A1(n211), .A2(n210), .A3(n209), .ZN(N397) );
  AOI22D1BWP30P140LVT U252 ( .A1(n212), .A2(i_data_bus[207]), .B1(n2), .B2(
        i_data_bus[175]), .ZN(n213) );
  IOA21D1BWP30P140LVT U253 ( .A1(n18), .A2(i_data_bus[239]), .B(n213), .ZN(
        n214) );
  AOI21D1BWP30P140LVT U254 ( .A1(n3), .A2(i_data_bus[15]), .B(n214), .ZN(n222)
         );
  INVD1BWP30P140LVT U255 ( .I(i_data_bus[79]), .ZN(n217) );
  INVD1BWP30P140LVT U256 ( .I(i_data_bus[47]), .ZN(n215) );
  OA22D1BWP30P140LVT U257 ( .A1(n218), .A2(n217), .B1(n216), .B2(n215), .Z(
        n221) );
  AOI22D1BWP30P140LVT U258 ( .A1(n219), .A2(i_data_bus[111]), .B1(n4), .B2(
        i_data_bus[143]), .ZN(n220) );
  ND3D1BWP30P140LVT U259 ( .A1(n222), .A2(n221), .A3(n220), .ZN(N384) );
  INVD1BWP30P140LVT U260 ( .I(i_data_bus[208]), .ZN(n223) );
  MAOI22D1BWP30P140LVT U261 ( .A1(n2), .A2(i_data_bus[176]), .B1(n224), .B2(
        n223), .ZN(n225) );
  IOA21D1BWP30P140LVT U262 ( .A1(n18), .A2(i_data_bus[240]), .B(n225), .ZN(
        n226) );
  AOI21D1BWP30P140LVT U263 ( .A1(n3), .A2(i_data_bus[16]), .B(n226), .ZN(n231)
         );
  AOI22D1BWP30P140LVT U264 ( .A1(n208), .A2(i_data_bus[80]), .B1(n227), .B2(
        i_data_bus[48]), .ZN(n230) );
  AOI22D1BWP30P140LVT U265 ( .A1(n228), .A2(i_data_bus[112]), .B1(n4), .B2(
        i_data_bus[144]), .ZN(n229) );
  ND3D1BWP30P140LVT U266 ( .A1(n231), .A2(n230), .A3(n229), .ZN(N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_7 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  AOI21D1BWP30P140LVT U3 ( .A1(n3), .A2(i_data_bus[17]), .B(n142), .ZN(n145)
         );
  INVD6BWP30P140LVT U4 ( .I(n209), .ZN(n1) );
  OR2D1BWP30P140LVT U5 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n32) );
  CKND2D3BWP30P140LVT U6 ( .A1(n15), .A2(n14), .ZN(n22) );
  INVD6BWP30P140LVT U7 ( .I(n225), .ZN(n2) );
  INVD3BWP30P140LVT U8 ( .I(n50), .ZN(n3) );
  ND2OPTIBD1BWP30P140LVT U9 ( .A1(n42), .A2(n10), .ZN(n50) );
  ND2OPTIBD2BWP30P140LVT U10 ( .A1(n7), .A2(n6), .ZN(n27) );
  INVD1BWP30P140LVT U11 ( .I(i_valid[6]), .ZN(n17) );
  NR2D1BWP30P140LVT U12 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n28) );
  NR2D1BWP30P140LVT U13 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .ZN(n4) );
  NR2OPTPAD1BWP30P140LVT U14 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .ZN(n7) );
  INR2D1BWP30P140LVT U15 ( .A1(i_en), .B1(rst), .ZN(n5) );
  INR2D1BWP30P140LVT U16 ( .A1(n5), .B1(i_cmd[6]), .ZN(n6) );
  NR3D1P5BWP30P140LVT U17 ( .A1(n32), .A2(n27), .A3(i_cmd[1]), .ZN(n42) );
  INR2D1BWP30P140LVT U18 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n8) );
  INVD1BWP30P140LVT U19 ( .I(n8), .ZN(n9) );
  INR2D1BWP30P140LVT U20 ( .A1(i_cmd[0]), .B1(n9), .ZN(n10) );
  ND2OPTIBD1BWP30P140LVT U21 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n11) );
  NR3D0P7BWP30P140LVT U22 ( .A1(n11), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n16)
         );
  NR3D1P5BWP30P140LVT U23 ( .A1(i_cmd[2]), .A2(i_cmd[0]), .A3(i_cmd[3]), .ZN(
        n15) );
  INR2D1BWP30P140LVT U24 ( .A1(i_en), .B1(rst), .ZN(n12) );
  INVD1BWP30P140LVT U25 ( .I(n12), .ZN(n13) );
  NR3D1P5BWP30P140LVT U26 ( .A1(i_cmd[1]), .A2(i_cmd[4]), .A3(n13), .ZN(n14)
         );
  INR2D2BWP30P140LVT U27 ( .A1(n16), .B1(n22), .ZN(n228) );
  INVD1BWP30P140LVT U28 ( .I(i_cmd[6]), .ZN(n18) );
  NR4D1BWP30P140LVT U29 ( .A1(n18), .A2(n17), .A3(i_cmd[5]), .A4(i_cmd[7]), 
        .ZN(n19) );
  INR2D2BWP30P140LVT U30 ( .A1(n19), .B1(n22), .ZN(n20) );
  INVD3BWP30P140LVT U31 ( .I(n20), .ZN(n225) );
  INVD1BWP30P140LVT U32 ( .I(i_cmd[5]), .ZN(n21) );
  INR4D1BWP30P140LVT U33 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n21), .ZN(n23) );
  INR2D2BWP30P140LVT U34 ( .A1(n23), .B1(n22), .ZN(n24) );
  INVD2BWP30P140LVT U35 ( .I(n24), .ZN(n180) );
  INVD3BWP30P140LVT U36 ( .I(n180), .ZN(n226) );
  AOI22D1BWP30P140LVT U37 ( .A1(n2), .A2(i_data_bus[206]), .B1(n226), .B2(
        i_data_bus[174]), .ZN(n25) );
  IOA21D1BWP30P140LVT U38 ( .A1(n228), .A2(i_data_bus[238]), .B(n25), .ZN(n26)
         );
  AOI21OPTREPBD1BWP30P140LVT U39 ( .A1(n3), .A2(i_data_bus[14]), .B(n26), .ZN(
        n45) );
  INR2D2BWP30P140LVT U40 ( .A1(n28), .B1(n27), .ZN(n38) );
  INVD1BWP30P140LVT U41 ( .I(i_cmd[1]), .ZN(n29) );
  INVD1BWP30P140LVT U42 ( .I(i_cmd[3]), .ZN(n36) );
  ND4D1BWP30P140LVT U43 ( .A1(n29), .A2(n36), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n30) );
  INR2D1BWP30P140LVT U44 ( .A1(n38), .B1(n30), .ZN(n31) );
  INVD2BWP30P140LVT U45 ( .I(n31), .ZN(n211) );
  INVD2BWP30P140LVT U46 ( .I(n211), .ZN(n219) );
  INVD1BWP30P140LVT U47 ( .I(n32), .ZN(n33) );
  ND3D1BWP30P140LVT U48 ( .A1(n33), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n34)
         );
  INR2D1BWP30P140LVT U49 ( .A1(n38), .B1(n34), .ZN(n35) );
  INVD2BWP30P140LVT U50 ( .I(n35), .ZN(n209) );
  AOI22D1BWP30P140LVT U51 ( .A1(n219), .A2(i_data_bus[78]), .B1(n1), .B2(
        i_data_bus[46]), .ZN(n44) );
  ND3D1BWP30P140LVT U52 ( .A1(n4), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n37) );
  INR2D1BWP30P140LVT U53 ( .A1(n38), .B1(n37), .ZN(n39) );
  INVD2BWP30P140LVT U54 ( .I(n39), .ZN(n56) );
  INVD2BWP30P140LVT U55 ( .I(n56), .ZN(n220) );
  IND3D1BWP30P140LVT U56 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n40) );
  INVD1BWP30P140LVT U57 ( .I(n40), .ZN(n41) );
  ND2OPTIBD2BWP30P140LVT U58 ( .A1(n42), .A2(n41), .ZN(n57) );
  INVD2BWP30P140LVT U59 ( .I(n57), .ZN(n231) );
  AOI22D1BWP30P140LVT U60 ( .A1(n220), .A2(i_data_bus[110]), .B1(n231), .B2(
        i_data_bus[142]), .ZN(n43) );
  ND3D1BWP30P140LVT U61 ( .A1(n45), .A2(n44), .A3(n43), .ZN(N383) );
  NR4D0BWP30P140LVT U62 ( .A1(n3), .A2(n228), .A3(n2), .A4(n226), .ZN(n48) );
  INVD1BWP30P140LVT U63 ( .I(n211), .ZN(n230) );
  NR2D1BWP30P140LVT U64 ( .A1(n230), .A2(n1), .ZN(n47) );
  INVD1BWP30P140LVT U65 ( .I(n56), .ZN(n232) );
  NR2D1BWP30P140LVT U66 ( .A1(n232), .A2(n231), .ZN(n46) );
  ND3D1BWP30P140LVT U67 ( .A1(n48), .A2(n47), .A3(n46), .ZN(N402) );
  INVD1BWP30P140LVT U68 ( .I(n228), .ZN(n55) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[224]), .ZN(n54) );
  INVD3BWP30P140LVT U70 ( .I(n180), .ZN(n216) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[192]), .ZN(n49) );
  MAOI22D1BWP30P140LVT U72 ( .A1(n216), .A2(i_data_bus[160]), .B1(n225), .B2(
        n49), .ZN(n53) );
  INR2D1BWP30P140LVT U73 ( .A1(i_data_bus[0]), .B1(n50), .ZN(n51) );
  INVD1BWP30P140LVT U74 ( .I(n51), .ZN(n52) );
  OA211D1BWP30P140LVT U75 ( .A1(n55), .A2(n54), .B(n53), .C(n52), .Z(n60) );
  INVD2BWP30P140LVT U76 ( .I(n211), .ZN(n161) );
  AOI22D1BWP30P140LVT U77 ( .A1(n161), .A2(i_data_bus[64]), .B1(n1), .B2(
        i_data_bus[32]), .ZN(n59) );
  INVD2BWP30P140LVT U78 ( .I(n56), .ZN(n163) );
  INVD2BWP30P140LVT U79 ( .I(n57), .ZN(n162) );
  AOI22D1BWP30P140LVT U80 ( .A1(n163), .A2(i_data_bus[96]), .B1(n162), .B2(
        i_data_bus[128]), .ZN(n58) );
  ND3D1BWP30P140LVT U81 ( .A1(n60), .A2(n59), .A3(n58), .ZN(N369) );
  AOI22D1BWP30P140LVT U82 ( .A1(n2), .A2(i_data_bus[203]), .B1(n226), .B2(
        i_data_bus[171]), .ZN(n61) );
  IOA21D1BWP30P140LVT U83 ( .A1(n228), .A2(i_data_bus[235]), .B(n61), .ZN(n62)
         );
  AOI21D1BWP30P140LVT U84 ( .A1(n3), .A2(i_data_bus[11]), .B(n62), .ZN(n65) );
  AOI22D1BWP30P140LVT U85 ( .A1(n161), .A2(i_data_bus[75]), .B1(n1), .B2(
        i_data_bus[43]), .ZN(n64) );
  AOI22D1BWP30P140LVT U86 ( .A1(n163), .A2(i_data_bus[107]), .B1(n162), .B2(
        i_data_bus[139]), .ZN(n63) );
  ND3D1BWP30P140LVT U87 ( .A1(n65), .A2(n64), .A3(n63), .ZN(N380) );
  AOI22D1BWP30P140LVT U88 ( .A1(n2), .A2(i_data_bus[200]), .B1(n226), .B2(
        i_data_bus[168]), .ZN(n66) );
  IOA21D1BWP30P140LVT U89 ( .A1(n228), .A2(i_data_bus[232]), .B(n66), .ZN(n67)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n3), .A2(i_data_bus[8]), .B(n67), .ZN(n70) );
  AOI22D1BWP30P140LVT U91 ( .A1(n161), .A2(i_data_bus[72]), .B1(n1), .B2(
        i_data_bus[40]), .ZN(n69) );
  AOI22D1BWP30P140LVT U92 ( .A1(n163), .A2(i_data_bus[104]), .B1(n162), .B2(
        i_data_bus[136]), .ZN(n68) );
  ND3D1BWP30P140LVT U93 ( .A1(n70), .A2(n69), .A3(n68), .ZN(N377) );
  AOI22D1BWP30P140LVT U94 ( .A1(n2), .A2(i_data_bus[202]), .B1(n226), .B2(
        i_data_bus[170]), .ZN(n71) );
  IOA21D1BWP30P140LVT U95 ( .A1(n228), .A2(i_data_bus[234]), .B(n71), .ZN(n72)
         );
  AOI21D1BWP30P140LVT U96 ( .A1(n3), .A2(i_data_bus[10]), .B(n72), .ZN(n75) );
  AOI22D1BWP30P140LVT U97 ( .A1(n161), .A2(i_data_bus[74]), .B1(n1), .B2(
        i_data_bus[42]), .ZN(n74) );
  AOI22D1BWP30P140LVT U98 ( .A1(n163), .A2(i_data_bus[106]), .B1(n162), .B2(
        i_data_bus[138]), .ZN(n73) );
  ND3D1BWP30P140LVT U99 ( .A1(n75), .A2(n74), .A3(n73), .ZN(N379) );
  AOI22D1BWP30P140LVT U100 ( .A1(n2), .A2(i_data_bus[199]), .B1(n226), .B2(
        i_data_bus[167]), .ZN(n76) );
  IOA21D1BWP30P140LVT U101 ( .A1(n228), .A2(i_data_bus[231]), .B(n76), .ZN(n77) );
  AOI21D1BWP30P140LVT U102 ( .A1(n3), .A2(i_data_bus[7]), .B(n77), .ZN(n80) );
  AOI22D1BWP30P140LVT U103 ( .A1(n161), .A2(i_data_bus[71]), .B1(n1), .B2(
        i_data_bus[39]), .ZN(n79) );
  AOI22D1BWP30P140LVT U104 ( .A1(n163), .A2(i_data_bus[103]), .B1(n162), .B2(
        i_data_bus[135]), .ZN(n78) );
  ND3D1BWP30P140LVT U105 ( .A1(n80), .A2(n79), .A3(n78), .ZN(N376) );
  AOI22D1BWP30P140LVT U106 ( .A1(n2), .A2(i_data_bus[198]), .B1(n226), .B2(
        i_data_bus[166]), .ZN(n81) );
  IOA21D1BWP30P140LVT U107 ( .A1(n228), .A2(i_data_bus[230]), .B(n81), .ZN(n82) );
  AOI21D1BWP30P140LVT U108 ( .A1(n3), .A2(i_data_bus[6]), .B(n82), .ZN(n85) );
  AOI22D1BWP30P140LVT U109 ( .A1(n161), .A2(i_data_bus[70]), .B1(n1), .B2(
        i_data_bus[38]), .ZN(n84) );
  AOI22D1BWP30P140LVT U110 ( .A1(n163), .A2(i_data_bus[102]), .B1(n162), .B2(
        i_data_bus[134]), .ZN(n83) );
  ND3D1BWP30P140LVT U111 ( .A1(n85), .A2(n84), .A3(n83), .ZN(N375) );
  AOI22D1BWP30P140LVT U112 ( .A1(n2), .A2(i_data_bus[204]), .B1(n226), .B2(
        i_data_bus[172]), .ZN(n86) );
  IOA21D1BWP30P140LVT U113 ( .A1(n228), .A2(i_data_bus[236]), .B(n86), .ZN(n87) );
  AOI21D1BWP30P140LVT U114 ( .A1(n3), .A2(i_data_bus[12]), .B(n87), .ZN(n90)
         );
  AOI22D1BWP30P140LVT U115 ( .A1(n161), .A2(i_data_bus[76]), .B1(n1), .B2(
        i_data_bus[44]), .ZN(n89) );
  AOI22D1BWP30P140LVT U116 ( .A1(n163), .A2(i_data_bus[108]), .B1(n162), .B2(
        i_data_bus[140]), .ZN(n88) );
  ND3D1BWP30P140LVT U117 ( .A1(n90), .A2(n89), .A3(n88), .ZN(N381) );
  AOI22D1BWP30P140LVT U118 ( .A1(n2), .A2(i_data_bus[197]), .B1(n226), .B2(
        i_data_bus[165]), .ZN(n91) );
  IOA21D1BWP30P140LVT U119 ( .A1(n228), .A2(i_data_bus[229]), .B(n91), .ZN(n92) );
  AOI21D1BWP30P140LVT U120 ( .A1(n3), .A2(i_data_bus[5]), .B(n92), .ZN(n95) );
  AOI22D1BWP30P140LVT U121 ( .A1(n161), .A2(i_data_bus[69]), .B1(n1), .B2(
        i_data_bus[37]), .ZN(n94) );
  AOI22D1BWP30P140LVT U122 ( .A1(n163), .A2(i_data_bus[101]), .B1(n162), .B2(
        i_data_bus[133]), .ZN(n93) );
  ND3D1BWP30P140LVT U123 ( .A1(n95), .A2(n94), .A3(n93), .ZN(N374) );
  AOI22D1BWP30P140LVT U124 ( .A1(n2), .A2(i_data_bus[196]), .B1(n226), .B2(
        i_data_bus[164]), .ZN(n96) );
  IOA21D1BWP30P140LVT U125 ( .A1(n228), .A2(i_data_bus[228]), .B(n96), .ZN(n97) );
  AOI21D1BWP30P140LVT U126 ( .A1(n3), .A2(i_data_bus[4]), .B(n97), .ZN(n100)
         );
  AOI22D1BWP30P140LVT U127 ( .A1(n161), .A2(i_data_bus[68]), .B1(n1), .B2(
        i_data_bus[36]), .ZN(n99) );
  AOI22D1BWP30P140LVT U128 ( .A1(n163), .A2(i_data_bus[100]), .B1(n162), .B2(
        i_data_bus[132]), .ZN(n98) );
  ND3D1BWP30P140LVT U129 ( .A1(n100), .A2(n99), .A3(n98), .ZN(N373) );
  AOI22D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[201]), .B1(n226), .B2(
        i_data_bus[169]), .ZN(n101) );
  IOA21D1BWP30P140LVT U131 ( .A1(n228), .A2(i_data_bus[233]), .B(n101), .ZN(
        n102) );
  AOI21D1BWP30P140LVT U132 ( .A1(n3), .A2(i_data_bus[9]), .B(n102), .ZN(n105)
         );
  AOI22D1BWP30P140LVT U133 ( .A1(n161), .A2(i_data_bus[73]), .B1(n1), .B2(
        i_data_bus[41]), .ZN(n104) );
  AOI22D1BWP30P140LVT U134 ( .A1(n163), .A2(i_data_bus[105]), .B1(n162), .B2(
        i_data_bus[137]), .ZN(n103) );
  ND3D1BWP30P140LVT U135 ( .A1(n105), .A2(n104), .A3(n103), .ZN(N378) );
  AOI22D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[214]), .B1(n216), .B2(
        i_data_bus[182]), .ZN(n106) );
  IOA21D1BWP30P140LVT U137 ( .A1(n228), .A2(i_data_bus[246]), .B(n106), .ZN(
        n107) );
  AOI21D1BWP30P140LVT U138 ( .A1(n3), .A2(i_data_bus[22]), .B(n107), .ZN(n110)
         );
  AOI22D1BWP30P140LVT U139 ( .A1(n219), .A2(i_data_bus[86]), .B1(n1), .B2(
        i_data_bus[54]), .ZN(n109) );
  AOI22D1BWP30P140LVT U140 ( .A1(n220), .A2(i_data_bus[118]), .B1(n231), .B2(
        i_data_bus[150]), .ZN(n108) );
  ND3D1BWP30P140LVT U141 ( .A1(n110), .A2(n109), .A3(n108), .ZN(N391) );
  AOI22D1BWP30P140LVT U142 ( .A1(n2), .A2(i_data_bus[210]), .B1(n216), .B2(
        i_data_bus[178]), .ZN(n111) );
  IOA21D1BWP30P140LVT U143 ( .A1(n228), .A2(i_data_bus[242]), .B(n111), .ZN(
        n112) );
  AOI21OPTREPBD1BWP30P140LVT U144 ( .A1(n3), .A2(i_data_bus[18]), .B(n112), 
        .ZN(n115) );
  AOI22D1BWP30P140LVT U145 ( .A1(n219), .A2(i_data_bus[82]), .B1(n1), .B2(
        i_data_bus[50]), .ZN(n114) );
  AOI22D1BWP30P140LVT U146 ( .A1(n220), .A2(i_data_bus[114]), .B1(n231), .B2(
        i_data_bus[146]), .ZN(n113) );
  ND3D1BWP30P140LVT U147 ( .A1(n115), .A2(n114), .A3(n113), .ZN(N387) );
  AOI22D1BWP30P140LVT U148 ( .A1(n2), .A2(i_data_bus[215]), .B1(n216), .B2(
        i_data_bus[183]), .ZN(n116) );
  IOA21D1BWP30P140LVT U149 ( .A1(n228), .A2(i_data_bus[247]), .B(n116), .ZN(
        n117) );
  AOI21D1BWP30P140LVT U150 ( .A1(n3), .A2(i_data_bus[23]), .B(n117), .ZN(n120)
         );
  AOI22D1BWP30P140LVT U151 ( .A1(n219), .A2(i_data_bus[87]), .B1(n1), .B2(
        i_data_bus[55]), .ZN(n119) );
  AOI22D1BWP30P140LVT U152 ( .A1(n220), .A2(i_data_bus[119]), .B1(n231), .B2(
        i_data_bus[151]), .ZN(n118) );
  ND3D1BWP30P140LVT U153 ( .A1(n120), .A2(n119), .A3(n118), .ZN(N392) );
  AOI22D1BWP30P140LVT U154 ( .A1(n2), .A2(i_data_bus[216]), .B1(n216), .B2(
        i_data_bus[184]), .ZN(n121) );
  IOA21D1BWP30P140LVT U155 ( .A1(n228), .A2(i_data_bus[248]), .B(n121), .ZN(
        n122) );
  AOI21D1BWP30P140LVT U156 ( .A1(n3), .A2(i_data_bus[24]), .B(n122), .ZN(n125)
         );
  AOI22D1BWP30P140LVT U157 ( .A1(n219), .A2(i_data_bus[88]), .B1(n1), .B2(
        i_data_bus[56]), .ZN(n124) );
  AOI22D1BWP30P140LVT U158 ( .A1(n220), .A2(i_data_bus[120]), .B1(n231), .B2(
        i_data_bus[152]), .ZN(n123) );
  ND3D1BWP30P140LVT U159 ( .A1(n125), .A2(n124), .A3(n123), .ZN(N393) );
  AOI22D1BWP30P140LVT U160 ( .A1(n2), .A2(i_data_bus[213]), .B1(n216), .B2(
        i_data_bus[181]), .ZN(n126) );
  IOA21D1BWP30P140LVT U161 ( .A1(n228), .A2(i_data_bus[245]), .B(n126), .ZN(
        n127) );
  AOI21D1BWP30P140LVT U162 ( .A1(n3), .A2(i_data_bus[21]), .B(n127), .ZN(n130)
         );
  AOI22D1BWP30P140LVT U163 ( .A1(n219), .A2(i_data_bus[85]), .B1(n1), .B2(
        i_data_bus[53]), .ZN(n129) );
  AOI22D1BWP30P140LVT U164 ( .A1(n220), .A2(i_data_bus[117]), .B1(n231), .B2(
        i_data_bus[149]), .ZN(n128) );
  ND3D1BWP30P140LVT U165 ( .A1(n130), .A2(n129), .A3(n128), .ZN(N390) );
  AOI22D1BWP30P140LVT U166 ( .A1(n2), .A2(i_data_bus[211]), .B1(n216), .B2(
        i_data_bus[179]), .ZN(n131) );
  IOA21D1BWP30P140LVT U167 ( .A1(n228), .A2(i_data_bus[243]), .B(n131), .ZN(
        n132) );
  AOI21D1BWP30P140LVT U168 ( .A1(n3), .A2(i_data_bus[19]), .B(n132), .ZN(n135)
         );
  AOI22D1BWP30P140LVT U169 ( .A1(n219), .A2(i_data_bus[83]), .B1(n1), .B2(
        i_data_bus[51]), .ZN(n134) );
  AOI22D1BWP30P140LVT U170 ( .A1(n220), .A2(i_data_bus[115]), .B1(n231), .B2(
        i_data_bus[147]), .ZN(n133) );
  ND3D1BWP30P140LVT U171 ( .A1(n135), .A2(n134), .A3(n133), .ZN(N388) );
  AOI22D1BWP30P140LVT U172 ( .A1(n2), .A2(i_data_bus[212]), .B1(n216), .B2(
        i_data_bus[180]), .ZN(n136) );
  IOA21D1BWP30P140LVT U173 ( .A1(n228), .A2(i_data_bus[244]), .B(n136), .ZN(
        n137) );
  AOI21D1BWP30P140LVT U174 ( .A1(n3), .A2(i_data_bus[20]), .B(n137), .ZN(n140)
         );
  AOI22D1BWP30P140LVT U175 ( .A1(n219), .A2(i_data_bus[84]), .B1(n1), .B2(
        i_data_bus[52]), .ZN(n139) );
  AOI22D1BWP30P140LVT U176 ( .A1(n220), .A2(i_data_bus[116]), .B1(n231), .B2(
        i_data_bus[148]), .ZN(n138) );
  ND3D1BWP30P140LVT U177 ( .A1(n140), .A2(n139), .A3(n138), .ZN(N389) );
  AOI22D1BWP30P140LVT U178 ( .A1(n2), .A2(i_data_bus[209]), .B1(n216), .B2(
        i_data_bus[177]), .ZN(n141) );
  IOA21D1BWP30P140LVT U179 ( .A1(n228), .A2(i_data_bus[241]), .B(n141), .ZN(
        n142) );
  AOI22D1BWP30P140LVT U180 ( .A1(n219), .A2(i_data_bus[81]), .B1(n1), .B2(
        i_data_bus[49]), .ZN(n144) );
  AOI22D1BWP30P140LVT U181 ( .A1(n220), .A2(i_data_bus[113]), .B1(n231), .B2(
        i_data_bus[145]), .ZN(n143) );
  ND3D1BWP30P140LVT U182 ( .A1(n145), .A2(n144), .A3(n143), .ZN(N386) );
  INVD1BWP30P140LVT U183 ( .I(i_data_bus[195]), .ZN(n146) );
  MAOI22D1BWP30P140LVT U184 ( .A1(n226), .A2(i_data_bus[163]), .B1(n225), .B2(
        n146), .ZN(n147) );
  IOA21D1BWP30P140LVT U185 ( .A1(n228), .A2(i_data_bus[227]), .B(n147), .ZN(
        n148) );
  AOI21D1BWP30P140LVT U186 ( .A1(n3), .A2(i_data_bus[3]), .B(n148), .ZN(n151)
         );
  AOI22D1BWP30P140LVT U187 ( .A1(n161), .A2(i_data_bus[67]), .B1(n1), .B2(
        i_data_bus[35]), .ZN(n150) );
  AOI22D1BWP30P140LVT U188 ( .A1(n163), .A2(i_data_bus[99]), .B1(n162), .B2(
        i_data_bus[131]), .ZN(n149) );
  ND3D1BWP30P140LVT U189 ( .A1(n151), .A2(n150), .A3(n149), .ZN(N372) );
  INVD1BWP30P140LVT U190 ( .I(i_data_bus[194]), .ZN(n152) );
  MAOI22D1BWP30P140LVT U191 ( .A1(n226), .A2(i_data_bus[162]), .B1(n225), .B2(
        n152), .ZN(n153) );
  IOA21D1BWP30P140LVT U192 ( .A1(n228), .A2(i_data_bus[226]), .B(n153), .ZN(
        n154) );
  AOI21D1BWP30P140LVT U193 ( .A1(n3), .A2(i_data_bus[2]), .B(n154), .ZN(n157)
         );
  AOI22D1BWP30P140LVT U194 ( .A1(n161), .A2(i_data_bus[66]), .B1(n1), .B2(
        i_data_bus[34]), .ZN(n156) );
  AOI22D1BWP30P140LVT U195 ( .A1(n163), .A2(i_data_bus[98]), .B1(n162), .B2(
        i_data_bus[130]), .ZN(n155) );
  ND3D1BWP30P140LVT U196 ( .A1(n157), .A2(n156), .A3(n155), .ZN(N371) );
  INVD1BWP30P140LVT U197 ( .I(i_data_bus[193]), .ZN(n158) );
  MAOI22D1BWP30P140LVT U198 ( .A1(n226), .A2(i_data_bus[161]), .B1(n225), .B2(
        n158), .ZN(n159) );
  IOA21D1BWP30P140LVT U199 ( .A1(n228), .A2(i_data_bus[225]), .B(n159), .ZN(
        n160) );
  AOI21D1BWP30P140LVT U200 ( .A1(n3), .A2(i_data_bus[1]), .B(n160), .ZN(n166)
         );
  AOI22D1BWP30P140LVT U201 ( .A1(n161), .A2(i_data_bus[65]), .B1(n1), .B2(
        i_data_bus[33]), .ZN(n165) );
  AOI22D1BWP30P140LVT U202 ( .A1(n163), .A2(i_data_bus[97]), .B1(n162), .B2(
        i_data_bus[129]), .ZN(n164) );
  ND3D1BWP30P140LVT U203 ( .A1(n166), .A2(n165), .A3(n164), .ZN(N370) );
  INVD1BWP30P140LVT U204 ( .I(i_data_bus[221]), .ZN(n167) );
  MAOI22D1BWP30P140LVT U205 ( .A1(n226), .A2(i_data_bus[189]), .B1(n225), .B2(
        n167), .ZN(n168) );
  IOA21D1BWP30P140LVT U206 ( .A1(n228), .A2(i_data_bus[253]), .B(n168), .ZN(
        n169) );
  AOI21D1BWP30P140LVT U207 ( .A1(n3), .A2(i_data_bus[29]), .B(n169), .ZN(n172)
         );
  AOI22D1BWP30P140LVT U208 ( .A1(n230), .A2(i_data_bus[93]), .B1(n1), .B2(
        i_data_bus[61]), .ZN(n171) );
  AOI22D1BWP30P140LVT U209 ( .A1(n232), .A2(i_data_bus[125]), .B1(n231), .B2(
        i_data_bus[157]), .ZN(n170) );
  ND3D1BWP30P140LVT U210 ( .A1(n172), .A2(n171), .A3(n170), .ZN(N398) );
  INVD1BWP30P140LVT U211 ( .I(i_data_bus[222]), .ZN(n173) );
  MAOI22D1BWP30P140LVT U212 ( .A1(n226), .A2(i_data_bus[190]), .B1(n225), .B2(
        n173), .ZN(n174) );
  IOA21D1BWP30P140LVT U213 ( .A1(n228), .A2(i_data_bus[254]), .B(n174), .ZN(
        n175) );
  AOI21D1BWP30P140LVT U214 ( .A1(n3), .A2(i_data_bus[30]), .B(n175), .ZN(n178)
         );
  AOI22D1BWP30P140LVT U215 ( .A1(n230), .A2(i_data_bus[94]), .B1(n1), .B2(
        i_data_bus[62]), .ZN(n177) );
  AOI22D1BWP30P140LVT U216 ( .A1(n232), .A2(i_data_bus[126]), .B1(n231), .B2(
        i_data_bus[158]), .ZN(n176) );
  ND3D1BWP30P140LVT U217 ( .A1(n178), .A2(n177), .A3(n176), .ZN(N399) );
  INVD1BWP30P140LVT U218 ( .I(i_data_bus[173]), .ZN(n179) );
  MAOI22D1BWP30P140LVT U219 ( .A1(n2), .A2(i_data_bus[205]), .B1(n180), .B2(
        n179), .ZN(n181) );
  IOA21D1BWP30P140LVT U220 ( .A1(n228), .A2(i_data_bus[237]), .B(n181), .ZN(
        n182) );
  AOI21D1BWP30P140LVT U221 ( .A1(n3), .A2(i_data_bus[13]), .B(n182), .ZN(n185)
         );
  AOI22D1BWP30P140LVT U222 ( .A1(n219), .A2(i_data_bus[77]), .B1(n1), .B2(
        i_data_bus[45]), .ZN(n184) );
  AOI22D1BWP30P140LVT U223 ( .A1(n220), .A2(i_data_bus[109]), .B1(n231), .B2(
        i_data_bus[141]), .ZN(n183) );
  ND3D1BWP30P140LVT U224 ( .A1(n185), .A2(n184), .A3(n183), .ZN(N382) );
  AOI22D1BWP30P140LVT U225 ( .A1(n2), .A2(i_data_bus[217]), .B1(n216), .B2(
        i_data_bus[185]), .ZN(n186) );
  IOA21D1BWP30P140LVT U226 ( .A1(n228), .A2(i_data_bus[249]), .B(n186), .ZN(
        n187) );
  AOI21D1BWP30P140LVT U227 ( .A1(n3), .A2(i_data_bus[25]), .B(n187), .ZN(n190)
         );
  AOI22D1BWP30P140LVT U228 ( .A1(n219), .A2(i_data_bus[89]), .B1(n1), .B2(
        i_data_bus[57]), .ZN(n189) );
  AOI22D1BWP30P140LVT U229 ( .A1(n220), .A2(i_data_bus[121]), .B1(n231), .B2(
        i_data_bus[153]), .ZN(n188) );
  ND3D1BWP30P140LVT U230 ( .A1(n190), .A2(n189), .A3(n188), .ZN(N394) );
  AOI22D1BWP30P140LVT U231 ( .A1(n2), .A2(i_data_bus[218]), .B1(n216), .B2(
        i_data_bus[186]), .ZN(n191) );
  IOA21D1BWP30P140LVT U232 ( .A1(n228), .A2(i_data_bus[250]), .B(n191), .ZN(
        n192) );
  AOI21D1BWP30P140LVT U233 ( .A1(n3), .A2(i_data_bus[26]), .B(n192), .ZN(n195)
         );
  AOI22D1BWP30P140LVT U234 ( .A1(n230), .A2(i_data_bus[90]), .B1(n1), .B2(
        i_data_bus[58]), .ZN(n194) );
  AOI22D1BWP30P140LVT U235 ( .A1(n232), .A2(i_data_bus[122]), .B1(n231), .B2(
        i_data_bus[154]), .ZN(n193) );
  ND3D1BWP30P140LVT U236 ( .A1(n195), .A2(n194), .A3(n193), .ZN(N395) );
  AOI22D1BWP30P140LVT U237 ( .A1(n2), .A2(i_data_bus[219]), .B1(n216), .B2(
        i_data_bus[187]), .ZN(n196) );
  IOA21D1BWP30P140LVT U238 ( .A1(n228), .A2(i_data_bus[251]), .B(n196), .ZN(
        n197) );
  AOI21D1BWP30P140LVT U239 ( .A1(n3), .A2(i_data_bus[27]), .B(n197), .ZN(n200)
         );
  AOI22D1BWP30P140LVT U240 ( .A1(n230), .A2(i_data_bus[91]), .B1(n1), .B2(
        i_data_bus[59]), .ZN(n199) );
  AOI22D1BWP30P140LVT U241 ( .A1(n232), .A2(i_data_bus[123]), .B1(n231), .B2(
        i_data_bus[155]), .ZN(n198) );
  ND3D1BWP30P140LVT U242 ( .A1(n200), .A2(n199), .A3(n198), .ZN(N396) );
  AOI22D1BWP30P140LVT U243 ( .A1(n2), .A2(i_data_bus[220]), .B1(n216), .B2(
        i_data_bus[188]), .ZN(n201) );
  IOA21D1BWP30P140LVT U244 ( .A1(n228), .A2(i_data_bus[252]), .B(n201), .ZN(
        n202) );
  AOI21D1BWP30P140LVT U245 ( .A1(n3), .A2(i_data_bus[28]), .B(n202), .ZN(n205)
         );
  AOI22D1BWP30P140LVT U246 ( .A1(n230), .A2(i_data_bus[92]), .B1(n1), .B2(
        i_data_bus[60]), .ZN(n204) );
  AOI22D1BWP30P140LVT U247 ( .A1(n232), .A2(i_data_bus[124]), .B1(n231), .B2(
        i_data_bus[156]), .ZN(n203) );
  ND3D1BWP30P140LVT U248 ( .A1(n205), .A2(n204), .A3(n203), .ZN(N397) );
  AOI22D1BWP30P140LVT U249 ( .A1(n2), .A2(i_data_bus[207]), .B1(n216), .B2(
        i_data_bus[175]), .ZN(n206) );
  IOA21D1BWP30P140LVT U250 ( .A1(n228), .A2(i_data_bus[239]), .B(n206), .ZN(
        n207) );
  AOI21D1BWP30P140LVT U251 ( .A1(n3), .A2(i_data_bus[15]), .B(n207), .ZN(n214)
         );
  INVD1BWP30P140LVT U252 ( .I(i_data_bus[79]), .ZN(n210) );
  INVD1BWP30P140LVT U253 ( .I(i_data_bus[47]), .ZN(n208) );
  OA22D1BWP30P140LVT U254 ( .A1(n211), .A2(n210), .B1(n209), .B2(n208), .Z(
        n213) );
  AOI22D1BWP30P140LVT U255 ( .A1(n220), .A2(i_data_bus[111]), .B1(n231), .B2(
        i_data_bus[143]), .ZN(n212) );
  ND3D1BWP30P140LVT U256 ( .A1(n214), .A2(n213), .A3(n212), .ZN(N384) );
  INVD1BWP30P140LVT U257 ( .I(i_data_bus[208]), .ZN(n215) );
  MAOI22D1BWP30P140LVT U258 ( .A1(n216), .A2(i_data_bus[176]), .B1(n225), .B2(
        n215), .ZN(n217) );
  IOA21D1BWP30P140LVT U259 ( .A1(n228), .A2(i_data_bus[240]), .B(n217), .ZN(
        n218) );
  AOI21D1BWP30P140LVT U260 ( .A1(n3), .A2(i_data_bus[16]), .B(n218), .ZN(n223)
         );
  AOI22D1BWP30P140LVT U261 ( .A1(n219), .A2(i_data_bus[80]), .B1(n1), .B2(
        i_data_bus[48]), .ZN(n222) );
  AOI22D1BWP30P140LVT U262 ( .A1(n220), .A2(i_data_bus[112]), .B1(n231), .B2(
        i_data_bus[144]), .ZN(n221) );
  ND3D1BWP30P140LVT U263 ( .A1(n223), .A2(n222), .A3(n221), .ZN(N385) );
  INVD1BWP30P140LVT U264 ( .I(i_data_bus[223]), .ZN(n224) );
  MAOI22D1BWP30P140LVT U265 ( .A1(n226), .A2(i_data_bus[191]), .B1(n225), .B2(
        n224), .ZN(n227) );
  IOA21D1BWP30P140LVT U266 ( .A1(n228), .A2(i_data_bus[255]), .B(n227), .ZN(
        n229) );
  AOI21D1BWP30P140LVT U267 ( .A1(n3), .A2(i_data_bus[31]), .B(n229), .ZN(n235)
         );
  AOI22D1BWP30P140LVT U268 ( .A1(n230), .A2(i_data_bus[95]), .B1(n1), .B2(
        i_data_bus[63]), .ZN(n234) );
  AOI22D1BWP30P140LVT U269 ( .A1(n232), .A2(i_data_bus[127]), .B1(n231), .B2(
        i_data_bus[159]), .ZN(n233) );
  ND3D1BWP30P140LVT U270 ( .A1(n235), .A2(n234), .A3(n233), .ZN(N400) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule


module crossbar_one_hot_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [63:0] i_cmd;
  input clk, rst, i_en;

  wire   [63:0] inner_valid_wire;
  wire   [2047:0] inner_data_wire;
  wire   [0:7] i_cmd_id_0__inner_cmd_wire;
  wire   [0:7] i_cmd_id_1__inner_cmd_wire;
  wire   [0:7] i_cmd_id_2__inner_cmd_wire;
  wire   [0:7] i_cmd_id_3__inner_cmd_wire;
  wire   [0:7] i_cmd_id_4__inner_cmd_wire;
  wire   [0:7] i_cmd_id_5__inner_cmd_wire;
  wire   [0:7] i_cmd_id_6__inner_cmd_wire;
  wire   [0:7] i_cmd_id_7__inner_cmd_wire;
  wire   [7:0] o_valid_wire;
  wire   [255:0] o_data_bus_wire;
  wire   [7:0] output_shift_def_0__o_valid_reg_shift;
  wire   [255:0] output_shift_def_0__o_data_bus_reg_shift;
  wire   [7:0] output_shift_def_1__o_valid_reg_shift;
  wire   [255:0] output_shift_def_1__o_data_bus_reg_shift;

  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 top_half_0__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[0]), .i_data_bus(
        i_data_bus[31:0]), .o_valid(inner_valid_wire[7:0]), .o_data_bus(
        inner_data_wire[255:0]), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 top_half_1__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[1]), .i_data_bus(
        i_data_bus[63:32]), .o_valid(inner_valid_wire[15:8]), .o_data_bus(
        inner_data_wire[511:256]), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 top_half_2__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[2]), .i_data_bus(
        i_data_bus[95:64]), .o_valid(inner_valid_wire[23:16]), .o_data_bus(
        inner_data_wire[767:512]), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 top_half_3__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[3]), .i_data_bus(
        i_data_bus[127:96]), .o_valid(inner_valid_wire[31:24]), .o_data_bus(
        inner_data_wire[1023:768]), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 top_half_4__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[4]), .i_data_bus(
        i_data_bus[159:128]), .o_valid(inner_valid_wire[39:32]), .o_data_bus(
        inner_data_wire[1279:1024]), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 top_half_5__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[5]), .i_data_bus(
        i_data_bus[191:160]), .o_valid(inner_valid_wire[47:40]), .o_data_bus(
        inner_data_wire[1535:1280]), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 top_half_6__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[6]), .i_data_bus(
        i_data_bus[223:192]), .o_valid(inner_valid_wire[55:48]), .o_data_bus(
        inner_data_wire[1791:1536]), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 top_half_7__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[7]), .i_data_bus(
        i_data_bus[255:224]), .o_valid(inner_valid_wire[63:56]), .o_data_bus(
        inner_data_wire[2047:1792]), .i_en(i_en) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 i_cmd_id_0__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(i_cmd_id_0__inner_cmd_wire[0]), 
        .o_cmd_1(i_cmd_id_0__inner_cmd_wire[1]), .o_cmd_2(
        i_cmd_id_0__inner_cmd_wire[2]), .o_cmd_3(i_cmd_id_0__inner_cmd_wire[3]), .o_cmd_4(i_cmd_id_0__inner_cmd_wire[4]), .o_cmd_5(
        i_cmd_id_0__inner_cmd_wire[5]), .o_cmd_6(i_cmd_id_0__inner_cmd_wire[6]), .o_cmd_7(i_cmd_id_0__inner_cmd_wire[7]), .i_en(i_en), .i_cmd(i_cmd[7:0]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 i_cmd_id_1__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(i_cmd_id_1__inner_cmd_wire[0]), 
        .o_cmd_1(i_cmd_id_1__inner_cmd_wire[1]), .o_cmd_2(
        i_cmd_id_1__inner_cmd_wire[2]), .o_cmd_3(i_cmd_id_1__inner_cmd_wire[3]), .o_cmd_4(i_cmd_id_1__inner_cmd_wire[4]), .o_cmd_5(
        i_cmd_id_1__inner_cmd_wire[5]), .o_cmd_6(i_cmd_id_1__inner_cmd_wire[6]), .o_cmd_7(i_cmd_id_1__inner_cmd_wire[7]), .i_en(i_en), .i_cmd(i_cmd[15:8]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 i_cmd_id_2__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(i_cmd_id_2__inner_cmd_wire[0]), 
        .o_cmd_1(i_cmd_id_2__inner_cmd_wire[1]), .o_cmd_2(
        i_cmd_id_2__inner_cmd_wire[2]), .o_cmd_3(i_cmd_id_2__inner_cmd_wire[3]), .o_cmd_4(i_cmd_id_2__inner_cmd_wire[4]), .o_cmd_5(
        i_cmd_id_2__inner_cmd_wire[5]), .o_cmd_6(i_cmd_id_2__inner_cmd_wire[6]), .o_cmd_7(i_cmd_id_2__inner_cmd_wire[7]), .i_en(i_en), .i_cmd(i_cmd[23:16])
         );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 i_cmd_id_3__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(i_cmd_id_3__inner_cmd_wire[0]), 
        .o_cmd_1(i_cmd_id_3__inner_cmd_wire[1]), .o_cmd_2(
        i_cmd_id_3__inner_cmd_wire[2]), .o_cmd_3(i_cmd_id_3__inner_cmd_wire[3]), .o_cmd_4(i_cmd_id_3__inner_cmd_wire[4]), .o_cmd_5(
        i_cmd_id_3__inner_cmd_wire[5]), .o_cmd_6(i_cmd_id_3__inner_cmd_wire[6]), .o_cmd_7(i_cmd_id_3__inner_cmd_wire[7]), .i_en(i_en), .i_cmd(i_cmd[31:24])
         );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 i_cmd_id_4__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(i_cmd_id_4__inner_cmd_wire[0]), 
        .o_cmd_1(i_cmd_id_4__inner_cmd_wire[1]), .o_cmd_2(
        i_cmd_id_4__inner_cmd_wire[2]), .o_cmd_3(i_cmd_id_4__inner_cmd_wire[3]), .o_cmd_4(i_cmd_id_4__inner_cmd_wire[4]), .o_cmd_5(
        i_cmd_id_4__inner_cmd_wire[5]), .o_cmd_6(i_cmd_id_4__inner_cmd_wire[6]), .o_cmd_7(i_cmd_id_4__inner_cmd_wire[7]), .i_en(i_en), .i_cmd(i_cmd[39:32])
         );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 i_cmd_id_5__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(i_cmd_id_5__inner_cmd_wire[0]), 
        .o_cmd_1(i_cmd_id_5__inner_cmd_wire[1]), .o_cmd_2(
        i_cmd_id_5__inner_cmd_wire[2]), .o_cmd_3(i_cmd_id_5__inner_cmd_wire[3]), .o_cmd_4(i_cmd_id_5__inner_cmd_wire[4]), .o_cmd_5(
        i_cmd_id_5__inner_cmd_wire[5]), .o_cmd_6(i_cmd_id_5__inner_cmd_wire[6]), .o_cmd_7(i_cmd_id_5__inner_cmd_wire[7]), .i_en(i_en), .i_cmd(i_cmd[47:40])
         );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 i_cmd_id_6__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(i_cmd_id_6__inner_cmd_wire[0]), 
        .o_cmd_1(i_cmd_id_6__inner_cmd_wire[1]), .o_cmd_2(
        i_cmd_id_6__inner_cmd_wire[2]), .o_cmd_3(i_cmd_id_6__inner_cmd_wire[3]), .o_cmd_4(i_cmd_id_6__inner_cmd_wire[4]), .o_cmd_5(
        i_cmd_id_6__inner_cmd_wire[5]), .o_cmd_6(i_cmd_id_6__inner_cmd_wire[6]), .o_cmd_7(i_cmd_id_6__inner_cmd_wire[7]), .i_en(i_en), .i_cmd(i_cmd[55:48])
         );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 i_cmd_id_7__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(i_cmd_id_7__inner_cmd_wire[0]), 
        .o_cmd_1(i_cmd_id_7__inner_cmd_wire[1]), .o_cmd_2(
        i_cmd_id_7__inner_cmd_wire[2]), .o_cmd_3(i_cmd_id_7__inner_cmd_wire[3]), .o_cmd_4(i_cmd_id_7__inner_cmd_wire[4]), .o_cmd_5(
        i_cmd_id_7__inner_cmd_wire[5]), .o_cmd_6(i_cmd_id_7__inner_cmd_wire[6]), .o_cmd_7(i_cmd_id_7__inner_cmd_wire[7]), .i_en(i_en), .i_cmd(i_cmd[63:56])
         );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_0 bottom_half_0__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid({inner_valid_wire[56], 
        inner_valid_wire[48], inner_valid_wire[40], inner_valid_wire[32], 
        inner_valid_wire[24], inner_valid_wire[16], inner_valid_wire[8], 
        inner_valid_wire[0]}), .i_data_bus({inner_data_wire[1823:1792], 
        inner_data_wire[1567:1536], inner_data_wire[1311:1280], 
        inner_data_wire[1055:1024], inner_data_wire[799:768], 
        inner_data_wire[543:512], inner_data_wire[287:256], 
        inner_data_wire[31:0]}), .o_valid(o_valid_wire[0]), .o_data_bus(
        o_data_bus_wire[31:0]), .i_en(i_en), .i_cmd({
        i_cmd_id_7__inner_cmd_wire[0], i_cmd_id_6__inner_cmd_wire[0], 
        i_cmd_id_5__inner_cmd_wire[0], i_cmd_id_4__inner_cmd_wire[0], 
        i_cmd_id_3__inner_cmd_wire[0], i_cmd_id_2__inner_cmd_wire[0], 
        i_cmd_id_1__inner_cmd_wire[0], i_cmd_id_0__inner_cmd_wire[0]}) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_7 bottom_half_1__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid({inner_valid_wire[57], 
        inner_valid_wire[49], inner_valid_wire[41], inner_valid_wire[33], 
        inner_valid_wire[25], inner_valid_wire[17], inner_valid_wire[9], 
        inner_valid_wire[1]}), .i_data_bus({inner_data_wire[1855:1824], 
        inner_data_wire[1599:1568], inner_data_wire[1343:1312], 
        inner_data_wire[1087:1056], inner_data_wire[831:800], 
        inner_data_wire[575:544], inner_data_wire[319:288], 
        inner_data_wire[63:32]}), .o_valid(o_valid_wire[1]), .o_data_bus(
        o_data_bus_wire[63:32]), .i_en(i_en), .i_cmd({
        i_cmd_id_7__inner_cmd_wire[1], i_cmd_id_6__inner_cmd_wire[1], 
        i_cmd_id_5__inner_cmd_wire[1], i_cmd_id_4__inner_cmd_wire[1], 
        i_cmd_id_3__inner_cmd_wire[1], i_cmd_id_2__inner_cmd_wire[1], 
        i_cmd_id_1__inner_cmd_wire[1], i_cmd_id_0__inner_cmd_wire[1]}) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_6 bottom_half_2__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid({inner_valid_wire[58], 
        inner_valid_wire[50], inner_valid_wire[42], inner_valid_wire[34], 
        inner_valid_wire[26], inner_valid_wire[18], inner_valid_wire[10], 
        inner_valid_wire[2]}), .i_data_bus({inner_data_wire[1887:1856], 
        inner_data_wire[1631:1600], inner_data_wire[1375:1344], 
        inner_data_wire[1119:1088], inner_data_wire[863:832], 
        inner_data_wire[607:576], inner_data_wire[351:320], 
        inner_data_wire[95:64]}), .o_valid(o_valid_wire[2]), .o_data_bus(
        o_data_bus_wire[95:64]), .i_en(i_en), .i_cmd({
        i_cmd_id_7__inner_cmd_wire[2], i_cmd_id_6__inner_cmd_wire[2], 
        i_cmd_id_5__inner_cmd_wire[2], i_cmd_id_4__inner_cmd_wire[2], 
        i_cmd_id_3__inner_cmd_wire[2], i_cmd_id_2__inner_cmd_wire[2], 
        i_cmd_id_1__inner_cmd_wire[2], i_cmd_id_0__inner_cmd_wire[2]}) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_5 bottom_half_3__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid({inner_valid_wire[59], 
        inner_valid_wire[51], inner_valid_wire[43], inner_valid_wire[35], 
        inner_valid_wire[27], inner_valid_wire[19], inner_valid_wire[11], 
        inner_valid_wire[3]}), .i_data_bus({inner_data_wire[1919:1888], 
        inner_data_wire[1663:1632], inner_data_wire[1407:1376], 
        inner_data_wire[1151:1120], inner_data_wire[895:864], 
        inner_data_wire[639:608], inner_data_wire[383:352], 
        inner_data_wire[127:96]}), .o_valid(o_valid_wire[3]), .o_data_bus(
        o_data_bus_wire[127:96]), .i_en(i_en), .i_cmd({
        i_cmd_id_7__inner_cmd_wire[3], i_cmd_id_6__inner_cmd_wire[3], 
        i_cmd_id_5__inner_cmd_wire[3], i_cmd_id_4__inner_cmd_wire[3], 
        i_cmd_id_3__inner_cmd_wire[3], i_cmd_id_2__inner_cmd_wire[3], 
        i_cmd_id_1__inner_cmd_wire[3], i_cmd_id_0__inner_cmd_wire[3]}) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_4 bottom_half_4__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid({inner_valid_wire[60], 
        inner_valid_wire[52], inner_valid_wire[44], inner_valid_wire[36], 
        inner_valid_wire[28], inner_valid_wire[20], inner_valid_wire[12], 
        inner_valid_wire[4]}), .i_data_bus({inner_data_wire[1951:1920], 
        inner_data_wire[1695:1664], inner_data_wire[1439:1408], 
        inner_data_wire[1183:1152], inner_data_wire[927:896], 
        inner_data_wire[671:640], inner_data_wire[415:384], 
        inner_data_wire[159:128]}), .o_valid(o_valid_wire[4]), .o_data_bus(
        o_data_bus_wire[159:128]), .i_en(i_en), .i_cmd({
        i_cmd_id_7__inner_cmd_wire[4], i_cmd_id_6__inner_cmd_wire[4], 
        i_cmd_id_5__inner_cmd_wire[4], i_cmd_id_4__inner_cmd_wire[4], 
        i_cmd_id_3__inner_cmd_wire[4], i_cmd_id_2__inner_cmd_wire[4], 
        i_cmd_id_1__inner_cmd_wire[4], i_cmd_id_0__inner_cmd_wire[4]}) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_3 bottom_half_5__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid({inner_valid_wire[61], 
        inner_valid_wire[53], inner_valid_wire[45], inner_valid_wire[37], 
        inner_valid_wire[29], inner_valid_wire[21], inner_valid_wire[13], 
        inner_valid_wire[5]}), .i_data_bus({inner_data_wire[1983:1952], 
        inner_data_wire[1727:1696], inner_data_wire[1471:1440], 
        inner_data_wire[1215:1184], inner_data_wire[959:928], 
        inner_data_wire[703:672], inner_data_wire[447:416], 
        inner_data_wire[191:160]}), .o_valid(o_valid_wire[5]), .o_data_bus(
        o_data_bus_wire[191:160]), .i_en(i_en), .i_cmd({
        i_cmd_id_7__inner_cmd_wire[5], i_cmd_id_6__inner_cmd_wire[5], 
        i_cmd_id_5__inner_cmd_wire[5], i_cmd_id_4__inner_cmd_wire[5], 
        i_cmd_id_3__inner_cmd_wire[5], i_cmd_id_2__inner_cmd_wire[5], 
        i_cmd_id_1__inner_cmd_wire[5], i_cmd_id_0__inner_cmd_wire[5]}) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_2 bottom_half_6__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid({inner_valid_wire[62], 
        inner_valid_wire[54], inner_valid_wire[46], inner_valid_wire[38], 
        inner_valid_wire[30], inner_valid_wire[22], inner_valid_wire[14], 
        inner_valid_wire[6]}), .i_data_bus({inner_data_wire[2015:1984], 
        inner_data_wire[1759:1728], inner_data_wire[1503:1472], 
        inner_data_wire[1247:1216], inner_data_wire[991:960], 
        inner_data_wire[735:704], inner_data_wire[479:448], 
        inner_data_wire[223:192]}), .o_valid(o_valid_wire[6]), .o_data_bus(
        o_data_bus_wire[223:192]), .i_en(i_en), .i_cmd({
        i_cmd_id_7__inner_cmd_wire[6], i_cmd_id_6__inner_cmd_wire[6], 
        i_cmd_id_5__inner_cmd_wire[6], i_cmd_id_4__inner_cmd_wire[6], 
        i_cmd_id_3__inner_cmd_wire[6], i_cmd_id_2__inner_cmd_wire[6], 
        i_cmd_id_1__inner_cmd_wire[6], i_cmd_id_0__inner_cmd_wire[6]}) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_1 bottom_half_7__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid({inner_valid_wire[63], 
        inner_valid_wire[55], inner_valid_wire[47], inner_valid_wire[39], 
        inner_valid_wire[31], inner_valid_wire[23], inner_valid_wire[15], 
        inner_valid_wire[7]}), .i_data_bus({inner_data_wire[2047:2016], 
        inner_data_wire[1791:1760], inner_data_wire[1535:1504], 
        inner_data_wire[1279:1248], inner_data_wire[1023:992], 
        inner_data_wire[767:736], inner_data_wire[511:480], 
        inner_data_wire[255:224]}), .o_valid(o_valid_wire[7]), .o_data_bus(
        o_data_bus_wire[255:224]), .i_en(i_en), .i_cmd({
        i_cmd_id_7__inner_cmd_wire[7], i_cmd_id_6__inner_cmd_wire[7], 
        i_cmd_id_5__inner_cmd_wire[7], i_cmd_id_4__inner_cmd_wire[7], 
        i_cmd_id_3__inner_cmd_wire[7], i_cmd_id_2__inner_cmd_wire[7], 
        i_cmd_id_1__inner_cmd_wire[7], i_cmd_id_0__inner_cmd_wire[7]}) );
  DFQD1BWP30P140LVT output_shift_def_0__o_valid_reg_shift_reg_7_ ( .D(
        o_valid_wire[7]), .CP(clk), .Q(
        output_shift_def_0__o_valid_reg_shift[7]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_valid_reg_shift_reg_6_ ( .D(
        o_valid_wire[6]), .CP(clk), .Q(
        output_shift_def_0__o_valid_reg_shift[6]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_valid_reg_shift_reg_5_ ( .D(
        o_valid_wire[5]), .CP(clk), .Q(
        output_shift_def_0__o_valid_reg_shift[5]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_valid_reg_shift_reg_4_ ( .D(
        o_valid_wire[4]), .CP(clk), .Q(
        output_shift_def_0__o_valid_reg_shift[4]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_valid_reg_shift_reg_3_ ( .D(
        o_valid_wire[3]), .CP(clk), .Q(
        output_shift_def_0__o_valid_reg_shift[3]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_valid_reg_shift_reg_2_ ( .D(
        o_valid_wire[2]), .CP(clk), .Q(
        output_shift_def_0__o_valid_reg_shift[2]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_valid_reg_shift_reg_1_ ( .D(
        o_valid_wire[1]), .CP(clk), .Q(
        output_shift_def_0__o_valid_reg_shift[1]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_valid_reg_shift_reg_0_ ( .D(
        o_valid_wire[0]), .CP(clk), .Q(
        output_shift_def_0__o_valid_reg_shift[0]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_255_ ( .D(
        o_data_bus_wire[255]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[255]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_254_ ( .D(
        o_data_bus_wire[254]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[254]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_253_ ( .D(
        o_data_bus_wire[253]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[253]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_252_ ( .D(
        o_data_bus_wire[252]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[252]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_251_ ( .D(
        o_data_bus_wire[251]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[251]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_250_ ( .D(
        o_data_bus_wire[250]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[250]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_249_ ( .D(
        o_data_bus_wire[249]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[249]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_248_ ( .D(
        o_data_bus_wire[248]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[248]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_247_ ( .D(
        o_data_bus_wire[247]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[247]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_246_ ( .D(
        o_data_bus_wire[246]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[246]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_245_ ( .D(
        o_data_bus_wire[245]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[245]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_244_ ( .D(
        o_data_bus_wire[244]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[244]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_243_ ( .D(
        o_data_bus_wire[243]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[243]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_242_ ( .D(
        o_data_bus_wire[242]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[242]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_241_ ( .D(
        o_data_bus_wire[241]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[241]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_240_ ( .D(
        o_data_bus_wire[240]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[240]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_239_ ( .D(
        o_data_bus_wire[239]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[239]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_238_ ( .D(
        o_data_bus_wire[238]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[238]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_237_ ( .D(
        o_data_bus_wire[237]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[237]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_236_ ( .D(
        o_data_bus_wire[236]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[236]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_235_ ( .D(
        o_data_bus_wire[235]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[235]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_234_ ( .D(
        o_data_bus_wire[234]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[234]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_233_ ( .D(
        o_data_bus_wire[233]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[233]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_232_ ( .D(
        o_data_bus_wire[232]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[232]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_231_ ( .D(
        o_data_bus_wire[231]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[231]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_230_ ( .D(
        o_data_bus_wire[230]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[230]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_229_ ( .D(
        o_data_bus_wire[229]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[229]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_228_ ( .D(
        o_data_bus_wire[228]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[228]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_227_ ( .D(
        o_data_bus_wire[227]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[227]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_226_ ( .D(
        o_data_bus_wire[226]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[226]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_225_ ( .D(
        o_data_bus_wire[225]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[225]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_224_ ( .D(
        o_data_bus_wire[224]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[224]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_223_ ( .D(
        o_data_bus_wire[223]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[223]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_222_ ( .D(
        o_data_bus_wire[222]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[222]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_221_ ( .D(
        o_data_bus_wire[221]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[221]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_220_ ( .D(
        o_data_bus_wire[220]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[220]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_219_ ( .D(
        o_data_bus_wire[219]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[219]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_218_ ( .D(
        o_data_bus_wire[218]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[218]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_217_ ( .D(
        o_data_bus_wire[217]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[217]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_216_ ( .D(
        o_data_bus_wire[216]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[216]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_215_ ( .D(
        o_data_bus_wire[215]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[215]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_214_ ( .D(
        o_data_bus_wire[214]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[214]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_213_ ( .D(
        o_data_bus_wire[213]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[213]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_212_ ( .D(
        o_data_bus_wire[212]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[212]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_211_ ( .D(
        o_data_bus_wire[211]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[211]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_210_ ( .D(
        o_data_bus_wire[210]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[210]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_209_ ( .D(
        o_data_bus_wire[209]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[209]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_208_ ( .D(
        o_data_bus_wire[208]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[208]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_207_ ( .D(
        o_data_bus_wire[207]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[207]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_206_ ( .D(
        o_data_bus_wire[206]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[206]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_205_ ( .D(
        o_data_bus_wire[205]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[205]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_204_ ( .D(
        o_data_bus_wire[204]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[204]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_203_ ( .D(
        o_data_bus_wire[203]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[203]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_202_ ( .D(
        o_data_bus_wire[202]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[202]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_201_ ( .D(
        o_data_bus_wire[201]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[201]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_200_ ( .D(
        o_data_bus_wire[200]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[200]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_199_ ( .D(
        o_data_bus_wire[199]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[199]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_198_ ( .D(
        o_data_bus_wire[198]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[198]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_197_ ( .D(
        o_data_bus_wire[197]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[197]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_196_ ( .D(
        o_data_bus_wire[196]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[196]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_195_ ( .D(
        o_data_bus_wire[195]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[195]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_194_ ( .D(
        o_data_bus_wire[194]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[194]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_193_ ( .D(
        o_data_bus_wire[193]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[193]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_192_ ( .D(
        o_data_bus_wire[192]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[192]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_191_ ( .D(
        o_data_bus_wire[191]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[191]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_190_ ( .D(
        o_data_bus_wire[190]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[190]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_189_ ( .D(
        o_data_bus_wire[189]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[189]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_188_ ( .D(
        o_data_bus_wire[188]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[188]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_187_ ( .D(
        o_data_bus_wire[187]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[187]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_186_ ( .D(
        o_data_bus_wire[186]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[186]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_185_ ( .D(
        o_data_bus_wire[185]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[185]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_184_ ( .D(
        o_data_bus_wire[184]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[184]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_183_ ( .D(
        o_data_bus_wire[183]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[183]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_182_ ( .D(
        o_data_bus_wire[182]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[182]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_181_ ( .D(
        o_data_bus_wire[181]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[181]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_180_ ( .D(
        o_data_bus_wire[180]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[180]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_179_ ( .D(
        o_data_bus_wire[179]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[179]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_178_ ( .D(
        o_data_bus_wire[178]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[178]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_177_ ( .D(
        o_data_bus_wire[177]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[177]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_176_ ( .D(
        o_data_bus_wire[176]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[176]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_175_ ( .D(
        o_data_bus_wire[175]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[175]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_174_ ( .D(
        o_data_bus_wire[174]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[174]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_173_ ( .D(
        o_data_bus_wire[173]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[173]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_172_ ( .D(
        o_data_bus_wire[172]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[172]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_171_ ( .D(
        o_data_bus_wire[171]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[171]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_170_ ( .D(
        o_data_bus_wire[170]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[170]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_169_ ( .D(
        o_data_bus_wire[169]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[169]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_168_ ( .D(
        o_data_bus_wire[168]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[168]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_167_ ( .D(
        o_data_bus_wire[167]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[167]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_166_ ( .D(
        o_data_bus_wire[166]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[166]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_165_ ( .D(
        o_data_bus_wire[165]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[165]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_164_ ( .D(
        o_data_bus_wire[164]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[164]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_163_ ( .D(
        o_data_bus_wire[163]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[163]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_162_ ( .D(
        o_data_bus_wire[162]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[162]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_161_ ( .D(
        o_data_bus_wire[161]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[161]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_160_ ( .D(
        o_data_bus_wire[160]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[160]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_159_ ( .D(
        o_data_bus_wire[159]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[159]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_158_ ( .D(
        o_data_bus_wire[158]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[158]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_157_ ( .D(
        o_data_bus_wire[157]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[157]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_156_ ( .D(
        o_data_bus_wire[156]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[156]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_155_ ( .D(
        o_data_bus_wire[155]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[155]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_154_ ( .D(
        o_data_bus_wire[154]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[154]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_153_ ( .D(
        o_data_bus_wire[153]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[153]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_152_ ( .D(
        o_data_bus_wire[152]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[152]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_151_ ( .D(
        o_data_bus_wire[151]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[151]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_150_ ( .D(
        o_data_bus_wire[150]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[150]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_149_ ( .D(
        o_data_bus_wire[149]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[149]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_148_ ( .D(
        o_data_bus_wire[148]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[148]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_147_ ( .D(
        o_data_bus_wire[147]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[147]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_146_ ( .D(
        o_data_bus_wire[146]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[146]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_145_ ( .D(
        o_data_bus_wire[145]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[145]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_144_ ( .D(
        o_data_bus_wire[144]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[144]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_143_ ( .D(
        o_data_bus_wire[143]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[143]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_142_ ( .D(
        o_data_bus_wire[142]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[142]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_141_ ( .D(
        o_data_bus_wire[141]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[141]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_140_ ( .D(
        o_data_bus_wire[140]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[140]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_139_ ( .D(
        o_data_bus_wire[139]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[139]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_138_ ( .D(
        o_data_bus_wire[138]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[138]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_137_ ( .D(
        o_data_bus_wire[137]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[137]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_136_ ( .D(
        o_data_bus_wire[136]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[136]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_135_ ( .D(
        o_data_bus_wire[135]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[135]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_134_ ( .D(
        o_data_bus_wire[134]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[134]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_133_ ( .D(
        o_data_bus_wire[133]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[133]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_132_ ( .D(
        o_data_bus_wire[132]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[132]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_131_ ( .D(
        o_data_bus_wire[131]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[131]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_130_ ( .D(
        o_data_bus_wire[130]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[130]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_129_ ( .D(
        o_data_bus_wire[129]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[129]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_128_ ( .D(
        o_data_bus_wire[128]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[128]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_127_ ( .D(
        o_data_bus_wire[127]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[127]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_126_ ( .D(
        o_data_bus_wire[126]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[126]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_125_ ( .D(
        o_data_bus_wire[125]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[125]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_124_ ( .D(
        o_data_bus_wire[124]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[124]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_123_ ( .D(
        o_data_bus_wire[123]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[123]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_122_ ( .D(
        o_data_bus_wire[122]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[122]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_121_ ( .D(
        o_data_bus_wire[121]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[121]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_120_ ( .D(
        o_data_bus_wire[120]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[120]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_119_ ( .D(
        o_data_bus_wire[119]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[119]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_118_ ( .D(
        o_data_bus_wire[118]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[118]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_117_ ( .D(
        o_data_bus_wire[117]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[117]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_116_ ( .D(
        o_data_bus_wire[116]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[116]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_115_ ( .D(
        o_data_bus_wire[115]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[115]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_114_ ( .D(
        o_data_bus_wire[114]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[114]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_113_ ( .D(
        o_data_bus_wire[113]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[113]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_112_ ( .D(
        o_data_bus_wire[112]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[112]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_111_ ( .D(
        o_data_bus_wire[111]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[111]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_110_ ( .D(
        o_data_bus_wire[110]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[110]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_109_ ( .D(
        o_data_bus_wire[109]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[109]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_108_ ( .D(
        o_data_bus_wire[108]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[108]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_107_ ( .D(
        o_data_bus_wire[107]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[107]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_106_ ( .D(
        o_data_bus_wire[106]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[106]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_105_ ( .D(
        o_data_bus_wire[105]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[105]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_104_ ( .D(
        o_data_bus_wire[104]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[104]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_103_ ( .D(
        o_data_bus_wire[103]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[103]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_102_ ( .D(
        o_data_bus_wire[102]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[102]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_101_ ( .D(
        o_data_bus_wire[101]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[101]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_100_ ( .D(
        o_data_bus_wire[100]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[100]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_99_ ( .D(
        o_data_bus_wire[99]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[99]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_98_ ( .D(
        o_data_bus_wire[98]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[98]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_97_ ( .D(
        o_data_bus_wire[97]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[97]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_96_ ( .D(
        o_data_bus_wire[96]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[96]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_95_ ( .D(
        o_data_bus_wire[95]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[95]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_94_ ( .D(
        o_data_bus_wire[94]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[94]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_93_ ( .D(
        o_data_bus_wire[93]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[93]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_92_ ( .D(
        o_data_bus_wire[92]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[92]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_91_ ( .D(
        o_data_bus_wire[91]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[91]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_90_ ( .D(
        o_data_bus_wire[90]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[90]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_89_ ( .D(
        o_data_bus_wire[89]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[89]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_88_ ( .D(
        o_data_bus_wire[88]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[88]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_87_ ( .D(
        o_data_bus_wire[87]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[87]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_86_ ( .D(
        o_data_bus_wire[86]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[86]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_85_ ( .D(
        o_data_bus_wire[85]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[85]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_84_ ( .D(
        o_data_bus_wire[84]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[84]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_83_ ( .D(
        o_data_bus_wire[83]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[83]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_82_ ( .D(
        o_data_bus_wire[82]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[82]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_81_ ( .D(
        o_data_bus_wire[81]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[81]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_80_ ( .D(
        o_data_bus_wire[80]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[80]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_79_ ( .D(
        o_data_bus_wire[79]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[79]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_78_ ( .D(
        o_data_bus_wire[78]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[78]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_77_ ( .D(
        o_data_bus_wire[77]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[77]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_76_ ( .D(
        o_data_bus_wire[76]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[76]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_75_ ( .D(
        o_data_bus_wire[75]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[75]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_74_ ( .D(
        o_data_bus_wire[74]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[74]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_73_ ( .D(
        o_data_bus_wire[73]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[73]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_72_ ( .D(
        o_data_bus_wire[72]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[72]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_71_ ( .D(
        o_data_bus_wire[71]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[71]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_70_ ( .D(
        o_data_bus_wire[70]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[70]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_69_ ( .D(
        o_data_bus_wire[69]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[69]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_68_ ( .D(
        o_data_bus_wire[68]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[68]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_67_ ( .D(
        o_data_bus_wire[67]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[67]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_66_ ( .D(
        o_data_bus_wire[66]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[66]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_65_ ( .D(
        o_data_bus_wire[65]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[65]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_64_ ( .D(
        o_data_bus_wire[64]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[64]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_63_ ( .D(
        o_data_bus_wire[63]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[63]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_62_ ( .D(
        o_data_bus_wire[62]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[62]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_61_ ( .D(
        o_data_bus_wire[61]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[61]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_60_ ( .D(
        o_data_bus_wire[60]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[60]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_59_ ( .D(
        o_data_bus_wire[59]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[59]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_58_ ( .D(
        o_data_bus_wire[58]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[58]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_57_ ( .D(
        o_data_bus_wire[57]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[57]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_56_ ( .D(
        o_data_bus_wire[56]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[56]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_55_ ( .D(
        o_data_bus_wire[55]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[55]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_54_ ( .D(
        o_data_bus_wire[54]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[54]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_53_ ( .D(
        o_data_bus_wire[53]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[53]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_52_ ( .D(
        o_data_bus_wire[52]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[52]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_51_ ( .D(
        o_data_bus_wire[51]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[51]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_50_ ( .D(
        o_data_bus_wire[50]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[50]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_49_ ( .D(
        o_data_bus_wire[49]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[49]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_48_ ( .D(
        o_data_bus_wire[48]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[48]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_47_ ( .D(
        o_data_bus_wire[47]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[47]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_46_ ( .D(
        o_data_bus_wire[46]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[46]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_45_ ( .D(
        o_data_bus_wire[45]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[45]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_44_ ( .D(
        o_data_bus_wire[44]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[44]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_43_ ( .D(
        o_data_bus_wire[43]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[43]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_42_ ( .D(
        o_data_bus_wire[42]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[42]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_41_ ( .D(
        o_data_bus_wire[41]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[41]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_40_ ( .D(
        o_data_bus_wire[40]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[40]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_39_ ( .D(
        o_data_bus_wire[39]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[39]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_38_ ( .D(
        o_data_bus_wire[38]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[38]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_37_ ( .D(
        o_data_bus_wire[37]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[37]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_36_ ( .D(
        o_data_bus_wire[36]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[36]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_35_ ( .D(
        o_data_bus_wire[35]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[35]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_34_ ( .D(
        o_data_bus_wire[34]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[34]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_33_ ( .D(
        o_data_bus_wire[33]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[33]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_32_ ( .D(
        o_data_bus_wire[32]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[32]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_31_ ( .D(
        o_data_bus_wire[31]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[31]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_30_ ( .D(
        o_data_bus_wire[30]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[30]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_29_ ( .D(
        o_data_bus_wire[29]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[29]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_28_ ( .D(
        o_data_bus_wire[28]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[28]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_27_ ( .D(
        o_data_bus_wire[27]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[27]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_26_ ( .D(
        o_data_bus_wire[26]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[26]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_25_ ( .D(
        o_data_bus_wire[25]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[25]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_24_ ( .D(
        o_data_bus_wire[24]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[24]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_23_ ( .D(
        o_data_bus_wire[23]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[23]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_22_ ( .D(
        o_data_bus_wire[22]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[22]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_21_ ( .D(
        o_data_bus_wire[21]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[21]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_20_ ( .D(
        o_data_bus_wire[20]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[20]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_19_ ( .D(
        o_data_bus_wire[19]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[19]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_18_ ( .D(
        o_data_bus_wire[18]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[18]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_17_ ( .D(
        o_data_bus_wire[17]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[17]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_16_ ( .D(
        o_data_bus_wire[16]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[16]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_15_ ( .D(
        o_data_bus_wire[15]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[15]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_14_ ( .D(
        o_data_bus_wire[14]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[14]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_13_ ( .D(
        o_data_bus_wire[13]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[13]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_12_ ( .D(
        o_data_bus_wire[12]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[12]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_11_ ( .D(
        o_data_bus_wire[11]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[11]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_10_ ( .D(
        o_data_bus_wire[10]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[10]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_9_ ( .D(
        o_data_bus_wire[9]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[9]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_8_ ( .D(
        o_data_bus_wire[8]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[8]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_7_ ( .D(
        o_data_bus_wire[7]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[7]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_6_ ( .D(
        o_data_bus_wire[6]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[6]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_5_ ( .D(
        o_data_bus_wire[5]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[5]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_4_ ( .D(
        o_data_bus_wire[4]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[4]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_3_ ( .D(
        o_data_bus_wire[3]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[3]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_2_ ( .D(
        o_data_bus_wire[2]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[2]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_1_ ( .D(
        o_data_bus_wire[1]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[1]) );
  DFQD1BWP30P140LVT output_shift_def_0__o_data_bus_reg_shift_reg_0_ ( .D(
        o_data_bus_wire[0]), .CP(clk), .Q(
        output_shift_def_0__o_data_bus_reg_shift[0]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_valid_reg_shift_reg_7_ ( .D(
        output_shift_def_0__o_valid_reg_shift[7]), .CP(clk), .Q(
        output_shift_def_1__o_valid_reg_shift[7]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_valid_reg_shift_reg_6_ ( .D(
        output_shift_def_0__o_valid_reg_shift[6]), .CP(clk), .Q(
        output_shift_def_1__o_valid_reg_shift[6]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_valid_reg_shift_reg_5_ ( .D(
        output_shift_def_0__o_valid_reg_shift[5]), .CP(clk), .Q(
        output_shift_def_1__o_valid_reg_shift[5]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_valid_reg_shift_reg_4_ ( .D(
        output_shift_def_0__o_valid_reg_shift[4]), .CP(clk), .Q(
        output_shift_def_1__o_valid_reg_shift[4]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_valid_reg_shift_reg_3_ ( .D(
        output_shift_def_0__o_valid_reg_shift[3]), .CP(clk), .Q(
        output_shift_def_1__o_valid_reg_shift[3]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_valid_reg_shift_reg_2_ ( .D(
        output_shift_def_0__o_valid_reg_shift[2]), .CP(clk), .Q(
        output_shift_def_1__o_valid_reg_shift[2]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_valid_reg_shift_reg_1_ ( .D(
        output_shift_def_0__o_valid_reg_shift[1]), .CP(clk), .Q(
        output_shift_def_1__o_valid_reg_shift[1]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_valid_reg_shift_reg_0_ ( .D(
        output_shift_def_0__o_valid_reg_shift[0]), .CP(clk), .Q(
        output_shift_def_1__o_valid_reg_shift[0]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_255_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[255]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[255]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_254_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[254]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[254]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_253_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[253]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[253]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_252_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[252]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[252]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_251_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[251]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[251]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_250_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[250]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[250]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_249_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[249]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[249]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_248_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[248]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[248]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_247_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[247]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[247]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_246_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[246]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[246]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_245_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[245]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[245]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_244_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[244]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[244]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_243_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[243]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[243]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_242_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[242]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[242]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_241_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[241]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[241]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_240_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[240]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[240]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_239_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[239]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[239]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_238_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[238]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[238]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_237_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[237]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[237]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_236_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[236]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[236]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_235_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[235]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[235]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_234_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[234]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[234]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_233_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[233]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[233]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_232_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[232]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[232]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_231_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[231]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[231]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_230_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[230]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[230]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_229_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[229]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[229]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_228_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[228]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[228]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_227_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[227]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[227]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_226_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[226]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[226]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_225_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[225]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[225]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_224_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[224]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[224]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_223_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[223]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[223]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_222_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[222]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[222]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_221_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[221]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[221]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_220_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[220]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[220]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_219_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[219]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[219]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_218_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[218]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[218]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_217_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[217]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[217]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_216_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[216]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[216]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_215_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[215]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[215]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_214_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[214]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[214]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_213_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[213]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[213]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_212_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[212]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[212]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_211_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[211]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[211]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_210_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[210]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[210]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_209_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[209]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[209]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_208_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[208]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[208]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_207_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[207]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[207]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_206_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[206]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[206]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_205_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[205]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[205]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_204_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[204]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[204]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_203_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[203]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[203]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_202_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[202]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[202]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_201_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[201]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[201]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_200_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[200]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[200]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_199_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[199]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[199]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_198_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[198]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[198]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_197_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[197]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[197]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_196_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[196]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[196]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_195_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[195]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[195]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_194_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[194]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[194]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_193_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[193]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[193]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_192_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[192]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[192]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_191_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[191]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[191]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_190_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[190]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[190]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_189_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[189]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[189]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_188_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[188]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[188]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_187_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[187]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[187]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_186_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[186]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[186]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_185_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[185]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[185]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_184_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[184]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[184]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_183_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[183]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[183]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_182_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[182]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[182]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_181_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[181]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[181]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_180_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[180]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[180]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_179_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[179]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[179]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_178_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[178]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[178]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_177_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[177]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[177]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_176_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[176]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[176]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_175_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[175]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[175]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_174_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[174]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[174]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_173_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[173]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[173]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_172_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[172]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[172]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_171_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[171]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[171]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_170_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[170]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[170]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_169_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[169]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[169]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_168_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[168]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[168]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_167_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[167]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[167]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_166_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[166]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[166]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_165_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[165]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[165]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_164_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[164]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[164]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_163_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[163]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[163]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_162_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[162]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[162]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_161_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[161]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[161]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_160_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[160]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[160]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_159_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[159]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[159]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_158_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[158]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[158]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_157_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[157]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[157]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_156_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[156]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[156]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_155_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[155]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[155]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_154_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[154]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[154]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_153_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[153]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[153]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_152_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[152]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[152]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_151_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[151]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[151]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_150_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[150]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[150]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_149_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[149]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[149]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_148_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[148]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[148]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_147_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[147]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[147]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_146_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[146]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[146]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_145_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[145]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[145]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_144_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[144]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[144]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_143_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[143]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[143]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_142_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[142]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[142]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_141_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[141]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[141]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_140_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[140]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[140]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_139_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[139]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[139]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_138_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[138]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[138]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_137_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[137]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[137]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_136_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[136]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[136]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_135_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[135]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[135]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_134_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[134]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[134]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_133_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[133]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[133]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_132_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[132]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[132]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_131_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[131]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[131]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_130_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[130]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[130]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_129_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[129]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[129]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_128_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[128]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[128]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_127_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[127]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[127]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_126_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[126]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[126]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_125_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[125]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[125]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_124_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[124]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[124]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_123_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[123]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[123]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_122_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[122]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[122]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_121_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[121]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[121]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_120_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[120]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[120]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_119_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[119]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[119]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_118_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[118]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[118]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_117_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[117]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[117]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_116_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[116]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[116]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_115_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[115]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[115]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_114_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[114]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[114]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_113_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[113]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[113]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_112_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[112]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[112]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_111_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[111]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[111]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_110_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[110]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[110]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_109_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[109]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[109]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_108_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[108]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[108]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_107_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[107]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[107]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_106_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[106]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[106]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_105_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[105]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[105]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_104_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[104]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[104]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_103_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[103]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[103]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_102_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[102]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[102]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_101_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[101]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[101]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_100_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[100]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[100]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_99_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[99]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[99]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_98_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[98]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[98]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_97_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[97]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[97]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_96_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[96]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[96]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_95_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[95]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[95]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_94_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[94]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[94]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_93_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[93]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[93]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_92_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[92]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[92]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_91_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[91]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[91]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_90_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[90]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[90]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_89_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[89]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[89]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_88_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[88]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[88]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_87_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[87]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[87]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_86_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[86]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[86]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_85_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[85]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[85]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_84_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[84]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[84]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_83_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[83]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[83]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_82_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[82]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[82]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_81_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[81]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[81]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_80_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[80]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[80]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_79_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[79]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[79]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_78_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[78]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[78]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_77_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[77]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[77]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_76_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[76]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[76]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_75_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[75]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[75]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_74_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[74]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[74]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_73_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[73]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[73]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_72_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[72]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[72]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_71_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[71]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[71]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_70_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[70]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[70]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_69_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[69]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[69]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_68_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[68]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[68]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_67_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[67]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[67]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_66_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[66]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[66]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_65_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[65]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[65]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_64_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[64]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[64]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_63_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[63]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[63]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_62_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[62]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[62]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_61_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[61]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[61]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_60_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[60]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[60]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_59_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[59]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[59]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_58_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[58]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[58]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_57_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[57]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[57]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_56_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[56]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[56]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_55_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[55]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[55]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_54_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[54]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[54]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_53_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[53]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[53]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_52_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[52]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[52]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_51_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[51]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[51]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_50_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[50]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[50]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_49_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[49]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[49]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_48_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[48]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[48]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_47_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[47]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[47]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_46_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[46]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[46]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_45_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[45]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[45]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_44_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[44]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[44]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_43_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[43]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[43]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_42_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[42]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[42]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_41_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[41]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[41]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_40_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[40]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[40]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_39_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[39]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[39]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_38_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[38]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[38]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_37_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[37]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[37]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_36_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[36]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[36]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_35_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[35]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[35]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_34_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[34]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[34]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_33_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[33]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[33]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_32_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[32]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[32]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_31_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[31]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[31]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_30_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[30]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[30]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_29_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[29]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[29]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_28_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[28]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[28]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_27_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[27]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[27]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_26_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[26]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[26]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_25_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[25]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[25]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_24_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[24]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[24]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_23_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[23]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[23]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_22_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[22]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[22]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_21_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[21]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[21]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_20_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[20]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[20]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_19_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[19]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[19]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_18_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[18]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[18]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_17_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[17]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[17]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_16_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[16]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[16]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_15_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[15]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[15]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_14_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[14]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[14]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_13_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[13]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[13]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_12_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[12]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[12]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_11_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[11]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[11]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_10_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[10]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[10]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_9_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[9]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[9]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_8_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[8]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[8]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_7_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[7]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[7]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_6_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[6]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[6]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_5_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[5]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[5]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_4_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[4]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[4]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_3_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[3]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[3]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_2_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[2]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[2]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_1_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[1]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[1]) );
  DFQD1BWP30P140LVT output_shift_def_1__o_data_bus_reg_shift_reg_0_ ( .D(
        output_shift_def_0__o_data_bus_reg_shift[0]), .CP(clk), .Q(
        output_shift_def_1__o_data_bus_reg_shift[0]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_7_ ( .D(
        output_shift_def_1__o_valid_reg_shift[7]), .CP(clk), .Q(o_valid[7]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_6_ ( .D(
        output_shift_def_1__o_valid_reg_shift[6]), .CP(clk), .Q(o_valid[6]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_5_ ( .D(
        output_shift_def_1__o_valid_reg_shift[5]), .CP(clk), .Q(o_valid[5]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_4_ ( .D(
        output_shift_def_1__o_valid_reg_shift[4]), .CP(clk), .Q(o_valid[4]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_3_ ( .D(
        output_shift_def_1__o_valid_reg_shift[3]), .CP(clk), .Q(o_valid[3]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_2_ ( .D(
        output_shift_def_1__o_valid_reg_shift[2]), .CP(clk), .Q(o_valid[2]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_1_ ( .D(
        output_shift_def_1__o_valid_reg_shift[1]), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_0_ ( .D(
        output_shift_def_1__o_valid_reg_shift[0]), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[255]), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[254]), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[253]), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[252]), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[251]), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[250]), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[249]), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[248]), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[247]), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[246]), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[245]), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[244]), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[243]), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[242]), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[241]), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[240]), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[239]), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[238]), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[237]), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[236]), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[235]), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[234]), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[233]), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[232]), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[231]), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[230]), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[229]), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[228]), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[227]), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[226]), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[225]), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[224]), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[223]), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[222]), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[221]), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[220]), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[219]), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[218]), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[217]), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[216]), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[215]), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[214]), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[213]), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[212]), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[211]), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[210]), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[209]), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[208]), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[207]), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[206]), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[205]), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[204]), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[203]), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[202]), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[201]), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[200]), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[199]), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[198]), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[197]), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[196]), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[195]), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[194]), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[193]), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[192]), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[191]), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[190]), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[189]), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[188]), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[187]), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[186]), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[185]), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[184]), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[183]), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[182]), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[181]), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[180]), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[179]), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[178]), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[177]), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[176]), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[175]), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[174]), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[173]), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[172]), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[171]), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[170]), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[169]), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[168]), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[167]), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[166]), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[165]), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[164]), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[163]), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[162]), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[161]), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[160]), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[159]), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[158]), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[157]), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[156]), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[155]), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[154]), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[153]), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[152]), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[151]), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[150]), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[149]), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[148]), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[147]), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[146]), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[145]), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[144]), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[143]), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[142]), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[141]), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[140]), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[139]), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[138]), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[137]), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[136]), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[135]), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[134]), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[133]), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[132]), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[131]), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[130]), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[129]), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[128]), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[127]), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[126]), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[125]), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[124]), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[123]), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[122]), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[121]), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[120]), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[119]), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[118]), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[117]), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[116]), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[115]), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[114]), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[113]), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[112]), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[111]), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[110]), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[109]), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[108]), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[107]), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[106]), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[105]), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[104]), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[103]), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[102]), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[101]), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[100]), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[99]), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[98]), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[97]), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[96]), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[95]), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[94]), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[93]), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[92]), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[91]), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[90]), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[89]), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[88]), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[87]), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[86]), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[85]), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[84]), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[83]), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[82]), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[81]), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[80]), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[79]), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[78]), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[77]), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[76]), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[75]), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[74]), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[73]), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[72]), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[71]), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[70]), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[69]), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[68]), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[67]), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[66]), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[65]), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[64]), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[63]), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[62]), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[61]), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[60]), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[59]), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[58]), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[57]), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[56]), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[55]), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[54]), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[53]), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[52]), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[51]), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[50]), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[49]), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[48]), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[47]), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[46]), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[45]), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[44]), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[43]), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[42]), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[41]), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[40]), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[39]), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[38]), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[37]), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[36]), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[35]), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[34]), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[33]), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[32]), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[31]), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[30]), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[29]), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[28]), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[27]), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[26]), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[25]), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[24]), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[23]), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[22]), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[21]), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[20]), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[19]), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[18]), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[17]), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[16]), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[15]), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[14]), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[13]), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[12]), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[11]), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[10]), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[9]), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[8]), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[7]), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[6]), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[5]), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[4]), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[3]), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[2]), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[1]), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(
        output_shift_def_1__o_data_bus_reg_shift[0]), .CP(clk), .Q(
        o_data_bus[0]) );
endmodule

