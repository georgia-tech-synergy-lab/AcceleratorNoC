`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 03/31/2021 
// System Name: accelerator
// Module Name: table parse engine 
// Project Name: ARION DRBE
// Description: Decode elements of delay table
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module table_parse_engine(CLK, reset, boot_up, table_parse, input_valid, glob_scen_noc_input_valid, delay_matrix_element, obj_id_element, local_controller_id, calc_glob_controller_delay, calc_glob_dest_addr, tapping_loc_packet, scenario_update);

    // parameter
    	parameter N_sample = 256;
	parameter datawidth = 16;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for small tapeout
	parameter N_obj = 8; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 4; // 16 local controllers in subscaled system
	parameter sample_address_width = 8; /// assuming 256 words: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	parameter delay_length = 12; // log(id_width*N_sample)
	parameter obj_id_width = 3; // log(N_obj)
	parameter tapping_loc_packet_width = sample_address_width + obj_id_width; // log(N_obj)
	

//=== IO Ports ===//


    // input
    	input CLK; // system clock, generated by VCO
	input reset;
	input [delay_length - 1:0] delay_matrix_element;
	input [obj_id_width - 1:0] obj_id_element;
	input boot_up;
	input table_parse;
	input input_valid;
	input glob_scen_noc_input_valid;
	input scenario_update;
    // output

	output reg [address_vector_width - 1:0] calc_glob_dest_addr;
	output reg [sample_address_width - 1:0] calc_glob_controller_delay;
	//output reg [sample_address_width - 1:0] calc_glob_prefetch_stop;
	output reg [tapping_loc_packet_width - 1:0] tapping_loc_packet;
	output reg [id_width - 1:0] local_controller_id;




//////////// internal status regs/signals //////////////////////////////////
	reg done;
	reg [obj_id_width - 1:0] group_header;
	reg [obj_id_width - 1:0] table_ptr;
	reg [obj_id_width - 1:0] pointer;
	reg [obj_id_width - 1:0] ptr_next;
	wire [obj_id_width - 1:0] index;
	reg [delay_length - 1:0] delay_matrix_N_1[N_obj - 1:0];
	reg [delay_length - 1:0] delay_matrix_N_1_next[N_obj - 1:0];
	reg [obj_id_width - 1:0] obj_id[N_obj - 1:0];
	reg [obj_id_width - 1:0] obj_id_next[N_obj - 1:0];
	reg [9:0] scenario_counter;

	integer i;
	integer j;
	integer k;



///////////////////////////////////////////////////////////////////////////////    

////////// logic part ///////////////////////////////////////////////////////  

	assign index = obj_id[table_ptr];


////////////sequential logic
//
//


	always @(posedge CLK) begin
		if (reset) begin
			for (i = 0; i < N_obj; i = i + 1) begin
				delay_matrix_N_1[i] <= 12'hfff;
				obj_id[i] <= 0;
				pointer <= 0;
			end
		end
		else if (scenario_update) begin
			for (i=0;i<N_obj;i=i+1) begin
				delay_matrix_N_1[i] <= delay_matrix_N_1_next[i];
				obj_id[i] <= obj_id_next[i];
			end
			pointer <= 0;

		end

		else if (boot_up) begin
			if (input_valid) begin
				for (k = 0; k< N_obj ; k=k+1) begin
					if (k[2:0]==pointer) begin
						delay_matrix_N_1[k] <= delay_matrix_element;
						obj_id[k] <= obj_id_element;
					end
					else begin
						delay_matrix_N_1[k] <= delay_matrix_N_1[k];
						obj_id[k] <= obj_id[k];
					end
				end
				pointer <= pointer + 1;
			end
			else begin
				for (i=0;i<N_obj;i=i+1) begin
					delay_matrix_N_1[i] <= delay_matrix_N_1[i];
					obj_id[i] <= obj_id[i];
				end
				pointer <= pointer;
			end
			
		end
		else begin
			for (i=0;i<N_obj;i=i+1) begin
				delay_matrix_N_1[i] <= delay_matrix_N_1[i];
				obj_id[i] <= obj_id[i];
			end
			pointer <= pointer;
		end

	end

	always @(posedge CLK) begin
//		if (reset) begin
			for (i = 0; i < N_obj; i = i + 1) begin
				delay_matrix_N_1_next[i] <= 12'hfff;
				obj_id_next[i] <= 0;
				ptr_next <= 0;
			end
//		end

//		else if (glob_scen_noc_input_valid) begin
		//	if (input_valid) begin
//				delay_matrix_N_1_next[ptr_next] <= delay_matrix_element;
//				obj_id_next[ptr_next] <= obj_id_element;
//				ptr_next <= ptr_next + 1;
		//	end
		//	else begin
		//		delay_matrix_N_1[pointer] <= delay_matrix_N_1[pointer];
		//		obj_id[pointer] <= obj_id[pointer];
		//		pointer <= pointer;
		//	end
			
//		end
//		else begin
//			delay_matrix_N_1_next[ptr_next] <= delay_matrix_N_1_next[ptr_next];
//			obj_id_next[ptr_next] <= obj_id[ptr_next];
//			ptr_next <= ptr_next;
//		end

	end





        always @(posedge CLK) begin
		if (reset | scenario_update) begin
			table_ptr <= 0;
			done <= 0;
		end
		else if (table_parse) begin
			if (done) begin
				table_ptr <= 0;
				done <= done;
			end
			else begin
				if (table_ptr == N_obj - 1 || delay_matrix_N_1[table_ptr] == 12'hfff ) begin
					table_ptr <= 0;
					done <= 1;
				end
				else  begin
					table_ptr <= table_ptr + 1;
					done <= done;
				end
			end

		end
		else begin
			table_ptr <= 0;
			done <= 0;
		end



	end


	always @(posedge CLK) begin	
		if (reset) begin
			group_header <= 0;
			tapping_loc_packet <= 11'bz;
			calc_glob_dest_addr <= 8'b0;
			calc_glob_controller_delay <= 8'bz;
			local_controller_id <= 4'bz;
		end
		else if (table_parse)begin
			if (done) begin    ////indicates table parsing done
					group_header <= group_header;
					calc_glob_dest_addr <= calc_glob_dest_addr;
					tapping_loc_packet <= 11'bz;
					calc_glob_controller_delay <= 8'bz;
					local_controller_id <= 4'bz;
			end
			else begin
				if (table_ptr == 0 ) begin
						group_header <= table_ptr;
						tapping_loc_packet <= {8'b0,index};   //no need to send this really
						calc_glob_controller_delay <= delay_matrix_N_1[table_ptr][7:0];
						local_controller_id <= delay_matrix_N_1[table_ptr][11:8];
						for (i=0;i<N_obj;i=i+1) begin
							if (i == index) begin
								calc_glob_dest_addr[i] <= 1;
							end
							else begin
								calc_glob_dest_addr[i] <= 0;
							end
						end

				end

				else if (delay_matrix_N_1[table_ptr] - delay_matrix_N_1[group_header] >= N_sample) begin
						group_header <= table_ptr;
						tapping_loc_packet <= {8'b0,index};   //no need to send this really
						calc_glob_controller_delay <= delay_matrix_N_1[table_ptr][7:0];
						local_controller_id <= delay_matrix_N_1[table_ptr][11:8];
						for (i=0;i<N_obj;i=i+1) begin
							if (i == index) begin
								calc_glob_dest_addr[i] <= 1;
							end
							else begin
								calc_glob_dest_addr[i] <= 0;
							end
						end

				end
				else if (delay_matrix_N_1[table_ptr] - delay_matrix_N_1[group_header] < N_sample) begin
						for (i=0;i<N_obj;i=i+1) begin
							if (i == index) begin
								calc_glob_dest_addr[i] <= 1;
							end
							else begin
								calc_glob_dest_addr[i] <= calc_glob_dest_addr[i] ;
							end
						end

						tapping_loc_packet <=  {(delay_matrix_N_1[table_ptr] - delay_matrix_N_1[group_header]),index};
						group_header <= group_header;
						calc_glob_controller_delay <= 8'bz;
						local_controller_id <= 4'bz;
				end
				else begin
						group_header <= group_header;
						calc_glob_dest_addr <= calc_glob_dest_addr;
						tapping_loc_packet <= 11'bz;
						calc_glob_controller_delay <= 8'bz;
						local_controller_id <= 4'bz;


				end
			end
		end
		else begin
			group_header <= 0;
			tapping_loc_packet <= 11'bz;
			calc_glob_dest_addr <= 8'b0;
			calc_glob_controller_delay <= 8'bz;
			local_controller_id <= 4'bz;
		end


	end
	 
	 


   
endmodule
    

