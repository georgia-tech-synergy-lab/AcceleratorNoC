`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module small_trial(clk, reset, a, b, out );
    // parameter
       
    // input
    	input clk; // system clock, generated by VCO
	input reset;
	input a;
	input b;



    // output
	output reg out;	
	

    // internal status regs/signals



	//sequential logic
    always @ (posedge clk) begin
        if (reset) begin
		out <= 0;	
        end
	else begin
		out <= a + b;

	end  
     end
	 
	 


   
endmodule
    
