`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module local_controller_v1(clk, reset, init, controller_id, write_flag, data_from_sram, input_boundary_flag, prev_dest_address, from_glob_dest_addr, packet_out, boundary_next);
    // parameter
    parameter N_row = 1024;
	parameter datawidth = 32;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for subscaled system
	parameter id_width = 11; // 1221 local controllers in subscaled system
	parameter row_address_width = 10; /// assuming 1024 rows and 64 columns: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	
	
	
        
    // input
    input clk; // system clock, generated by VCO
	input reset;
	input init;
	input [2*datawidth - 1:0] data_from_sram;
	input [id_width - 1:0] controller_id;
	input input_boundary_flag;
	input write_flag;
	input [address_vector_width - 1:0] prev_dest_address;
	input [address_vector_width - 1:0] from_glob_dest_addr;

    // output
    output [packet_width-1:0] packet_out; 
    output reg boundary_next; 
	
	

    // internal status regs/signals
    reg [row_address_width-1:0] row_address;
	reg id; 
	reg [packet_width-1:0] packet_out_internal;
	reg [address_vector_width - 1:0] dest_address;
	reg coeff_num;
    

    // logic part  
    assign packet_out = packet_out_internal;

	//sequential logic
    always @ (posedge clk) begin
        if (reset) begin
			id <= 0;
			row_address <= 0;
			packet_out_internal <= 0;
			dest_address <= 0;
			
        end
        else if (init) begin
			id <= controller_id;
			row_address <= row_address;
			packet_out_internal <= 0;
			dest_address <= 0;
			
        end
		else begin
			if (coeff_num == 1 && write_flag == 0) begin
				packet_out_internal <= {data_from_sram, dest_address};
				
			end
			else if (coeff_num == 1 && write_flag == 1) begin
				packet_out_internal <= {64'b0, dest_address};				
			end
			else if (coeff_num == 0) begin
				packet_out_internal <= 264'bz;
			end
			id <= id;
			row_address <= row_address + 1;
			dest_address <= dest_address;
		end  
     end
	 
	 always @ (posedge clk) begin
		if (row_address == N_row - 1) begin
			boundary_next <= 1;
		end
		else begin
			boundary_next <= 0;
		end
	 end
	 
	 
	 always @ (negedge clk) begin
		boundary_next <= 0;
		if (input_boundary_flag == 1) begin
			coeff_num <= 1;
			row_address <= 0;
			dest_address <= prev_dest_address;
		end
		else if (input_boundary_flag == 0) begin
			if (boundary_next == 1) begin
				coeff_num <= 0;
			end
			else begin
				coeff_num <= 1;
			end
			row_address <= row_address;
			dest_address <= dest_address;
			
		end
	 end
	 
	 


   
endmodule
    
