
module crossbar_one_hot_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(n561) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(n562) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(n563) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(n564) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(n565) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(n566) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(n567) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(n568) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(n569) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(n570) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(n571) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(n572) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(n573) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(n574) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(n575) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(n576) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(n577) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(n578) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(n579) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(n580) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(n581) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(n582) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(n583) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(n584) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(n585) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(n586) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(n587) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(n588) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(n589) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(n590) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(n591) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(n592) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(n593) );
  INVD4BWP30P140LVT U197 ( .I(n406), .ZN(n165) );
  INVD3BWP30P140LVT U198 ( .I(n231), .ZN(n408) );
  INVD1BWP30P140LVT U199 ( .I(n234), .ZN(n166) );
  CKND2D2BWP30P140LVT U200 ( .A1(n221), .A2(n220), .ZN(n222) );
  NR2OPTPAD1BWP30P140LVT U201 ( .A1(n218), .A2(n217), .ZN(n221) );
  NR3D1P5BWP30P140LVT U202 ( .A1(rst), .A2(n244), .A3(n243), .ZN(n245) );
  ND2OPTIBD1BWP30P140LVT U203 ( .A1(i_cmd[6]), .A2(n257), .ZN(n241) );
  NR3D2BWP30P140LVT U204 ( .A1(rst), .A2(i_cmd[0]), .A3(i_cmd[1]), .ZN(n234)
         );
  NR2D1BWP30P140LVT U205 ( .A1(n249), .A2(i_cmd[7]), .ZN(n250) );
  INVD1BWP30P140LVT U206 ( .I(rst), .ZN(n213) );
  INVD2BWP30P140LVT U207 ( .I(i_cmd[4]), .ZN(n232) );
  INVD1BWP30P140LVT U208 ( .I(i_cmd[1]), .ZN(n228) );
  NR2OPTPAD4BWP30P140LVT U209 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n257) );
  NR2OPTPAD1BWP30P140LVT U210 ( .A1(i_cmd[1]), .A2(i_cmd[4]), .ZN(n238) );
  NR2D2BWP30P140LVT U211 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .ZN(n215) );
  NR2OPTPAD1BWP30P140LVT U212 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .ZN(n216) );
  INVD6BWP30P140LVT U213 ( .I(i_en), .ZN(n169) );
  NR2OPTPAD4BWP30P140LVT U214 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n224) );
  INVD2BWP30P140LVT U215 ( .I(n225), .ZN(n226) );
  ND3D2BWP30P140LVT U216 ( .A1(n259), .A2(i_valid[3]), .A3(i_cmd[3]), .ZN(n260) );
  CKAN2D4BWP30P140LVT U217 ( .A1(n258), .A2(n170), .Z(n162) );
  ND2OPTPAD4BWP30P140LVT U218 ( .A1(n226), .A2(n168), .ZN(n261) );
  INVD12BWP30P140LVT U219 ( .I(n288), .ZN(n163) );
  INVD6BWP30P140LVT U220 ( .I(n408), .ZN(n164) );
  INVD8BWP30P140LVT U221 ( .I(n173), .ZN(n524) );
  INVD4BWP30P140LVT U222 ( .I(n222), .ZN(n288) );
  INVD6BWP30P140LVT U223 ( .I(n167), .ZN(n172) );
  INVD2BWP30P140LVT U224 ( .I(n251), .ZN(n253) );
  NR2D3BWP30P140LVT U225 ( .A1(n241), .A2(n240), .ZN(n246) );
  AN2D4BWP30P140LVT U226 ( .A1(n211), .A2(n212), .Z(n171) );
  NR3D3BWP30P140LVT U227 ( .A1(n166), .A2(n233), .A3(n236), .ZN(n523) );
  NR2OPTPAD1BWP30P140LVT U228 ( .A1(i_cmd[3]), .A2(i_cmd[5]), .ZN(n214) );
  ND2D1BWP30P140LVT U229 ( .A1(n215), .A2(n214), .ZN(n208) );
  ND2D1BWP30P140LVT U230 ( .A1(n242), .A2(i_cmd[4]), .ZN(n210) );
  INR2D4BWP30P140LVT U231 ( .A1(n234), .B1(n233), .ZN(n252) );
  ND3OPTPAD6BWP30P140LVT U232 ( .A1(n257), .A2(i_en), .A3(n232), .ZN(n233) );
  ND2D1BWP30P140LVT U233 ( .A1(n248), .A2(n247), .ZN(n255) );
  ND2D1BWP30P140LVT U234 ( .A1(n172), .A2(i_data_bus[198]), .ZN(n247) );
  ND2D1BWP30P140LVT U235 ( .A1(n164), .A2(i_data_bus[74]), .ZN(n276) );
  ND2D1BWP30P140LVT U236 ( .A1(n165), .A2(i_data_bus[170]), .ZN(n277) );
  ND2D1BWP30P140LVT U237 ( .A1(n164), .A2(i_data_bus[76]), .ZN(n491) );
  ND2D1BWP30P140LVT U238 ( .A1(n165), .A2(i_data_bus[172]), .ZN(n492) );
  ND2OPTIBD2BWP30P140LVT U239 ( .A1(n242), .A2(i_en), .ZN(n244) );
  INVD1BWP30P140LVT U240 ( .I(i_valid[6]), .ZN(n243) );
  ND2OPTIBD2BWP30P140LVT U241 ( .A1(n239), .A2(n238), .ZN(n240) );
  NR2D1BWP30P140LVT U242 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .ZN(n239) );
  ND2OPTIBD1BWP30P140LVT U243 ( .A1(n216), .A2(n215), .ZN(n217) );
  ND2D1BWP30P140LVT U244 ( .A1(n164), .A2(i_data_bus[64]), .ZN(n390) );
  ND2D1BWP30P140LVT U245 ( .A1(n165), .A2(i_data_bus[160]), .ZN(n391) );
  ND2D1BWP30P140LVT U246 ( .A1(n164), .A2(i_data_bus[65]), .ZN(n382) );
  ND2D1BWP30P140LVT U247 ( .A1(n165), .A2(i_data_bus[161]), .ZN(n383) );
  ND2D1BWP30P140LVT U248 ( .A1(n164), .A2(i_data_bus[66]), .ZN(n374) );
  ND2D1BWP30P140LVT U249 ( .A1(n165), .A2(i_data_bus[162]), .ZN(n375) );
  ND2D1BWP30P140LVT U250 ( .A1(n164), .A2(i_data_bus[67]), .ZN(n366) );
  ND2D1BWP30P140LVT U251 ( .A1(n165), .A2(i_data_bus[163]), .ZN(n367) );
  ND2D1BWP30P140LVT U252 ( .A1(n164), .A2(i_data_bus[68]), .ZN(n358) );
  ND2D1BWP30P140LVT U253 ( .A1(n165), .A2(i_data_bus[164]), .ZN(n359) );
  ND2D1BWP30P140LVT U254 ( .A1(n164), .A2(i_data_bus[69]), .ZN(n350) );
  ND2D1BWP30P140LVT U255 ( .A1(n165), .A2(i_data_bus[165]), .ZN(n351) );
  OAI22D1BWP30P140LVT U256 ( .A1(n269), .A2(n268), .B1(n167), .B2(n267), .ZN(
        n270) );
  ND2D1BWP30P140LVT U257 ( .A1(n164), .A2(i_data_bus[72]), .ZN(n515) );
  ND2D1BWP30P140LVT U258 ( .A1(n165), .A2(i_data_bus[168]), .ZN(n516) );
  ND2D1BWP30P140LVT U259 ( .A1(n164), .A2(i_data_bus[73]), .ZN(n507) );
  ND2D1BWP30P140LVT U260 ( .A1(n165), .A2(i_data_bus[169]), .ZN(n508) );
  ND2D1BWP30P140LVT U261 ( .A1(n164), .A2(i_data_bus[75]), .ZN(n499) );
  ND2D1BWP30P140LVT U262 ( .A1(n165), .A2(i_data_bus[171]), .ZN(n500) );
  ND2D1BWP30P140LVT U263 ( .A1(n165), .A2(i_data_bus[186]), .ZN(n294) );
  ND2D1BWP30P140LVT U264 ( .A1(n165), .A2(i_data_bus[187]), .ZN(n434) );
  ND2D1BWP30P140LVT U265 ( .A1(n165), .A2(i_data_bus[188]), .ZN(n426) );
  ND2D1BWP30P140LVT U266 ( .A1(n164), .A2(i_data_bus[93]), .ZN(n417) );
  ND2D1BWP30P140LVT U267 ( .A1(n165), .A2(i_data_bus[189]), .ZN(n418) );
  ND2OPTIBD1BWP30P140LVT U268 ( .A1(n410), .A2(n409), .ZN(n411) );
  ND2OPTIBD1BWP30P140LVT U269 ( .A1(n172), .A2(i_data_bus[222]), .ZN(n409) );
  ND2OPTIBD1BWP30P140LVT U270 ( .A1(n523), .A2(i_data_bus[254]), .ZN(n410) );
  OAI22D1BWP30P140LVT U271 ( .A1(n408), .A2(n407), .B1(n406), .B2(n405), .ZN(
        n412) );
  INVD1BWP30P140LVT U272 ( .I(i_data_bus[94]), .ZN(n407) );
  INVD1BWP30P140LVT U273 ( .I(i_data_bus[190]), .ZN(n405) );
  ND2D1BWP30P140LVT U274 ( .A1(n164), .A2(i_data_bus[95]), .ZN(n397) );
  ND2D1BWP30P140LVT U275 ( .A1(n165), .A2(i_data_bus[191]), .ZN(n398) );
  ND2D1BWP30P140LVT U276 ( .A1(i_en), .A2(i_valid[4]), .ZN(n209) );
  AOI21D1BWP30P140LVT U277 ( .A1(i_data_bus[38]), .A2(n162), .B(n201), .ZN(
        n262) );
  AOI21D1BWP30P140LVT U278 ( .A1(i_data_bus[42]), .A2(n162), .B(n202), .ZN(
        n283) );
  AOI21D1BWP30P140LVT U279 ( .A1(i_data_bus[44]), .A2(n162), .B(n203), .ZN(
        n498) );
  ND2OPTIBD4BWP30P140LVT U280 ( .A1(n246), .A2(n245), .ZN(n167) );
  NR3D3BWP30P140LVT U281 ( .A1(rst), .A2(i_cmd[7]), .A3(n169), .ZN(n168) );
  OR2D4BWP30P140LVT U282 ( .A1(n261), .A2(n260), .Z(n173) );
  CKAN2D1BWP30P140LVT U283 ( .A1(n257), .A2(n206), .Z(n170) );
  CKAN2D1BWP30P140LVT U284 ( .A1(n524), .A2(i_data_bus[120]), .Z(n174) );
  CKAN2D1BWP30P140LVT U285 ( .A1(n524), .A2(i_data_bus[122]), .Z(n175) );
  CKAN2D1BWP30P140LVT U286 ( .A1(n524), .A2(i_data_bus[113]), .Z(n176) );
  CKAN2D1BWP30P140LVT U287 ( .A1(n524), .A2(i_data_bus[118]), .Z(n177) );
  CKAN2D1BWP30P140LVT U288 ( .A1(n524), .A2(i_data_bus[121]), .Z(n178) );
  CKAN2D1BWP30P140LVT U289 ( .A1(n524), .A2(i_data_bus[111]), .Z(n179) );
  CKAN2D1BWP30P140LVT U290 ( .A1(n524), .A2(i_data_bus[117]), .Z(n180) );
  CKAN2D1BWP30P140LVT U291 ( .A1(n524), .A2(i_data_bus[116]), .Z(n181) );
  CKAN2D1BWP30P140LVT U292 ( .A1(n524), .A2(i_data_bus[100]), .Z(n182) );
  CKAN2D1BWP30P140LVT U293 ( .A1(n524), .A2(i_data_bus[99]), .Z(n183) );
  CKAN2D1BWP30P140LVT U294 ( .A1(n524), .A2(i_data_bus[98]), .Z(n184) );
  CKAN2D1BWP30P140LVT U295 ( .A1(n524), .A2(i_data_bus[97]), .Z(n185) );
  CKAN2D1BWP30P140LVT U296 ( .A1(n524), .A2(i_data_bus[96]), .Z(n186) );
  CKAN2D1BWP30P140LVT U297 ( .A1(n524), .A2(i_data_bus[127]), .Z(n187) );
  CKAN2D1BWP30P140LVT U298 ( .A1(n524), .A2(i_data_bus[126]), .Z(n188) );
  CKAN2D1BWP30P140LVT U299 ( .A1(n524), .A2(i_data_bus[125]), .Z(n189) );
  CKAN2D1BWP30P140LVT U300 ( .A1(n524), .A2(i_data_bus[124]), .Z(n190) );
  CKAN2D1BWP30P140LVT U301 ( .A1(n524), .A2(i_data_bus[123]), .Z(n191) );
  CKAN2D1BWP30P140LVT U302 ( .A1(n524), .A2(i_data_bus[119]), .Z(n192) );
  CKAN2D1BWP30P140LVT U303 ( .A1(n524), .A2(i_data_bus[115]), .Z(n193) );
  CKAN2D1BWP30P140LVT U304 ( .A1(n524), .A2(i_data_bus[114]), .Z(n194) );
  CKAN2D1BWP30P140LVT U305 ( .A1(n524), .A2(i_data_bus[112]), .Z(n195) );
  CKAN2D1BWP30P140LVT U306 ( .A1(n524), .A2(i_data_bus[110]), .Z(n196) );
  CKAN2D1BWP30P140LVT U307 ( .A1(n524), .A2(i_data_bus[109]), .Z(n197) );
  CKAN2D1BWP30P140LVT U308 ( .A1(n524), .A2(i_data_bus[107]), .Z(n198) );
  CKAN2D1BWP30P140LVT U309 ( .A1(n524), .A2(i_data_bus[105]), .Z(n199) );
  CKAN2D1BWP30P140LVT U310 ( .A1(n524), .A2(i_data_bus[104]), .Z(n200) );
  CKAN2D1BWP30P140LVT U311 ( .A1(n524), .A2(i_data_bus[102]), .Z(n201) );
  CKAN2D1BWP30P140LVT U312 ( .A1(n524), .A2(i_data_bus[106]), .Z(n202) );
  CKAN2D1BWP30P140LVT U313 ( .A1(n524), .A2(i_data_bus[108]), .Z(n203) );
  CKAN2D1BWP30P140LVT U314 ( .A1(n524), .A2(i_data_bus[103]), .Z(n204) );
  CKAN2D1BWP30P140LVT U315 ( .A1(n524), .A2(i_data_bus[101]), .Z(n205) );
  INVD1BWP30P140LVT U316 ( .I(i_cmd[6]), .ZN(n237) );
  CKAN2D1BWP30P140LVT U317 ( .A1(i_valid[1]), .A2(i_cmd[1]), .Z(n206) );
  BUFFD6BWP30P140LVT U318 ( .I(n593), .Z(o_data_bus[0]) );
  BUFFD6BWP30P140LVT U319 ( .I(n592), .Z(o_data_bus[1]) );
  BUFFD6BWP30P140LVT U320 ( .I(n591), .Z(o_data_bus[2]) );
  BUFFD6BWP30P140LVT U321 ( .I(n590), .Z(o_data_bus[3]) );
  BUFFD6BWP30P140LVT U322 ( .I(n589), .Z(o_data_bus[4]) );
  BUFFD6BWP30P140LVT U323 ( .I(n588), .Z(o_data_bus[5]) );
  BUFFD6BWP30P140LVT U324 ( .I(n587), .Z(o_data_bus[6]) );
  BUFFD6BWP30P140LVT U325 ( .I(n586), .Z(o_data_bus[7]) );
  BUFFD6BWP30P140LVT U326 ( .I(n585), .Z(o_data_bus[8]) );
  BUFFD6BWP30P140LVT U327 ( .I(n584), .Z(o_data_bus[9]) );
  BUFFD6BWP30P140LVT U328 ( .I(n583), .Z(o_data_bus[10]) );
  BUFFD6BWP30P140LVT U329 ( .I(n582), .Z(o_data_bus[11]) );
  BUFFD6BWP30P140LVT U330 ( .I(n581), .Z(o_data_bus[12]) );
  BUFFD6BWP30P140LVT U331 ( .I(n580), .Z(o_data_bus[13]) );
  BUFFD6BWP30P140LVT U332 ( .I(n579), .Z(o_data_bus[14]) );
  BUFFD6BWP30P140LVT U333 ( .I(n578), .Z(o_data_bus[15]) );
  BUFFD6BWP30P140LVT U334 ( .I(n577), .Z(o_data_bus[16]) );
  BUFFD6BWP30P140LVT U335 ( .I(n576), .Z(o_data_bus[17]) );
  BUFFD6BWP30P140LVT U336 ( .I(n575), .Z(o_data_bus[18]) );
  BUFFD6BWP30P140LVT U337 ( .I(n574), .Z(o_data_bus[19]) );
  BUFFD6BWP30P140LVT U338 ( .I(n573), .Z(o_data_bus[20]) );
  BUFFD6BWP30P140LVT U339 ( .I(n572), .Z(o_data_bus[21]) );
  BUFFD6BWP30P140LVT U340 ( .I(n571), .Z(o_data_bus[22]) );
  BUFFD6BWP30P140LVT U341 ( .I(n570), .Z(o_data_bus[23]) );
  BUFFD6BWP30P140LVT U342 ( .I(n569), .Z(o_data_bus[24]) );
  BUFFD6BWP30P140LVT U343 ( .I(n568), .Z(o_data_bus[25]) );
  BUFFD6BWP30P140LVT U344 ( .I(n567), .Z(o_data_bus[26]) );
  BUFFD6BWP30P140LVT U345 ( .I(n566), .Z(o_data_bus[27]) );
  BUFFD6BWP30P140LVT U346 ( .I(n565), .Z(o_data_bus[28]) );
  BUFFD6BWP30P140LVT U347 ( .I(n564), .Z(o_data_bus[29]) );
  BUFFD6BWP30P140LVT U348 ( .I(n563), .Z(o_data_bus[30]) );
  BUFFD6BWP30P140LVT U349 ( .I(n562), .Z(o_data_bus[31]) );
  BUFFD6BWP30P140LVT U350 ( .I(n561), .Z(o_valid[0]) );
  ND2OPTIBD1BWP30P140LVT U351 ( .A1(n216), .A2(n213), .ZN(n207) );
  NR2D1BWP30P140LVT U352 ( .A1(n208), .A2(n207), .ZN(n212) );
  NR2D1BWP30P140LVT U353 ( .A1(n210), .A2(n209), .ZN(n211) );
  ND3OPTPAD2BWP30P140LVT U354 ( .A1(n214), .A2(i_en), .A3(n213), .ZN(n218) );
  INVD1BWP30P140LVT U355 ( .I(i_valid[0]), .ZN(n219) );
  NR3D0P7BWP30P140LVT U356 ( .A1(n242), .A2(n219), .A3(i_cmd[4]), .ZN(n220) );
  INR2D1BWP30P140LVT U357 ( .A1(i_data_bus[6]), .B1(n163), .ZN(n223) );
  AOI21D1BWP30P140LVT U358 ( .A1(n171), .A2(i_data_bus[134]), .B(n223), .ZN(
        n264) );
  NR2OPTPAD12BWP30P140LVT U359 ( .A1(i_cmd[5]), .A2(i_cmd[6]), .ZN(n235) );
  ND2OPTPAD4BWP30P140LVT U360 ( .A1(n224), .A2(n235), .ZN(n225) );
  INVD1BWP30P140LVT U361 ( .I(i_cmd[2]), .ZN(n227) );
  NR2D1BWP30P140LVT U362 ( .A1(n227), .A2(i_cmd[3]), .ZN(n229) );
  ND3OPTPAD2BWP30P140LVT U363 ( .A1(n229), .A2(i_valid[2]), .A3(n228), .ZN(
        n230) );
  NR2D3BWP30P140LVT U364 ( .A1(n261), .A2(n230), .ZN(n231) );
  INR2D1BWP30P140LVT U365 ( .A1(i_data_bus[70]), .B1(n408), .ZN(n256) );
  ND3OPTPAD2BWP30P140LVT U366 ( .A1(n235), .A2(i_valid[7]), .A3(i_cmd[7]), 
        .ZN(n236) );
  ND2OPTIBD1BWP30P140LVT U367 ( .A1(n523), .A2(i_data_bus[230]), .ZN(n248) );
  INVD2BWP30P140LVT U368 ( .I(i_cmd[0]), .ZN(n242) );
  INVD1BWP30P140LVT U369 ( .I(i_valid[5]), .ZN(n249) );
  ND3OPTPAD2BWP30P140LVT U370 ( .A1(n250), .A2(n237), .A3(i_cmd[5]), .ZN(n251)
         );
  CKND2D4BWP30P140LVT U371 ( .A1(n253), .A2(n252), .ZN(n406) );
  INR2D1BWP30P140LVT U372 ( .A1(i_data_bus[166]), .B1(n406), .ZN(n254) );
  NR3D0P7BWP30P140LVT U373 ( .A1(n256), .A2(n255), .A3(n254), .ZN(n263) );
  INVD2BWP30P140LVT U374 ( .I(n261), .ZN(n258) );
  NR2D1BWP30P140LVT U375 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n259) );
  ND3D1BWP30P140LVT U376 ( .A1(n264), .A2(n263), .A3(n262), .ZN(N375) );
  INR2D1BWP30P140LVT U377 ( .A1(i_data_bus[7]), .B1(n163), .ZN(n265) );
  AOI21D1BWP30P140LVT U378 ( .A1(n171), .A2(i_data_bus[135]), .B(n265), .ZN(
        n275) );
  INR2D1BWP30P140LVT U379 ( .A1(i_data_bus[71]), .B1(n408), .ZN(n272) );
  INVD1BWP30P140LVT U380 ( .I(i_data_bus[167]), .ZN(n266) );
  NR2D1BWP30P140LVT U381 ( .A1(n406), .A2(n266), .ZN(n271) );
  INVD1BWP30P140LVT U382 ( .I(n523), .ZN(n269) );
  INVD1BWP30P140LVT U383 ( .I(i_data_bus[231]), .ZN(n268) );
  INVD1BWP30P140LVT U384 ( .I(i_data_bus[199]), .ZN(n267) );
  NR3D0P7BWP30P140LVT U385 ( .A1(n272), .A2(n271), .A3(n270), .ZN(n274) );
  AOI21D1BWP30P140LVT U386 ( .A1(i_data_bus[39]), .A2(n162), .B(n204), .ZN(
        n273) );
  ND3D1BWP30P140LVT U387 ( .A1(n275), .A2(n274), .A3(n273), .ZN(N376) );
  IOA21D1BWP30P140LVT U388 ( .A1(n523), .A2(i_data_bus[234]), .B(n276), .ZN(
        n279) );
  IOA21D1BWP30P140LVT U389 ( .A1(n172), .A2(i_data_bus[202]), .B(n277), .ZN(
        n278) );
  NR2D1BWP30P140LVT U390 ( .A1(n279), .A2(n278), .ZN(n282) );
  INR2D1BWP30P140LVT U391 ( .A1(i_data_bus[10]), .B1(n163), .ZN(n280) );
  AOI21D1BWP30P140LVT U392 ( .A1(n171), .A2(i_data_bus[138]), .B(n280), .ZN(
        n281) );
  ND3D1BWP30P140LVT U393 ( .A1(n283), .A2(n282), .A3(n281), .ZN(N379) );
  AOI21D1BWP30P140LVT U394 ( .A1(i_data_bus[56]), .A2(n162), .B(n174), .ZN(
        n292) );
  INVD4BWP30P140LVT U395 ( .I(n408), .ZN(n481) );
  ND2OPTIBD1BWP30P140LVT U396 ( .A1(n481), .A2(i_data_bus[88]), .ZN(n284) );
  IOA21D1BWP30P140LVT U397 ( .A1(n523), .A2(i_data_bus[248]), .B(n284), .ZN(
        n287) );
  INVD3BWP30P140LVT U398 ( .I(n406), .ZN(n483) );
  ND2OPTIBD1BWP30P140LVT U399 ( .A1(n483), .A2(i_data_bus[184]), .ZN(n285) );
  IOA21D1BWP30P140LVT U400 ( .A1(n172), .A2(i_data_bus[216]), .B(n285), .ZN(
        n286) );
  NR2D1BWP30P140LVT U401 ( .A1(n287), .A2(n286), .ZN(n291) );
  INR2D1BWP30P140LVT U402 ( .A1(i_data_bus[24]), .B1(n163), .ZN(n289) );
  AOI21D1BWP30P140LVT U403 ( .A1(n171), .A2(i_data_bus[152]), .B(n289), .ZN(
        n290) );
  ND3D1BWP30P140LVT U404 ( .A1(n292), .A2(n291), .A3(n290), .ZN(N393) );
  AOI21D1BWP30P140LVT U405 ( .A1(i_data_bus[58]), .A2(n162), .B(n175), .ZN(
        n300) );
  ND2OPTIBD1BWP30P140LVT U406 ( .A1(n164), .A2(i_data_bus[90]), .ZN(n293) );
  IOA21D1BWP30P140LVT U407 ( .A1(n523), .A2(i_data_bus[250]), .B(n293), .ZN(
        n296) );
  IOA21D1BWP30P140LVT U408 ( .A1(n172), .A2(i_data_bus[218]), .B(n294), .ZN(
        n295) );
  NR2D1BWP30P140LVT U409 ( .A1(n296), .A2(n295), .ZN(n299) );
  INR2D1BWP30P140LVT U410 ( .A1(i_data_bus[26]), .B1(n163), .ZN(n297) );
  AOI21D1BWP30P140LVT U411 ( .A1(n171), .A2(i_data_bus[154]), .B(n297), .ZN(
        n298) );
  ND3D1BWP30P140LVT U412 ( .A1(n300), .A2(n299), .A3(n298), .ZN(N395) );
  AOI21D1BWP30P140LVT U413 ( .A1(i_data_bus[49]), .A2(n162), .B(n176), .ZN(
        n308) );
  ND2OPTIBD1BWP30P140LVT U414 ( .A1(n481), .A2(i_data_bus[81]), .ZN(n301) );
  IOA21D1BWP30P140LVT U415 ( .A1(n523), .A2(i_data_bus[241]), .B(n301), .ZN(
        n304) );
  ND2OPTIBD1BWP30P140LVT U416 ( .A1(n483), .A2(i_data_bus[177]), .ZN(n302) );
  IOA21D1BWP30P140LVT U417 ( .A1(n172), .A2(i_data_bus[209]), .B(n302), .ZN(
        n303) );
  NR2D1BWP30P140LVT U418 ( .A1(n304), .A2(n303), .ZN(n307) );
  INR2D1BWP30P140LVT U419 ( .A1(i_data_bus[17]), .B1(n163), .ZN(n305) );
  AOI21D1BWP30P140LVT U420 ( .A1(n171), .A2(i_data_bus[145]), .B(n305), .ZN(
        n306) );
  ND3D1BWP30P140LVT U421 ( .A1(n308), .A2(n307), .A3(n306), .ZN(N386) );
  AOI21D1BWP30P140LVT U422 ( .A1(i_data_bus[54]), .A2(n162), .B(n177), .ZN(
        n316) );
  ND2OPTIBD1BWP30P140LVT U423 ( .A1(n481), .A2(i_data_bus[86]), .ZN(n309) );
  IOA21D1BWP30P140LVT U424 ( .A1(n523), .A2(i_data_bus[246]), .B(n309), .ZN(
        n312) );
  ND2OPTIBD1BWP30P140LVT U425 ( .A1(n483), .A2(i_data_bus[182]), .ZN(n310) );
  IOA21D1BWP30P140LVT U426 ( .A1(n172), .A2(i_data_bus[214]), .B(n310), .ZN(
        n311) );
  NR2D1BWP30P140LVT U427 ( .A1(n312), .A2(n311), .ZN(n315) );
  INR2D1BWP30P140LVT U428 ( .A1(i_data_bus[22]), .B1(n163), .ZN(n313) );
  AOI21D1BWP30P140LVT U429 ( .A1(n171), .A2(i_data_bus[150]), .B(n313), .ZN(
        n314) );
  ND3D1BWP30P140LVT U430 ( .A1(n316), .A2(n315), .A3(n314), .ZN(N391) );
  AOI21D1BWP30P140LVT U431 ( .A1(i_data_bus[57]), .A2(n162), .B(n178), .ZN(
        n324) );
  ND2OPTIBD1BWP30P140LVT U432 ( .A1(n481), .A2(i_data_bus[89]), .ZN(n317) );
  IOA21D1BWP30P140LVT U433 ( .A1(n523), .A2(i_data_bus[249]), .B(n317), .ZN(
        n320) );
  ND2OPTIBD1BWP30P140LVT U434 ( .A1(n483), .A2(i_data_bus[185]), .ZN(n318) );
  IOA21D1BWP30P140LVT U435 ( .A1(n172), .A2(i_data_bus[217]), .B(n318), .ZN(
        n319) );
  NR2D1BWP30P140LVT U436 ( .A1(n320), .A2(n319), .ZN(n323) );
  INR2D1BWP30P140LVT U437 ( .A1(i_data_bus[25]), .B1(n163), .ZN(n321) );
  AOI21D1BWP30P140LVT U438 ( .A1(n171), .A2(i_data_bus[153]), .B(n321), .ZN(
        n322) );
  ND3D1BWP30P140LVT U439 ( .A1(n324), .A2(n323), .A3(n322), .ZN(N394) );
  AOI21D1BWP30P140LVT U440 ( .A1(i_data_bus[47]), .A2(n162), .B(n179), .ZN(
        n332) );
  ND2OPTIBD1BWP30P140LVT U441 ( .A1(n481), .A2(i_data_bus[79]), .ZN(n325) );
  IOA21D1BWP30P140LVT U442 ( .A1(n523), .A2(i_data_bus[239]), .B(n325), .ZN(
        n328) );
  ND2OPTIBD1BWP30P140LVT U443 ( .A1(n483), .A2(i_data_bus[175]), .ZN(n326) );
  IOA21D1BWP30P140LVT U444 ( .A1(n172), .A2(i_data_bus[207]), .B(n326), .ZN(
        n327) );
  NR2D1BWP30P140LVT U445 ( .A1(n328), .A2(n327), .ZN(n331) );
  INR2D1BWP30P140LVT U446 ( .A1(i_data_bus[15]), .B1(n163), .ZN(n329) );
  AOI21D1BWP30P140LVT U447 ( .A1(n171), .A2(i_data_bus[143]), .B(n329), .ZN(
        n330) );
  ND3D1BWP30P140LVT U448 ( .A1(n332), .A2(n331), .A3(n330), .ZN(N384) );
  AOI21D1BWP30P140LVT U449 ( .A1(i_data_bus[53]), .A2(n162), .B(n180), .ZN(
        n340) );
  ND2OPTIBD1BWP30P140LVT U450 ( .A1(n481), .A2(i_data_bus[85]), .ZN(n333) );
  IOA21D1BWP30P140LVT U451 ( .A1(n523), .A2(i_data_bus[245]), .B(n333), .ZN(
        n336) );
  ND2OPTIBD1BWP30P140LVT U452 ( .A1(n483), .A2(i_data_bus[181]), .ZN(n334) );
  IOA21D1BWP30P140LVT U453 ( .A1(n172), .A2(i_data_bus[213]), .B(n334), .ZN(
        n335) );
  NR2D1BWP30P140LVT U454 ( .A1(n336), .A2(n335), .ZN(n339) );
  INR2D1BWP30P140LVT U455 ( .A1(i_data_bus[21]), .B1(n163), .ZN(n337) );
  AOI21D1BWP30P140LVT U456 ( .A1(n171), .A2(i_data_bus[149]), .B(n337), .ZN(
        n338) );
  ND3D1BWP30P140LVT U457 ( .A1(n340), .A2(n339), .A3(n338), .ZN(N390) );
  AOI21D1BWP30P140LVT U458 ( .A1(i_data_bus[52]), .A2(n162), .B(n181), .ZN(
        n348) );
  ND2OPTIBD1BWP30P140LVT U459 ( .A1(n481), .A2(i_data_bus[84]), .ZN(n341) );
  IOA21D1BWP30P140LVT U460 ( .A1(n523), .A2(i_data_bus[244]), .B(n341), .ZN(
        n344) );
  ND2OPTIBD1BWP30P140LVT U461 ( .A1(n483), .A2(i_data_bus[180]), .ZN(n342) );
  IOA21D1BWP30P140LVT U462 ( .A1(n172), .A2(i_data_bus[212]), .B(n342), .ZN(
        n343) );
  NR2D1BWP30P140LVT U463 ( .A1(n344), .A2(n343), .ZN(n347) );
  INR2D1BWP30P140LVT U464 ( .A1(i_data_bus[20]), .B1(n163), .ZN(n345) );
  AOI21D1BWP30P140LVT U465 ( .A1(n171), .A2(i_data_bus[148]), .B(n345), .ZN(
        n346) );
  ND3D1BWP30P140LVT U466 ( .A1(n348), .A2(n347), .A3(n346), .ZN(N389) );
  INR2D1BWP30P140LVT U467 ( .A1(i_data_bus[5]), .B1(n163), .ZN(n349) );
  AOI21D1BWP30P140LVT U468 ( .A1(n171), .A2(i_data_bus[133]), .B(n349), .ZN(
        n356) );
  IOA21D1BWP30P140LVT U469 ( .A1(n523), .A2(i_data_bus[229]), .B(n350), .ZN(
        n353) );
  IOA21D1BWP30P140LVT U470 ( .A1(n172), .A2(i_data_bus[197]), .B(n351), .ZN(
        n352) );
  NR2D1BWP30P140LVT U471 ( .A1(n353), .A2(n352), .ZN(n355) );
  AOI21D1BWP30P140LVT U472 ( .A1(i_data_bus[37]), .A2(n162), .B(n205), .ZN(
        n354) );
  ND3D1BWP30P140LVT U473 ( .A1(n356), .A2(n355), .A3(n354), .ZN(N374) );
  INR2D1BWP30P140LVT U474 ( .A1(i_data_bus[4]), .B1(n163), .ZN(n357) );
  AOI21D1BWP30P140LVT U475 ( .A1(n171), .A2(i_data_bus[132]), .B(n357), .ZN(
        n364) );
  IOA21D1BWP30P140LVT U476 ( .A1(n523), .A2(i_data_bus[228]), .B(n358), .ZN(
        n361) );
  IOA21D1BWP30P140LVT U477 ( .A1(n172), .A2(i_data_bus[196]), .B(n359), .ZN(
        n360) );
  NR2D1BWP30P140LVT U478 ( .A1(n361), .A2(n360), .ZN(n363) );
  AOI21D1BWP30P140LVT U479 ( .A1(i_data_bus[36]), .A2(n162), .B(n182), .ZN(
        n362) );
  ND3D1BWP30P140LVT U480 ( .A1(n364), .A2(n363), .A3(n362), .ZN(N373) );
  INR2D1BWP30P140LVT U481 ( .A1(i_data_bus[3]), .B1(n163), .ZN(n365) );
  AOI21D1BWP30P140LVT U482 ( .A1(n171), .A2(i_data_bus[131]), .B(n365), .ZN(
        n372) );
  IOA21D1BWP30P140LVT U483 ( .A1(n523), .A2(i_data_bus[227]), .B(n366), .ZN(
        n369) );
  IOA21D1BWP30P140LVT U484 ( .A1(n172), .A2(i_data_bus[195]), .B(n367), .ZN(
        n368) );
  NR2D1BWP30P140LVT U485 ( .A1(n369), .A2(n368), .ZN(n371) );
  AOI21D1BWP30P140LVT U486 ( .A1(i_data_bus[35]), .A2(n162), .B(n183), .ZN(
        n370) );
  ND3D1BWP30P140LVT U487 ( .A1(n372), .A2(n371), .A3(n370), .ZN(N372) );
  INR2D1BWP30P140LVT U488 ( .A1(i_data_bus[2]), .B1(n163), .ZN(n373) );
  AOI21D1BWP30P140LVT U489 ( .A1(n171), .A2(i_data_bus[130]), .B(n373), .ZN(
        n380) );
  IOA21D1BWP30P140LVT U490 ( .A1(n523), .A2(i_data_bus[226]), .B(n374), .ZN(
        n377) );
  IOA21D1BWP30P140LVT U491 ( .A1(n172), .A2(i_data_bus[194]), .B(n375), .ZN(
        n376) );
  NR2D1BWP30P140LVT U492 ( .A1(n377), .A2(n376), .ZN(n379) );
  AOI21D1BWP30P140LVT U493 ( .A1(i_data_bus[34]), .A2(n162), .B(n184), .ZN(
        n378) );
  ND3D1BWP30P140LVT U494 ( .A1(n380), .A2(n379), .A3(n378), .ZN(N371) );
  INR2D1BWP30P140LVT U495 ( .A1(i_data_bus[1]), .B1(n163), .ZN(n381) );
  AOI21D1BWP30P140LVT U496 ( .A1(n171), .A2(i_data_bus[129]), .B(n381), .ZN(
        n388) );
  IOA21D1BWP30P140LVT U497 ( .A1(n523), .A2(i_data_bus[225]), .B(n382), .ZN(
        n385) );
  IOA21D1BWP30P140LVT U498 ( .A1(n172), .A2(i_data_bus[193]), .B(n383), .ZN(
        n384) );
  NR2D1BWP30P140LVT U499 ( .A1(n385), .A2(n384), .ZN(n387) );
  AOI21D1BWP30P140LVT U500 ( .A1(i_data_bus[33]), .A2(n162), .B(n185), .ZN(
        n386) );
  ND3D1BWP30P140LVT U501 ( .A1(n388), .A2(n387), .A3(n386), .ZN(N370) );
  INR2D1BWP30P140LVT U502 ( .A1(i_data_bus[0]), .B1(n163), .ZN(n389) );
  AOI21D1BWP30P140LVT U503 ( .A1(n171), .A2(i_data_bus[128]), .B(n389), .ZN(
        n396) );
  IOA21D1BWP30P140LVT U504 ( .A1(n523), .A2(i_data_bus[224]), .B(n390), .ZN(
        n393) );
  IOA21D1BWP30P140LVT U505 ( .A1(n172), .A2(i_data_bus[192]), .B(n391), .ZN(
        n392) );
  NR2D1BWP30P140LVT U506 ( .A1(n393), .A2(n392), .ZN(n395) );
  AOI21D1BWP30P140LVT U507 ( .A1(i_data_bus[32]), .A2(n162), .B(n186), .ZN(
        n394) );
  ND3D1BWP30P140LVT U508 ( .A1(n396), .A2(n395), .A3(n394), .ZN(N369) );
  AOI21D1BWP30P140LVT U509 ( .A1(i_data_bus[63]), .A2(n162), .B(n187), .ZN(
        n404) );
  IOA21D1BWP30P140LVT U510 ( .A1(n523), .A2(i_data_bus[255]), .B(n397), .ZN(
        n400) );
  IOA21D1BWP30P140LVT U511 ( .A1(n172), .A2(i_data_bus[223]), .B(n398), .ZN(
        n399) );
  NR2D1BWP30P140LVT U512 ( .A1(n400), .A2(n399), .ZN(n403) );
  INR2D1BWP30P140LVT U513 ( .A1(i_data_bus[31]), .B1(n163), .ZN(n401) );
  AOI21D1BWP30P140LVT U514 ( .A1(n171), .A2(i_data_bus[159]), .B(n401), .ZN(
        n402) );
  ND3D1BWP30P140LVT U515 ( .A1(n404), .A2(n403), .A3(n402), .ZN(N400) );
  AOI21D1BWP30P140LVT U516 ( .A1(i_data_bus[62]), .A2(n162), .B(n188), .ZN(
        n416) );
  NR2D1BWP30P140LVT U517 ( .A1(n412), .A2(n411), .ZN(n415) );
  INR2D1BWP30P140LVT U518 ( .A1(i_data_bus[30]), .B1(n163), .ZN(n413) );
  AOI21D1BWP30P140LVT U519 ( .A1(n171), .A2(i_data_bus[158]), .B(n413), .ZN(
        n414) );
  ND3D1BWP30P140LVT U520 ( .A1(n416), .A2(n415), .A3(n414), .ZN(N399) );
  AOI21D1BWP30P140LVT U521 ( .A1(i_data_bus[61]), .A2(n162), .B(n189), .ZN(
        n424) );
  IOA21D1BWP30P140LVT U522 ( .A1(n523), .A2(i_data_bus[253]), .B(n417), .ZN(
        n420) );
  IOA21D1BWP30P140LVT U523 ( .A1(n172), .A2(i_data_bus[221]), .B(n418), .ZN(
        n419) );
  NR2D1BWP30P140LVT U524 ( .A1(n420), .A2(n419), .ZN(n423) );
  INR2D1BWP30P140LVT U525 ( .A1(i_data_bus[29]), .B1(n163), .ZN(n421) );
  AOI21D1BWP30P140LVT U526 ( .A1(n171), .A2(i_data_bus[157]), .B(n421), .ZN(
        n422) );
  ND3D1BWP30P140LVT U527 ( .A1(n424), .A2(n423), .A3(n422), .ZN(N398) );
  AOI21D1BWP30P140LVT U528 ( .A1(i_data_bus[60]), .A2(n162), .B(n190), .ZN(
        n432) );
  ND2OPTIBD1BWP30P140LVT U529 ( .A1(n164), .A2(i_data_bus[92]), .ZN(n425) );
  IOA21D1BWP30P140LVT U530 ( .A1(n523), .A2(i_data_bus[252]), .B(n425), .ZN(
        n428) );
  IOA21D1BWP30P140LVT U531 ( .A1(n172), .A2(i_data_bus[220]), .B(n426), .ZN(
        n427) );
  NR2D1BWP30P140LVT U532 ( .A1(n428), .A2(n427), .ZN(n431) );
  INR2D1BWP30P140LVT U533 ( .A1(i_data_bus[28]), .B1(n163), .ZN(n429) );
  AOI21D1BWP30P140LVT U534 ( .A1(n171), .A2(i_data_bus[156]), .B(n429), .ZN(
        n430) );
  ND3D1BWP30P140LVT U535 ( .A1(n432), .A2(n431), .A3(n430), .ZN(N397) );
  AOI21D1BWP30P140LVT U536 ( .A1(i_data_bus[59]), .A2(n162), .B(n191), .ZN(
        n440) );
  ND2OPTIBD1BWP30P140LVT U537 ( .A1(n164), .A2(i_data_bus[91]), .ZN(n433) );
  IOA21D1BWP30P140LVT U538 ( .A1(n523), .A2(i_data_bus[251]), .B(n433), .ZN(
        n436) );
  IOA21D1BWP30P140LVT U539 ( .A1(n172), .A2(i_data_bus[219]), .B(n434), .ZN(
        n435) );
  NR2D1BWP30P140LVT U540 ( .A1(n436), .A2(n435), .ZN(n439) );
  INR2D1BWP30P140LVT U541 ( .A1(i_data_bus[27]), .B1(n163), .ZN(n437) );
  AOI21D1BWP30P140LVT U542 ( .A1(n171), .A2(i_data_bus[155]), .B(n437), .ZN(
        n438) );
  ND3D1BWP30P140LVT U543 ( .A1(n440), .A2(n439), .A3(n438), .ZN(N396) );
  AOI21D1BWP30P140LVT U544 ( .A1(i_data_bus[55]), .A2(n162), .B(n192), .ZN(
        n448) );
  ND2OPTIBD1BWP30P140LVT U545 ( .A1(n481), .A2(i_data_bus[87]), .ZN(n441) );
  IOA21D1BWP30P140LVT U546 ( .A1(n523), .A2(i_data_bus[247]), .B(n441), .ZN(
        n444) );
  ND2OPTIBD1BWP30P140LVT U547 ( .A1(n483), .A2(i_data_bus[183]), .ZN(n442) );
  IOA21D1BWP30P140LVT U548 ( .A1(n172), .A2(i_data_bus[215]), .B(n442), .ZN(
        n443) );
  NR2D1BWP30P140LVT U549 ( .A1(n444), .A2(n443), .ZN(n447) );
  INR2D1BWP30P140LVT U550 ( .A1(i_data_bus[23]), .B1(n163), .ZN(n445) );
  AOI21D1BWP30P140LVT U551 ( .A1(n171), .A2(i_data_bus[151]), .B(n445), .ZN(
        n446) );
  ND3D1BWP30P140LVT U552 ( .A1(n448), .A2(n447), .A3(n446), .ZN(N392) );
  AOI21D1BWP30P140LVT U553 ( .A1(i_data_bus[51]), .A2(n162), .B(n193), .ZN(
        n456) );
  ND2OPTIBD1BWP30P140LVT U554 ( .A1(n481), .A2(i_data_bus[83]), .ZN(n449) );
  IOA21D1BWP30P140LVT U555 ( .A1(n523), .A2(i_data_bus[243]), .B(n449), .ZN(
        n452) );
  ND2OPTIBD1BWP30P140LVT U556 ( .A1(n483), .A2(i_data_bus[179]), .ZN(n450) );
  IOA21D1BWP30P140LVT U557 ( .A1(n172), .A2(i_data_bus[211]), .B(n450), .ZN(
        n451) );
  NR2D1BWP30P140LVT U558 ( .A1(n452), .A2(n451), .ZN(n455) );
  INR2D1BWP30P140LVT U559 ( .A1(i_data_bus[19]), .B1(n163), .ZN(n453) );
  AOI21D1BWP30P140LVT U560 ( .A1(n171), .A2(i_data_bus[147]), .B(n453), .ZN(
        n454) );
  ND3D1BWP30P140LVT U561 ( .A1(n456), .A2(n455), .A3(n454), .ZN(N388) );
  AOI21D1BWP30P140LVT U562 ( .A1(i_data_bus[50]), .A2(n162), .B(n194), .ZN(
        n464) );
  ND2OPTIBD1BWP30P140LVT U563 ( .A1(n481), .A2(i_data_bus[82]), .ZN(n457) );
  IOA21D1BWP30P140LVT U564 ( .A1(n523), .A2(i_data_bus[242]), .B(n457), .ZN(
        n460) );
  ND2OPTIBD1BWP30P140LVT U565 ( .A1(n483), .A2(i_data_bus[178]), .ZN(n458) );
  IOA21D1BWP30P140LVT U566 ( .A1(n172), .A2(i_data_bus[210]), .B(n458), .ZN(
        n459) );
  NR2D1BWP30P140LVT U567 ( .A1(n460), .A2(n459), .ZN(n463) );
  INR2D1BWP30P140LVT U568 ( .A1(i_data_bus[18]), .B1(n163), .ZN(n461) );
  AOI21D1BWP30P140LVT U569 ( .A1(n171), .A2(i_data_bus[146]), .B(n461), .ZN(
        n462) );
  ND3D1BWP30P140LVT U570 ( .A1(n464), .A2(n463), .A3(n462), .ZN(N387) );
  AOI21D1BWP30P140LVT U571 ( .A1(i_data_bus[48]), .A2(n162), .B(n195), .ZN(
        n472) );
  ND2OPTIBD1BWP30P140LVT U572 ( .A1(n481), .A2(i_data_bus[80]), .ZN(n465) );
  IOA21D1BWP30P140LVT U573 ( .A1(n523), .A2(i_data_bus[240]), .B(n465), .ZN(
        n468) );
  ND2OPTIBD1BWP30P140LVT U574 ( .A1(n483), .A2(i_data_bus[176]), .ZN(n466) );
  IOA21D1BWP30P140LVT U575 ( .A1(n172), .A2(i_data_bus[208]), .B(n466), .ZN(
        n467) );
  NR2D1BWP30P140LVT U576 ( .A1(n468), .A2(n467), .ZN(n471) );
  INR2D1BWP30P140LVT U577 ( .A1(i_data_bus[16]), .B1(n163), .ZN(n469) );
  AOI21D1BWP30P140LVT U578 ( .A1(n171), .A2(i_data_bus[144]), .B(n469), .ZN(
        n470) );
  ND3D1BWP30P140LVT U579 ( .A1(n472), .A2(n471), .A3(n470), .ZN(N385) );
  AOI21D1BWP30P140LVT U580 ( .A1(i_data_bus[46]), .A2(n162), .B(n196), .ZN(
        n480) );
  ND2OPTIBD1BWP30P140LVT U581 ( .A1(n481), .A2(i_data_bus[78]), .ZN(n473) );
  IOA21D1BWP30P140LVT U582 ( .A1(n523), .A2(i_data_bus[238]), .B(n473), .ZN(
        n476) );
  ND2OPTIBD1BWP30P140LVT U583 ( .A1(n483), .A2(i_data_bus[174]), .ZN(n474) );
  IOA21D1BWP30P140LVT U584 ( .A1(n172), .A2(i_data_bus[206]), .B(n474), .ZN(
        n475) );
  NR2D1BWP30P140LVT U585 ( .A1(n476), .A2(n475), .ZN(n479) );
  INR2D1BWP30P140LVT U586 ( .A1(i_data_bus[14]), .B1(n163), .ZN(n477) );
  AOI21D1BWP30P140LVT U587 ( .A1(n171), .A2(i_data_bus[142]), .B(n477), .ZN(
        n478) );
  ND3D1BWP30P140LVT U588 ( .A1(n480), .A2(n479), .A3(n478), .ZN(N383) );
  AOI21D1BWP30P140LVT U589 ( .A1(i_data_bus[45]), .A2(n162), .B(n197), .ZN(
        n490) );
  ND2OPTIBD1BWP30P140LVT U590 ( .A1(n481), .A2(i_data_bus[77]), .ZN(n482) );
  IOA21D1BWP30P140LVT U591 ( .A1(n523), .A2(i_data_bus[237]), .B(n482), .ZN(
        n486) );
  ND2OPTIBD1BWP30P140LVT U592 ( .A1(n483), .A2(i_data_bus[173]), .ZN(n484) );
  IOA21D1BWP30P140LVT U593 ( .A1(n172), .A2(i_data_bus[205]), .B(n484), .ZN(
        n485) );
  NR2D1BWP30P140LVT U594 ( .A1(n486), .A2(n485), .ZN(n489) );
  INR2D1BWP30P140LVT U595 ( .A1(i_data_bus[13]), .B1(n163), .ZN(n487) );
  AOI21D1BWP30P140LVT U596 ( .A1(n171), .A2(i_data_bus[141]), .B(n487), .ZN(
        n488) );
  ND3D1BWP30P140LVT U597 ( .A1(n490), .A2(n489), .A3(n488), .ZN(N382) );
  IOA21D1BWP30P140LVT U598 ( .A1(n523), .A2(i_data_bus[236]), .B(n491), .ZN(
        n494) );
  IOA21D1BWP30P140LVT U599 ( .A1(n172), .A2(i_data_bus[204]), .B(n492), .ZN(
        n493) );
  NR2D1BWP30P140LVT U600 ( .A1(n494), .A2(n493), .ZN(n497) );
  INR2D1BWP30P140LVT U601 ( .A1(i_data_bus[12]), .B1(n163), .ZN(n495) );
  AOI21D1BWP30P140LVT U602 ( .A1(n171), .A2(i_data_bus[140]), .B(n495), .ZN(
        n496) );
  ND3D1BWP30P140LVT U603 ( .A1(n498), .A2(n497), .A3(n496), .ZN(N381) );
  AOI21D1BWP30P140LVT U604 ( .A1(i_data_bus[43]), .A2(n162), .B(n198), .ZN(
        n506) );
  IOA21D1BWP30P140LVT U605 ( .A1(n523), .A2(i_data_bus[235]), .B(n499), .ZN(
        n502) );
  IOA21D1BWP30P140LVT U606 ( .A1(n172), .A2(i_data_bus[203]), .B(n500), .ZN(
        n501) );
  NR2D1BWP30P140LVT U607 ( .A1(n502), .A2(n501), .ZN(n505) );
  INR2D1BWP30P140LVT U608 ( .A1(i_data_bus[11]), .B1(n163), .ZN(n503) );
  AOI21D1BWP30P140LVT U609 ( .A1(n171), .A2(i_data_bus[139]), .B(n503), .ZN(
        n504) );
  ND3D1BWP30P140LVT U610 ( .A1(n506), .A2(n505), .A3(n504), .ZN(N380) );
  AOI21D1BWP30P140LVT U611 ( .A1(i_data_bus[41]), .A2(n162), .B(n199), .ZN(
        n514) );
  IOA21D1BWP30P140LVT U612 ( .A1(n523), .A2(i_data_bus[233]), .B(n507), .ZN(
        n510) );
  IOA21D1BWP30P140LVT U613 ( .A1(n172), .A2(i_data_bus[201]), .B(n508), .ZN(
        n509) );
  NR2D1BWP30P140LVT U614 ( .A1(n510), .A2(n509), .ZN(n513) );
  INR2D1BWP30P140LVT U615 ( .A1(i_data_bus[9]), .B1(n163), .ZN(n511) );
  AOI21D1BWP30P140LVT U616 ( .A1(n171), .A2(i_data_bus[137]), .B(n511), .ZN(
        n512) );
  ND3D1BWP30P140LVT U617 ( .A1(n514), .A2(n513), .A3(n512), .ZN(N378) );
  AOI21D1BWP30P140LVT U618 ( .A1(i_data_bus[40]), .A2(n162), .B(n200), .ZN(
        n522) );
  IOA21D1BWP30P140LVT U619 ( .A1(n523), .A2(i_data_bus[232]), .B(n515), .ZN(
        n518) );
  IOA21D1BWP30P140LVT U620 ( .A1(n172), .A2(i_data_bus[200]), .B(n516), .ZN(
        n517) );
  NR2D1BWP30P140LVT U621 ( .A1(n518), .A2(n517), .ZN(n521) );
  INR2D1BWP30P140LVT U622 ( .A1(i_data_bus[8]), .B1(n163), .ZN(n519) );
  AOI21D1BWP30P140LVT U623 ( .A1(n171), .A2(i_data_bus[136]), .B(n519), .ZN(
        n520) );
  ND3D1BWP30P140LVT U624 ( .A1(n522), .A2(n521), .A3(n520), .ZN(N377) );
  NR4D0BWP30P140LVT U625 ( .A1(n164), .A2(n172), .A3(n165), .A4(n523), .ZN(
        n527) );
  NR2D1BWP30P140LVT U626 ( .A1(n162), .A2(n524), .ZN(n526) );
  INVD1BWP30P140LVT U627 ( .I(n171), .ZN(n525) );
  ND4D1BWP30P140LVT U628 ( .A1(n527), .A2(n526), .A3(n525), .A4(n163), .ZN(
        N402) );
endmodule

