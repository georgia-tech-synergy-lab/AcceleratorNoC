

    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_0 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD6BWP30P140LVT U3 ( .I(n267), .ZN(n280) );
  INVD6BWP30P140LVT U4 ( .I(n123), .ZN(n261) );
  INVD3BWP30P140LVT U5 ( .I(n57), .ZN(n1) );
  INVD3BWP30P140LVT U6 ( .I(n122), .ZN(n2) );
  MOAI22D1BWP30P140LVT U7 ( .A1(n280), .A2(n3), .B1(n2), .B2(i_data_bus[174]), 
        .ZN(n268) );
  INVD1BWP30P140LVT U8 ( .I(i_data_bus[206]), .ZN(n3) );
  INVD6BWP30P140LVT U9 ( .I(n16), .ZN(n267) );
  INVD4BWP30P140LVT U10 ( .I(n2), .ZN(n278) );
  INVD2BWP30P140LVT U11 ( .I(n31), .ZN(n156) );
  ND2OPTIBD1BWP30P140LVT U12 ( .A1(n40), .A2(n7), .ZN(n32) );
  ND2D1BWP30P140LVT U13 ( .A1(n28), .A2(n27), .ZN(n38) );
  INVD1BWP30P140LVT U14 ( .I(n9), .ZN(n61) );
  INVD1BWP30P140LVT U15 ( .I(n156), .ZN(n252) );
  INVD1BWP30P140LVT U16 ( .I(n156), .ZN(n276) );
  ND2D1BWP30P140LVT U17 ( .A1(n6), .A2(n37), .ZN(n43) );
  INVD1BWP30P140LVT U18 ( .I(n139), .ZN(n269) );
  ND2D1BWP30P140LVT U19 ( .A1(n41), .A2(n40), .ZN(n48) );
  AOI21D1BWP30P140LVT U20 ( .A1(n282), .A2(i_data_bus[229]), .B(n117), .ZN(
        n119) );
  AOI21D1BWP30P140LVT U21 ( .A1(n282), .A2(i_data_bus[237]), .B(n281), .ZN(
        n285) );
  INR2D1BWP30P140LVT U22 ( .A1(n45), .B1(n44), .ZN(n155) );
  INVD1BWP30P140LVT U23 ( .I(i_cmd[0]), .ZN(n27) );
  INR3D0BWP30P140LVT U24 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n27), .ZN(n8)
         );
  INVD1BWP30P140LVT U25 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U26 ( .A1(n4), .A2(i_en), .ZN(n10) );
  NR2OPTPAD1BWP30P140LVT U27 ( .A1(i_cmd[5]), .A2(n10), .ZN(n5) );
  OR2D2BWP30P140LVT U28 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n18) );
  INR2D2BWP30P140LVT U29 ( .A1(n5), .B1(n18), .ZN(n40) );
  INVD1BWP30P140LVT U30 ( .I(i_cmd[3]), .ZN(n6) );
  INVD1BWP30P140LVT U31 ( .I(i_cmd[2]), .ZN(n37) );
  NR2D1BWP30P140LVT U32 ( .A1(n43), .A2(i_cmd[1]), .ZN(n7) );
  INR2D1BWP30P140LVT U33 ( .A1(n8), .B1(n32), .ZN(n9) );
  INVD2BWP30P140LVT U34 ( .I(n61), .ZN(n255) );
  OR2D4BWP30P140LVT U35 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n26) );
  NR3D0P7BWP30P140LVT U36 ( .A1(n26), .A2(i_cmd[3]), .A3(i_cmd[0]), .ZN(n12)
         );
  NR2D1BWP30P140LVT U37 ( .A1(i_cmd[4]), .A2(n10), .ZN(n11) );
  ND2OPTIBD2BWP30P140LVT U38 ( .A1(n12), .A2(n11), .ZN(n22) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(i_cmd[6]), .A2(i_valid[6]), .ZN(n14) );
  NR2D1BWP30P140LVT U40 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n13) );
  IND2D1BWP30P140LVT U41 ( .A1(n14), .B1(n13), .ZN(n15) );
  OR2D2BWP30P140LVT U42 ( .A1(n22), .A2(n15), .Z(n16) );
  ND2OPTIBD1BWP30P140LVT U43 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n17) );
  NR2D1BWP30P140LVT U44 ( .A1(n18), .A2(n17), .ZN(n19) );
  INVD1BWP30P140LVT U45 ( .I(n19), .ZN(n20) );
  OR2D4BWP30P140LVT U46 ( .A1(n22), .A2(n20), .Z(n122) );
  INVD1BWP30P140LVT U47 ( .I(i_cmd[7]), .ZN(n21) );
  INR4D0BWP30P140LVT U48 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n21), .ZN(n23) );
  INR2D1BWP30P140LVT U49 ( .A1(n23), .B1(n22), .ZN(n24) );
  INVD2BWP30P140LVT U50 ( .I(n24), .ZN(n139) );
  INVD2BWP30P140LVT U51 ( .I(n139), .ZN(n282) );
  NR4D0BWP30P140LVT U52 ( .A1(n255), .A2(n267), .A3(n2), .A4(n282), .ZN(n47)
         );
  ND2D1BWP30P140LVT U53 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n25) );
  NR2D1BWP30P140LVT U54 ( .A1(n26), .A2(n25), .ZN(n30) );
  INVD1BWP30P140LVT U55 ( .I(i_cmd[4]), .ZN(n28) );
  INVD1BWP30P140LVT U56 ( .I(n38), .ZN(n29) );
  ND2OPTIBD2BWP30P140LVT U57 ( .A1(n40), .A2(n29), .ZN(n44) );
  INR2D1BWP30P140LVT U58 ( .A1(n30), .B1(n44), .ZN(n31) );
  INVD1BWP30P140LVT U59 ( .I(n156), .ZN(n147) );
  INVD1BWP30P140LVT U60 ( .I(n32), .ZN(n35) );
  ND2OPTIBD1BWP30P140LVT U61 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n33) );
  NR2D1BWP30P140LVT U62 ( .A1(n33), .A2(i_cmd[0]), .ZN(n34) );
  ND2OPTIBD2BWP30P140LVT U63 ( .A1(n35), .A2(n34), .ZN(n49) );
  INVD3BWP30P140LVT U64 ( .I(n49), .ZN(n275) );
  NR2D1BWP30P140LVT U65 ( .A1(n147), .A2(n275), .ZN(n46) );
  NR2D1BWP30P140LVT U66 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .ZN(n36) );
  IND3D1BWP30P140LVT U67 ( .A1(n37), .B1(i_valid[2]), .B2(n36), .ZN(n39) );
  NR2D1BWP30P140LVT U68 ( .A1(n39), .A2(n38), .ZN(n41) );
  ND2D1BWP30P140LVT U69 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n42) );
  NR2D1BWP30P140LVT U70 ( .A1(n43), .A2(n42), .ZN(n45) );
  INVD1BWP30P140LVT U71 ( .I(n155), .ZN(n57) );
  ND4D1BWP30P140LVT U72 ( .A1(n47), .A2(n46), .A3(n48), .A4(n57), .ZN(N402) );
  INVD2BWP30P140LVT U73 ( .I(n48), .ZN(n274) );
  INVD2BWP30P140LVT U74 ( .I(n57), .ZN(n250) );
  AOI22D1BWP30P140LVT U75 ( .A1(n274), .A2(i_data_bus[68]), .B1(n250), .B2(
        i_data_bus[36]), .ZN(n56) );
  INVD2BWP30P140LVT U76 ( .I(n49), .ZN(n251) );
  AOI22D1BWP30P140LVT U77 ( .A1(n252), .A2(i_data_bus[100]), .B1(n251), .B2(
        i_data_bus[132]), .ZN(n55) );
  INVD1BWP30P140LVT U78 ( .I(i_data_bus[164]), .ZN(n51) );
  INVD4BWP30P140LVT U79 ( .I(n267), .ZN(n237) );
  INVD1BWP30P140LVT U80 ( .I(i_data_bus[196]), .ZN(n50) );
  OAI22D1BWP30P140LVT U81 ( .A1(n278), .A2(n51), .B1(n237), .B2(n50), .ZN(n52)
         );
  AOI21OPTREPBD1BWP30P140LVT U82 ( .A1(n282), .A2(i_data_bus[228]), .B(n52), 
        .ZN(n54) );
  ND2D1BWP30P140LVT U83 ( .A1(n255), .A2(i_data_bus[4]), .ZN(n53) );
  ND4D1BWP30P140LVT U84 ( .A1(n56), .A2(n55), .A3(n54), .A4(n53), .ZN(N373) );
  AOI22D1BWP30P140LVT U85 ( .A1(n274), .A2(i_data_bus[95]), .B1(n1), .B2(
        i_data_bus[63]), .ZN(n65) );
  AOI22D1BWP30P140LVT U86 ( .A1(n147), .A2(i_data_bus[127]), .B1(n275), .B2(
        i_data_bus[159]), .ZN(n64) );
  INVD1BWP30P140LVT U87 ( .I(i_data_bus[223]), .ZN(n59) );
  INVD1BWP30P140LVT U88 ( .I(i_data_bus[191]), .ZN(n58) );
  OAI22D1BWP30P140LVT U89 ( .A1(n237), .A2(n59), .B1(n122), .B2(n58), .ZN(n60)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n282), .A2(i_data_bus[255]), .B(n60), .ZN(n63)
         );
  INVD2BWP30P140LVT U91 ( .I(n61), .ZN(n283) );
  ND2D1BWP30P140LVT U92 ( .A1(n283), .A2(i_data_bus[31]), .ZN(n62) );
  ND4D1BWP30P140LVT U93 ( .A1(n65), .A2(n64), .A3(n63), .A4(n62), .ZN(N400) );
  AOI22D1BWP30P140LVT U94 ( .A1(n274), .A2(i_data_bus[94]), .B1(n1), .B2(
        i_data_bus[62]), .ZN(n72) );
  AOI22D1BWP30P140LVT U95 ( .A1(n147), .A2(i_data_bus[126]), .B1(n275), .B2(
        i_data_bus[158]), .ZN(n71) );
  INVD1BWP30P140LVT U96 ( .I(n139), .ZN(n134) );
  INVD1BWP30P140LVT U97 ( .I(i_data_bus[222]), .ZN(n67) );
  INVD1BWP30P140LVT U98 ( .I(i_data_bus[190]), .ZN(n66) );
  OAI22D1BWP30P140LVT U99 ( .A1(n237), .A2(n67), .B1(n122), .B2(n66), .ZN(n68)
         );
  AOI21D1BWP30P140LVT U100 ( .A1(n134), .A2(i_data_bus[254]), .B(n68), .ZN(n70) );
  ND2D1BWP30P140LVT U101 ( .A1(n283), .A2(i_data_bus[30]), .ZN(n69) );
  ND4D1BWP30P140LVT U102 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(N399)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n274), .A2(i_data_bus[76]), .B1(n250), .B2(
        i_data_bus[44]), .ZN(n79) );
  AOI22D1BWP30P140LVT U104 ( .A1(n252), .A2(i_data_bus[108]), .B1(n251), .B2(
        i_data_bus[140]), .ZN(n78) );
  INVD1BWP30P140LVT U105 ( .I(i_data_bus[204]), .ZN(n74) );
  INVD1BWP30P140LVT U106 ( .I(i_data_bus[172]), .ZN(n73) );
  OAI22D1BWP30P140LVT U107 ( .A1(n280), .A2(n74), .B1(n278), .B2(n73), .ZN(n75) );
  AOI21D1BWP30P140LVT U108 ( .A1(n282), .A2(i_data_bus[236]), .B(n75), .ZN(n77) );
  ND2D1BWP30P140LVT U109 ( .A1(n255), .A2(i_data_bus[12]), .ZN(n76) );
  ND4D1BWP30P140LVT U110 ( .A1(n79), .A2(n78), .A3(n77), .A4(n76), .ZN(N381)
         );
  AOI22D1BWP30P140LVT U111 ( .A1(n274), .A2(i_data_bus[75]), .B1(n250), .B2(
        i_data_bus[43]), .ZN(n86) );
  AOI22D1BWP30P140LVT U112 ( .A1(n252), .A2(i_data_bus[107]), .B1(n251), .B2(
        i_data_bus[139]), .ZN(n85) );
  INVD1BWP30P140LVT U113 ( .I(i_data_bus[203]), .ZN(n81) );
  INVD1BWP30P140LVT U114 ( .I(i_data_bus[171]), .ZN(n80) );
  OAI22D1BWP30P140LVT U115 ( .A1(n280), .A2(n81), .B1(n278), .B2(n80), .ZN(n82) );
  AOI21D1BWP30P140LVT U116 ( .A1(n282), .A2(i_data_bus[235]), .B(n82), .ZN(n84) );
  ND2D1BWP30P140LVT U117 ( .A1(n255), .A2(i_data_bus[11]), .ZN(n83) );
  ND4D1BWP30P140LVT U118 ( .A1(n86), .A2(n85), .A3(n84), .A4(n83), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U119 ( .A1(n274), .A2(i_data_bus[74]), .B1(n250), .B2(
        i_data_bus[42]), .ZN(n93) );
  AOI22D1BWP30P140LVT U120 ( .A1(n252), .A2(i_data_bus[106]), .B1(n251), .B2(
        i_data_bus[138]), .ZN(n92) );
  INVD1BWP30P140LVT U121 ( .I(i_data_bus[202]), .ZN(n88) );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[170]), .ZN(n87) );
  OAI22D1BWP30P140LVT U123 ( .A1(n280), .A2(n88), .B1(n278), .B2(n87), .ZN(n89) );
  AOI21D1BWP30P140LVT U124 ( .A1(n282), .A2(i_data_bus[234]), .B(n89), .ZN(n91) );
  ND2D1BWP30P140LVT U125 ( .A1(n255), .A2(i_data_bus[10]), .ZN(n90) );
  ND4D1BWP30P140LVT U126 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(N379)
         );
  AOI22D1BWP30P140LVT U127 ( .A1(n274), .A2(i_data_bus[73]), .B1(n250), .B2(
        i_data_bus[41]), .ZN(n100) );
  AOI22D1BWP30P140LVT U128 ( .A1(n252), .A2(i_data_bus[105]), .B1(n251), .B2(
        i_data_bus[137]), .ZN(n99) );
  INVD1BWP30P140LVT U129 ( .I(i_data_bus[201]), .ZN(n95) );
  INVD1BWP30P140LVT U130 ( .I(i_data_bus[169]), .ZN(n94) );
  OAI22D1BWP30P140LVT U131 ( .A1(n280), .A2(n95), .B1(n278), .B2(n94), .ZN(n96) );
  AOI21D1BWP30P140LVT U132 ( .A1(n282), .A2(i_data_bus[233]), .B(n96), .ZN(n98) );
  ND2D1BWP30P140LVT U133 ( .A1(n255), .A2(i_data_bus[9]), .ZN(n97) );
  ND4D1BWP30P140LVT U134 ( .A1(n100), .A2(n99), .A3(n98), .A4(n97), .ZN(N378)
         );
  AOI22D1BWP30P140LVT U135 ( .A1(n274), .A2(i_data_bus[71]), .B1(n250), .B2(
        i_data_bus[39]), .ZN(n107) );
  AOI22D1BWP30P140LVT U136 ( .A1(n252), .A2(i_data_bus[103]), .B1(n251), .B2(
        i_data_bus[135]), .ZN(n106) );
  INVD1BWP30P140LVT U137 ( .I(i_data_bus[199]), .ZN(n102) );
  INVD1BWP30P140LVT U138 ( .I(i_data_bus[167]), .ZN(n101) );
  OAI22D1BWP30P140LVT U139 ( .A1(n280), .A2(n102), .B1(n278), .B2(n101), .ZN(
        n103) );
  AOI21D1BWP30P140LVT U140 ( .A1(n282), .A2(i_data_bus[231]), .B(n103), .ZN(
        n105) );
  ND2D1BWP30P140LVT U141 ( .A1(n255), .A2(i_data_bus[7]), .ZN(n104) );
  ND4D1BWP30P140LVT U142 ( .A1(n107), .A2(n106), .A3(n105), .A4(n104), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U143 ( .A1(n274), .A2(i_data_bus[70]), .B1(n250), .B2(
        i_data_bus[38]), .ZN(n114) );
  AOI22D1BWP30P140LVT U144 ( .A1(n252), .A2(i_data_bus[102]), .B1(n251), .B2(
        i_data_bus[134]), .ZN(n113) );
  INVD1BWP30P140LVT U145 ( .I(i_data_bus[198]), .ZN(n109) );
  INVD1BWP30P140LVT U146 ( .I(i_data_bus[166]), .ZN(n108) );
  OAI22D1BWP30P140LVT U147 ( .A1(n280), .A2(n109), .B1(n278), .B2(n108), .ZN(
        n110) );
  AOI21D1BWP30P140LVT U148 ( .A1(n282), .A2(i_data_bus[230]), .B(n110), .ZN(
        n112) );
  ND2D1BWP30P140LVT U149 ( .A1(n255), .A2(i_data_bus[6]), .ZN(n111) );
  ND4D1BWP30P140LVT U150 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U151 ( .A1(n274), .A2(i_data_bus[69]), .B1(n250), .B2(
        i_data_bus[37]), .ZN(n121) );
  AOI22D1BWP30P140LVT U152 ( .A1(n252), .A2(i_data_bus[101]), .B1(n251), .B2(
        i_data_bus[133]), .ZN(n120) );
  INVD1BWP30P140LVT U153 ( .I(i_data_bus[197]), .ZN(n116) );
  INVD1BWP30P140LVT U154 ( .I(i_data_bus[165]), .ZN(n115) );
  OAI22D1BWP30P140LVT U155 ( .A1(n280), .A2(n116), .B1(n278), .B2(n115), .ZN(
        n117) );
  ND2D1BWP30P140LVT U156 ( .A1(n255), .A2(i_data_bus[5]), .ZN(n118) );
  ND4D1BWP30P140LVT U157 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U158 ( .A1(n274), .A2(i_data_bus[93]), .B1(n1), .B2(
        i_data_bus[61]), .ZN(n130) );
  AOI22D1BWP30P140LVT U159 ( .A1(n147), .A2(i_data_bus[125]), .B1(n275), .B2(
        i_data_bus[157]), .ZN(n129) );
  INVD1BWP30P140LVT U160 ( .I(i_data_bus[221]), .ZN(n125) );
  INVD2BWP30P140LVT U161 ( .I(n122), .ZN(n123) );
  INVD1BWP30P140LVT U162 ( .I(i_data_bus[189]), .ZN(n124) );
  OAI22D1BWP30P140LVT U163 ( .A1(n237), .A2(n125), .B1(n261), .B2(n124), .ZN(
        n126) );
  AOI21D1BWP30P140LVT U164 ( .A1(n134), .A2(i_data_bus[253]), .B(n126), .ZN(
        n128) );
  ND2D1BWP30P140LVT U165 ( .A1(n283), .A2(i_data_bus[29]), .ZN(n127) );
  ND4D1BWP30P140LVT U166 ( .A1(n130), .A2(n129), .A3(n128), .A4(n127), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U167 ( .A1(n274), .A2(i_data_bus[92]), .B1(n1), .B2(
        i_data_bus[60]), .ZN(n138) );
  AOI22D1BWP30P140LVT U168 ( .A1(n147), .A2(i_data_bus[124]), .B1(n275), .B2(
        i_data_bus[156]), .ZN(n137) );
  INVD1BWP30P140LVT U169 ( .I(i_data_bus[220]), .ZN(n132) );
  INVD1BWP30P140LVT U170 ( .I(i_data_bus[188]), .ZN(n131) );
  OAI22D1BWP30P140LVT U171 ( .A1(n237), .A2(n132), .B1(n261), .B2(n131), .ZN(
        n133) );
  AOI21D1BWP30P140LVT U172 ( .A1(n134), .A2(i_data_bus[252]), .B(n133), .ZN(
        n136) );
  ND2D1BWP30P140LVT U173 ( .A1(n283), .A2(i_data_bus[28]), .ZN(n135) );
  ND4D1BWP30P140LVT U174 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U175 ( .A1(n274), .A2(i_data_bus[91]), .B1(n1), .B2(
        i_data_bus[59]), .ZN(n146) );
  AOI22D1BWP30P140LVT U176 ( .A1(n147), .A2(i_data_bus[123]), .B1(n275), .B2(
        i_data_bus[155]), .ZN(n145) );
  INVD1BWP30P140LVT U177 ( .I(i_data_bus[219]), .ZN(n141) );
  INVD1BWP30P140LVT U178 ( .I(i_data_bus[187]), .ZN(n140) );
  OAI22D1BWP30P140LVT U179 ( .A1(n237), .A2(n141), .B1(n261), .B2(n140), .ZN(
        n142) );
  AOI21D1BWP30P140LVT U180 ( .A1(n269), .A2(i_data_bus[251]), .B(n142), .ZN(
        n144) );
  ND2D1BWP30P140LVT U181 ( .A1(n283), .A2(i_data_bus[27]), .ZN(n143) );
  ND4D1BWP30P140LVT U182 ( .A1(n146), .A2(n145), .A3(n144), .A4(n143), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U183 ( .A1(n274), .A2(i_data_bus[90]), .B1(n1), .B2(
        i_data_bus[58]), .ZN(n154) );
  AOI22D1BWP30P140LVT U184 ( .A1(n147), .A2(i_data_bus[122]), .B1(n275), .B2(
        i_data_bus[154]), .ZN(n153) );
  INVD1BWP30P140LVT U185 ( .I(i_data_bus[218]), .ZN(n149) );
  INVD1BWP30P140LVT U186 ( .I(i_data_bus[186]), .ZN(n148) );
  OAI22D1BWP30P140LVT U187 ( .A1(n237), .A2(n149), .B1(n261), .B2(n148), .ZN(
        n150) );
  AOI21D1BWP30P140LVT U188 ( .A1(n269), .A2(i_data_bus[250]), .B(n150), .ZN(
        n152) );
  ND2D1BWP30P140LVT U189 ( .A1(n255), .A2(i_data_bus[26]), .ZN(n151) );
  ND4D1BWP30P140LVT U190 ( .A1(n154), .A2(n153), .A3(n152), .A4(n151), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U191 ( .A1(n274), .A2(i_data_bus[89]), .B1(n1), .B2(
        i_data_bus[57]), .ZN(n163) );
  AOI22D1BWP30P140LVT U192 ( .A1(n276), .A2(i_data_bus[121]), .B1(n275), .B2(
        i_data_bus[153]), .ZN(n162) );
  INVD1BWP30P140LVT U193 ( .I(i_data_bus[217]), .ZN(n158) );
  INVD1BWP30P140LVT U194 ( .I(i_data_bus[185]), .ZN(n157) );
  OAI22D1BWP30P140LVT U195 ( .A1(n237), .A2(n158), .B1(n261), .B2(n157), .ZN(
        n159) );
  AOI21D1BWP30P140LVT U196 ( .A1(n269), .A2(i_data_bus[249]), .B(n159), .ZN(
        n161) );
  ND2D1BWP30P140LVT U197 ( .A1(n283), .A2(i_data_bus[25]), .ZN(n160) );
  ND4D1BWP30P140LVT U198 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U199 ( .A1(n274), .A2(i_data_bus[88]), .B1(n1), .B2(
        i_data_bus[56]), .ZN(n170) );
  AOI22D1BWP30P140LVT U200 ( .A1(n276), .A2(i_data_bus[120]), .B1(n275), .B2(
        i_data_bus[152]), .ZN(n169) );
  INVD1BWP30P140LVT U201 ( .I(i_data_bus[216]), .ZN(n165) );
  INVD1BWP30P140LVT U202 ( .I(i_data_bus[184]), .ZN(n164) );
  OAI22D1BWP30P140LVT U203 ( .A1(n280), .A2(n165), .B1(n261), .B2(n164), .ZN(
        n166) );
  AOI21D1BWP30P140LVT U204 ( .A1(n269), .A2(i_data_bus[248]), .B(n166), .ZN(
        n168) );
  ND2D1BWP30P140LVT U205 ( .A1(n283), .A2(i_data_bus[24]), .ZN(n167) );
  ND4D1BWP30P140LVT U206 ( .A1(n170), .A2(n169), .A3(n168), .A4(n167), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U207 ( .A1(n274), .A2(i_data_bus[87]), .B1(n1), .B2(
        i_data_bus[55]), .ZN(n177) );
  AOI22D1BWP30P140LVT U208 ( .A1(n276), .A2(i_data_bus[119]), .B1(n275), .B2(
        i_data_bus[151]), .ZN(n176) );
  INVD1BWP30P140LVT U209 ( .I(i_data_bus[215]), .ZN(n172) );
  INVD1BWP30P140LVT U210 ( .I(i_data_bus[183]), .ZN(n171) );
  OAI22D1BWP30P140LVT U211 ( .A1(n280), .A2(n172), .B1(n261), .B2(n171), .ZN(
        n173) );
  AOI21D1BWP30P140LVT U212 ( .A1(n269), .A2(i_data_bus[247]), .B(n173), .ZN(
        n175) );
  ND2D1BWP30P140LVT U213 ( .A1(n283), .A2(i_data_bus[23]), .ZN(n174) );
  ND4D1BWP30P140LVT U214 ( .A1(n177), .A2(n176), .A3(n175), .A4(n174), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U215 ( .A1(n274), .A2(i_data_bus[86]), .B1(n1), .B2(
        i_data_bus[54]), .ZN(n184) );
  AOI22D1BWP30P140LVT U216 ( .A1(n276), .A2(i_data_bus[118]), .B1(n275), .B2(
        i_data_bus[150]), .ZN(n183) );
  INVD1BWP30P140LVT U217 ( .I(i_data_bus[214]), .ZN(n179) );
  INVD1BWP30P140LVT U218 ( .I(i_data_bus[182]), .ZN(n178) );
  OAI22D1BWP30P140LVT U219 ( .A1(n280), .A2(n179), .B1(n261), .B2(n178), .ZN(
        n180) );
  AOI21D1BWP30P140LVT U220 ( .A1(n269), .A2(i_data_bus[246]), .B(n180), .ZN(
        n182) );
  ND2D1BWP30P140LVT U221 ( .A1(n283), .A2(i_data_bus[22]), .ZN(n181) );
  ND4D1BWP30P140LVT U222 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U223 ( .A1(n274), .A2(i_data_bus[85]), .B1(n1), .B2(
        i_data_bus[53]), .ZN(n191) );
  AOI22D1BWP30P140LVT U224 ( .A1(n276), .A2(i_data_bus[117]), .B1(n275), .B2(
        i_data_bus[149]), .ZN(n190) );
  INVD1BWP30P140LVT U225 ( .I(i_data_bus[213]), .ZN(n186) );
  INVD1BWP30P140LVT U226 ( .I(i_data_bus[181]), .ZN(n185) );
  OAI22D1BWP30P140LVT U227 ( .A1(n280), .A2(n186), .B1(n261), .B2(n185), .ZN(
        n187) );
  AOI21D1BWP30P140LVT U228 ( .A1(n269), .A2(i_data_bus[245]), .B(n187), .ZN(
        n189) );
  ND2D1BWP30P140LVT U229 ( .A1(n283), .A2(i_data_bus[21]), .ZN(n188) );
  ND4D1BWP30P140LVT U230 ( .A1(n191), .A2(n190), .A3(n189), .A4(n188), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U231 ( .A1(n274), .A2(i_data_bus[84]), .B1(n1), .B2(
        i_data_bus[52]), .ZN(n198) );
  AOI22D1BWP30P140LVT U232 ( .A1(n276), .A2(i_data_bus[116]), .B1(n275), .B2(
        i_data_bus[148]), .ZN(n197) );
  INVD1BWP30P140LVT U233 ( .I(i_data_bus[212]), .ZN(n193) );
  INVD1BWP30P140LVT U234 ( .I(i_data_bus[180]), .ZN(n192) );
  OAI22D1BWP30P140LVT U235 ( .A1(n280), .A2(n193), .B1(n261), .B2(n192), .ZN(
        n194) );
  AOI21D1BWP30P140LVT U236 ( .A1(n269), .A2(i_data_bus[244]), .B(n194), .ZN(
        n196) );
  ND2D1BWP30P140LVT U237 ( .A1(n283), .A2(i_data_bus[20]), .ZN(n195) );
  ND4D1BWP30P140LVT U238 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U239 ( .A1(n274), .A2(i_data_bus[83]), .B1(n1), .B2(
        i_data_bus[51]), .ZN(n205) );
  AOI22D1BWP30P140LVT U240 ( .A1(n276), .A2(i_data_bus[115]), .B1(n275), .B2(
        i_data_bus[147]), .ZN(n204) );
  INVD1BWP30P140LVT U241 ( .I(i_data_bus[211]), .ZN(n200) );
  INVD1BWP30P140LVT U242 ( .I(i_data_bus[179]), .ZN(n199) );
  OAI22D1BWP30P140LVT U243 ( .A1(n280), .A2(n200), .B1(n261), .B2(n199), .ZN(
        n201) );
  AOI21D1BWP30P140LVT U244 ( .A1(n269), .A2(i_data_bus[243]), .B(n201), .ZN(
        n203) );
  ND2D1BWP30P140LVT U245 ( .A1(n283), .A2(i_data_bus[19]), .ZN(n202) );
  ND4D1BWP30P140LVT U246 ( .A1(n205), .A2(n204), .A3(n203), .A4(n202), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U247 ( .A1(n274), .A2(i_data_bus[82]), .B1(n1), .B2(
        i_data_bus[50]), .ZN(n211) );
  AOI22D1BWP30P140LVT U248 ( .A1(n276), .A2(i_data_bus[114]), .B1(n275), .B2(
        i_data_bus[146]), .ZN(n210) );
  INVD1BWP30P140LVT U249 ( .I(i_data_bus[178]), .ZN(n206) );
  MOAI22D1BWP30P140LVT U250 ( .A1(n261), .A2(n206), .B1(n267), .B2(
        i_data_bus[210]), .ZN(n207) );
  AOI21D1BWP30P140LVT U251 ( .A1(n269), .A2(i_data_bus[242]), .B(n207), .ZN(
        n209) );
  ND2D1BWP30P140LVT U252 ( .A1(n283), .A2(i_data_bus[18]), .ZN(n208) );
  ND4D1BWP30P140LVT U253 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U254 ( .A1(n274), .A2(i_data_bus[67]), .B1(n250), .B2(
        i_data_bus[35]), .ZN(n217) );
  AOI22D1BWP30P140LVT U255 ( .A1(n252), .A2(i_data_bus[99]), .B1(n251), .B2(
        i_data_bus[131]), .ZN(n216) );
  INVD1BWP30P140LVT U256 ( .I(i_data_bus[163]), .ZN(n212) );
  MOAI22D1BWP30P140LVT U257 ( .A1(n278), .A2(n212), .B1(n267), .B2(
        i_data_bus[195]), .ZN(n213) );
  AOI21D1BWP30P140LVT U258 ( .A1(n282), .A2(i_data_bus[227]), .B(n213), .ZN(
        n215) );
  ND2D1BWP30P140LVT U259 ( .A1(n255), .A2(i_data_bus[3]), .ZN(n214) );
  ND4D1BWP30P140LVT U260 ( .A1(n217), .A2(n216), .A3(n215), .A4(n214), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U261 ( .A1(n274), .A2(i_data_bus[81]), .B1(n1), .B2(
        i_data_bus[49]), .ZN(n223) );
  AOI22D1BWP30P140LVT U262 ( .A1(n276), .A2(i_data_bus[113]), .B1(n275), .B2(
        i_data_bus[145]), .ZN(n222) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[177]), .ZN(n218) );
  MOAI22D1BWP30P140LVT U264 ( .A1(n261), .A2(n218), .B1(n267), .B2(
        i_data_bus[209]), .ZN(n219) );
  AOI21D1BWP30P140LVT U265 ( .A1(n269), .A2(i_data_bus[241]), .B(n219), .ZN(
        n221) );
  ND2D1BWP30P140LVT U266 ( .A1(n283), .A2(i_data_bus[17]), .ZN(n220) );
  ND4D1BWP30P140LVT U267 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U268 ( .A1(n274), .A2(i_data_bus[80]), .B1(n1), .B2(
        i_data_bus[48]), .ZN(n229) );
  AOI22D1BWP30P140LVT U269 ( .A1(n276), .A2(i_data_bus[112]), .B1(n275), .B2(
        i_data_bus[144]), .ZN(n228) );
  INVD1BWP30P140LVT U270 ( .I(i_data_bus[176]), .ZN(n224) );
  MOAI22D1BWP30P140LVT U271 ( .A1(n261), .A2(n224), .B1(n267), .B2(
        i_data_bus[208]), .ZN(n225) );
  AOI21D1BWP30P140LVT U272 ( .A1(n269), .A2(i_data_bus[240]), .B(n225), .ZN(
        n227) );
  ND2D1BWP30P140LVT U273 ( .A1(n283), .A2(i_data_bus[16]), .ZN(n226) );
  ND4D1BWP30P140LVT U274 ( .A1(n229), .A2(n228), .A3(n227), .A4(n226), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U275 ( .A1(n274), .A2(i_data_bus[66]), .B1(n250), .B2(
        i_data_bus[34]), .ZN(n235) );
  AOI22D1BWP30P140LVT U276 ( .A1(n252), .A2(i_data_bus[98]), .B1(n251), .B2(
        i_data_bus[130]), .ZN(n234) );
  INVD1BWP30P140LVT U277 ( .I(i_data_bus[162]), .ZN(n230) );
  MOAI22D1BWP30P140LVT U278 ( .A1(n278), .A2(n230), .B1(n267), .B2(
        i_data_bus[194]), .ZN(n231) );
  AOI21D1BWP30P140LVT U279 ( .A1(n282), .A2(i_data_bus[226]), .B(n231), .ZN(
        n233) );
  ND2D1BWP30P140LVT U280 ( .A1(n255), .A2(i_data_bus[2]), .ZN(n232) );
  ND4D1BWP30P140LVT U281 ( .A1(n235), .A2(n234), .A3(n233), .A4(n232), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U282 ( .A1(n274), .A2(i_data_bus[65]), .B1(n250), .B2(
        i_data_bus[33]), .ZN(n243) );
  AOI22D1BWP30P140LVT U283 ( .A1(n252), .A2(i_data_bus[97]), .B1(n251), .B2(
        i_data_bus[129]), .ZN(n242) );
  INVD1BWP30P140LVT U284 ( .I(i_data_bus[161]), .ZN(n238) );
  INVD1BWP30P140LVT U285 ( .I(i_data_bus[193]), .ZN(n236) );
  OAI22D1BWP30P140LVT U286 ( .A1(n278), .A2(n238), .B1(n237), .B2(n236), .ZN(
        n239) );
  AOI21OPTREPBD1BWP30P140LVT U287 ( .A1(n282), .A2(i_data_bus[225]), .B(n239), 
        .ZN(n241) );
  ND2D1BWP30P140LVT U288 ( .A1(n255), .A2(i_data_bus[1]), .ZN(n240) );
  ND4D1BWP30P140LVT U289 ( .A1(n243), .A2(n242), .A3(n241), .A4(n240), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U290 ( .A1(n274), .A2(i_data_bus[72]), .B1(n250), .B2(
        i_data_bus[40]), .ZN(n249) );
  AOI22D1BWP30P140LVT U291 ( .A1(n252), .A2(i_data_bus[104]), .B1(n251), .B2(
        i_data_bus[136]), .ZN(n248) );
  INVD1BWP30P140LVT U292 ( .I(i_data_bus[168]), .ZN(n244) );
  MOAI22D1BWP30P140LVT U293 ( .A1(n278), .A2(n244), .B1(n267), .B2(
        i_data_bus[200]), .ZN(n245) );
  AOI21D1BWP30P140LVT U294 ( .A1(n269), .A2(i_data_bus[232]), .B(n245), .ZN(
        n247) );
  ND2D1BWP30P140LVT U295 ( .A1(n255), .A2(i_data_bus[8]), .ZN(n246) );
  ND4D1BWP30P140LVT U296 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U297 ( .A1(n274), .A2(i_data_bus[64]), .B1(n250), .B2(
        i_data_bus[32]), .ZN(n259) );
  AOI22D1BWP30P140LVT U298 ( .A1(n252), .A2(i_data_bus[96]), .B1(n251), .B2(
        i_data_bus[128]), .ZN(n258) );
  INR2D1BWP30P140LVT U299 ( .A1(i_data_bus[192]), .B1(n280), .ZN(n254) );
  INR2D1BWP30P140LVT U300 ( .A1(i_data_bus[160]), .B1(n278), .ZN(n253) );
  AOI211D1BWP30P140LVT U301 ( .A1(i_data_bus[224]), .A2(n282), .B(n254), .C(
        n253), .ZN(n257) );
  ND2D1BWP30P140LVT U302 ( .A1(n255), .A2(i_data_bus[0]), .ZN(n256) );
  ND4D1BWP30P140LVT U303 ( .A1(n259), .A2(n258), .A3(n257), .A4(n256), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U304 ( .A1(n274), .A2(i_data_bus[79]), .B1(n1), .B2(
        i_data_bus[47]), .ZN(n266) );
  AOI22D1BWP30P140LVT U305 ( .A1(n276), .A2(i_data_bus[111]), .B1(n275), .B2(
        i_data_bus[143]), .ZN(n265) );
  INVD1BWP30P140LVT U306 ( .I(i_data_bus[175]), .ZN(n260) );
  MOAI22D1BWP30P140LVT U307 ( .A1(n261), .A2(n260), .B1(n267), .B2(
        i_data_bus[207]), .ZN(n262) );
  AOI21D1BWP30P140LVT U308 ( .A1(n269), .A2(i_data_bus[239]), .B(n262), .ZN(
        n264) );
  ND2D1BWP30P140LVT U309 ( .A1(n283), .A2(i_data_bus[15]), .ZN(n263) );
  ND4D1BWP30P140LVT U310 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U311 ( .A1(n274), .A2(i_data_bus[78]), .B1(n1), .B2(
        i_data_bus[46]), .ZN(n273) );
  AOI22D1BWP30P140LVT U312 ( .A1(n276), .A2(i_data_bus[110]), .B1(n275), .B2(
        i_data_bus[142]), .ZN(n272) );
  AOI21D1BWP30P140LVT U313 ( .A1(n269), .A2(i_data_bus[238]), .B(n268), .ZN(
        n271) );
  ND2D1BWP30P140LVT U314 ( .A1(n283), .A2(i_data_bus[14]), .ZN(n270) );
  ND4D1BWP30P140LVT U315 ( .A1(n273), .A2(n272), .A3(n271), .A4(n270), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U316 ( .A1(n274), .A2(i_data_bus[77]), .B1(n1), .B2(
        i_data_bus[45]), .ZN(n287) );
  AOI22D1BWP30P140LVT U317 ( .A1(n276), .A2(i_data_bus[109]), .B1(n275), .B2(
        i_data_bus[141]), .ZN(n286) );
  INVD1BWP30P140LVT U318 ( .I(i_data_bus[205]), .ZN(n279) );
  INVD1BWP30P140LVT U319 ( .I(i_data_bus[173]), .ZN(n277) );
  OAI22D1BWP30P140LVT U320 ( .A1(n280), .A2(n279), .B1(n278), .B2(n277), .ZN(
        n281) );
  ND2D1BWP30P140LVT U321 ( .A1(n283), .A2(i_data_bus[13]), .ZN(n284) );
  ND4D1BWP30P140LVT U322 ( .A1(n287), .A2(n286), .A3(n285), .A4(n284), .ZN(
        N382) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_9 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_10 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_11 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_12 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_13 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_14 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_15 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_9 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_10 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_11 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_12 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_13 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_14 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_15 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_9 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n211), .ZN(n1) );
  INVD4BWP30P140LVT U4 ( .I(n68), .ZN(n2) );
  ND2D1BWP30P140LVT U5 ( .A1(n2), .A2(i_data_bus[0]), .ZN(n256) );
  INR2D2BWP30P140LVT U6 ( .A1(n45), .B1(n44), .ZN(n284) );
  OR2D1BWP30P140LVT U7 ( .A1(n12), .A2(n28), .Z(n22) );
  ND2D1BWP30P140LVT U8 ( .A1(n11), .A2(n10), .ZN(n12) );
  CKBD1BWP30P140LVT U9 ( .I(n153), .Z(n288) );
  ND2D1BWP30P140LVT U10 ( .A1(n34), .A2(n33), .ZN(n48) );
  ND2D1BWP30P140LVT U11 ( .A1(n42), .A2(n7), .ZN(n49) );
  NR2D1BWP30P140LVT U12 ( .A1(n22), .A2(n20), .ZN(n21) );
  INVD1BWP30P140LVT U13 ( .I(n59), .ZN(n68) );
  OR3D1BWP30P140LVT U14 ( .A1(n40), .A2(n49), .A3(n39), .Z(n73) );
  INVD1BWP30P140LVT U15 ( .I(n37), .ZN(n177) );
  INVD1BWP30P140LVT U16 ( .I(n153), .ZN(n64) );
  ND2D1BWP30P140LVT U17 ( .A1(n26), .A2(n25), .ZN(n211) );
  BUFFD2BWP30P140LVT U18 ( .I(n284), .Z(n274) );
  INR2D4BWP30P140LVT U19 ( .A1(n52), .B1(n51), .ZN(n283) );
  INVD1BWP30P140LVT U20 ( .I(i_cmd[0]), .ZN(n33) );
  INR3D0BWP30P140LVT U21 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n33), .ZN(n3)
         );
  INVD1BWP30P140LVT U22 ( .I(n3), .ZN(n8) );
  OR2D4BWP30P140LVT U23 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n31) );
  NR2D1BWP30P140LVT U24 ( .A1(n31), .A2(i_cmd[5]), .ZN(n6) );
  INVD1BWP30P140LVT U25 ( .I(rst), .ZN(n4) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n4), .A2(i_en), .Z(n9) );
  INR2D1BWP30P140LVT U27 ( .A1(n9), .B1(i_cmd[1]), .ZN(n5) );
  ND2OPTIBD1BWP30P140LVT U28 ( .A1(n6), .A2(n5), .ZN(n39) );
  INVD1BWP30P140LVT U29 ( .I(i_cmd[2]), .ZN(n42) );
  INVD1BWP30P140LVT U30 ( .I(i_cmd[3]), .ZN(n7) );
  NR3D0P7BWP30P140LVT U31 ( .A1(n8), .A2(n39), .A3(n49), .ZN(n59) );
  NR2D1BWP30P140LVT U32 ( .A1(i_cmd[3]), .A2(i_cmd[4]), .ZN(n11) );
  INVD1BWP30P140LVT U33 ( .I(n9), .ZN(n29) );
  NR2D1BWP30P140LVT U34 ( .A1(i_cmd[0]), .A2(n29), .ZN(n10) );
  OR2D1BWP30P140LVT U35 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n28) );
  CKAN2D1BWP30P140LVT U36 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n14) );
  NR2D1BWP30P140LVT U37 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .ZN(n13) );
  ND2OPTIBD1BWP30P140LVT U38 ( .A1(n14), .A2(n13), .ZN(n15) );
  NR2OPTPAD1BWP30P140LVT U39 ( .A1(n22), .A2(n15), .ZN(n16) );
  INVD2BWP30P140LVT U40 ( .I(n16), .ZN(n207) );
  INVD2BWP30P140LVT U41 ( .I(n207), .ZN(n275) );
  INVD1BWP30P140LVT U42 ( .I(i_valid[5]), .ZN(n17) );
  IND2D1BWP30P140LVT U43 ( .A1(n17), .B1(i_cmd[5]), .ZN(n18) );
  NR2OPTPAD1BWP30P140LVT U44 ( .A1(n31), .A2(n18), .ZN(n19) );
  INVD1BWP30P140LVT U45 ( .I(n19), .ZN(n20) );
  INVD2BWP30P140LVT U46 ( .I(n21), .ZN(n153) );
  INVD1BWP30P140LVT U47 ( .I(n22), .ZN(n26) );
  INVD1BWP30P140LVT U48 ( .I(i_valid[7]), .ZN(n24) );
  INVD1BWP30P140LVT U49 ( .I(i_cmd[7]), .ZN(n23) );
  NR4D0BWP30P140LVT U50 ( .A1(n24), .A2(n23), .A3(i_cmd[6]), .A4(i_cmd[5]), 
        .ZN(n25) );
  NR4D0BWP30P140LVT U51 ( .A1(n59), .A2(n275), .A3(n64), .A4(n1), .ZN(n55) );
  ND2D1BWP30P140LVT U52 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n27) );
  NR2D1BWP30P140LVT U53 ( .A1(n28), .A2(n27), .ZN(n36) );
  NR2D1BWP30P140LVT U54 ( .A1(i_cmd[5]), .A2(n29), .ZN(n30) );
  INVD1BWP30P140LVT U55 ( .I(n30), .ZN(n32) );
  NR2OPTPAD1BWP30P140LVT U56 ( .A1(n32), .A2(n31), .ZN(n52) );
  INVD1BWP30P140LVT U57 ( .I(i_cmd[4]), .ZN(n34) );
  INVD1BWP30P140LVT U58 ( .I(n48), .ZN(n35) );
  ND2OPTIBD2BWP30P140LVT U59 ( .A1(n52), .A2(n35), .ZN(n44) );
  INR2D1BWP30P140LVT U60 ( .A1(n36), .B1(n44), .ZN(n37) );
  INVD1BWP30P140LVT U61 ( .I(n177), .ZN(n169) );
  ND2D1BWP30P140LVT U62 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n38) );
  OR2D1BWP30P140LVT U63 ( .A1(n38), .A2(i_cmd[0]), .Z(n40) );
  INVD3BWP30P140LVT U64 ( .I(n73), .ZN(n285) );
  NR2D1BWP30P140LVT U65 ( .A1(n169), .A2(n285), .ZN(n54) );
  NR2D1BWP30P140LVT U66 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .ZN(n41) );
  ND2D1BWP30P140LVT U67 ( .A1(n41), .A2(i_valid[2]), .ZN(n43) );
  NR2D1BWP30P140LVT U68 ( .A1(n43), .A2(n42), .ZN(n45) );
  INVD1BWP30P140LVT U69 ( .I(n284), .ZN(n46) );
  INVD1BWP30P140LVT U70 ( .I(n46), .ZN(n168) );
  ND2D1BWP30P140LVT U71 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n47) );
  NR3D0P7BWP30P140LVT U72 ( .A1(n49), .A2(n48), .A3(n47), .ZN(n50) );
  INVD1BWP30P140LVT U73 ( .I(n50), .ZN(n51) );
  NR2D1BWP30P140LVT U74 ( .A1(n168), .A2(n283), .ZN(n53) );
  ND3D1BWP30P140LVT U75 ( .A1(n55), .A2(n54), .A3(n53), .ZN(N402) );
  AOI22D1BWP30P140LVT U76 ( .A1(n168), .A2(i_data_bus[95]), .B1(n283), .B2(
        i_data_bus[63]), .ZN(n63) );
  AOI22D1BWP30P140LVT U77 ( .A1(n169), .A2(i_data_bus[127]), .B1(n285), .B2(
        i_data_bus[159]), .ZN(n62) );
  BUFFD4BWP30P140LVT U78 ( .I(n207), .Z(n290) );
  INVD1BWP30P140LVT U79 ( .I(i_data_bus[223]), .ZN(n57) );
  ND2D1BWP30P140LVT U80 ( .A1(n64), .A2(i_data_bus[191]), .ZN(n56) );
  OAI21D1BWP30P140LVT U81 ( .A1(n290), .A2(n57), .B(n56), .ZN(n58) );
  AOI21D1BWP30P140LVT U82 ( .A1(n1), .A2(i_data_bus[255]), .B(n58), .ZN(n61)
         );
  ND2D1BWP30P140LVT U83 ( .A1(n2), .A2(i_data_bus[31]), .ZN(n60) );
  ND4D1BWP30P140LVT U84 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(N400) );
  AOI22D1BWP30P140LVT U85 ( .A1(n168), .A2(i_data_bus[94]), .B1(n283), .B2(
        i_data_bus[62]), .ZN(n72) );
  AOI22D1BWP30P140LVT U86 ( .A1(n169), .A2(i_data_bus[126]), .B1(n285), .B2(
        i_data_bus[158]), .ZN(n71) );
  INVD1BWP30P140LVT U87 ( .I(i_data_bus[222]), .ZN(n66) );
  ND2D1BWP30P140LVT U88 ( .A1(n64), .A2(i_data_bus[190]), .ZN(n65) );
  OAI21D1BWP30P140LVT U89 ( .A1(n290), .A2(n66), .B(n65), .ZN(n67) );
  AOI21D1BWP30P140LVT U90 ( .A1(n1), .A2(i_data_bus[254]), .B(n67), .ZN(n70)
         );
  ND2D1BWP30P140LVT U91 ( .A1(n2), .A2(i_data_bus[30]), .ZN(n69) );
  ND4D1BWP30P140LVT U92 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(N399) );
  AOI22D1BWP30P140LVT U93 ( .A1(n274), .A2(i_data_bus[72]), .B1(n283), .B2(
        i_data_bus[40]), .ZN(n82) );
  INVD2BWP30P140LVT U94 ( .I(n177), .ZN(n267) );
  INVD2BWP30P140LVT U95 ( .I(n73), .ZN(n266) );
  AOI22D1BWP30P140LVT U96 ( .A1(n267), .A2(i_data_bus[104]), .B1(n266), .B2(
        i_data_bus[136]), .ZN(n81) );
  INVD1BWP30P140LVT U97 ( .I(i_data_bus[232]), .ZN(n74) );
  NR2D1BWP30P140LVT U98 ( .A1(n211), .A2(n74), .ZN(n78) );
  INVD2BWP30P140LVT U99 ( .I(n153), .ZN(n75) );
  INVD3BWP30P140LVT U100 ( .I(n75), .ZN(n277) );
  INVD1BWP30P140LVT U101 ( .I(i_data_bus[168]), .ZN(n76) );
  NR2D1BWP30P140LVT U102 ( .A1(n277), .A2(n76), .ZN(n77) );
  AOI211D1BWP30P140LVT U103 ( .A1(n275), .A2(i_data_bus[200]), .B(n78), .C(n77), .ZN(n80) );
  ND2D1BWP30P140LVT U104 ( .A1(n2), .A2(i_data_bus[8]), .ZN(n79) );
  ND4D1BWP30P140LVT U105 ( .A1(n82), .A2(n81), .A3(n80), .A4(n79), .ZN(N377)
         );
  AOI22D1BWP30P140LVT U106 ( .A1(n274), .A2(i_data_bus[76]), .B1(n283), .B2(
        i_data_bus[44]), .ZN(n89) );
  AOI22D1BWP30P140LVT U107 ( .A1(n267), .A2(i_data_bus[108]), .B1(n266), .B2(
        i_data_bus[140]), .ZN(n88) );
  INVD1BWP30P140LVT U108 ( .I(i_data_bus[204]), .ZN(n84) );
  INVD1BWP30P140LVT U109 ( .I(i_data_bus[172]), .ZN(n83) );
  OAI22D1BWP30P140LVT U110 ( .A1(n290), .A2(n84), .B1(n277), .B2(n83), .ZN(n85) );
  AOI21D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[236]), .B(n85), .ZN(n87)
         );
  ND2D1BWP30P140LVT U112 ( .A1(n2), .A2(i_data_bus[12]), .ZN(n86) );
  ND4D1BWP30P140LVT U113 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(N381)
         );
  AOI22D1BWP30P140LVT U114 ( .A1(n274), .A2(i_data_bus[75]), .B1(n283), .B2(
        i_data_bus[43]), .ZN(n96) );
  AOI22D1BWP30P140LVT U115 ( .A1(n267), .A2(i_data_bus[107]), .B1(n266), .B2(
        i_data_bus[139]), .ZN(n95) );
  INVD1BWP30P140LVT U116 ( .I(i_data_bus[203]), .ZN(n91) );
  INVD1BWP30P140LVT U117 ( .I(i_data_bus[171]), .ZN(n90) );
  OAI22D1BWP30P140LVT U118 ( .A1(n290), .A2(n91), .B1(n277), .B2(n90), .ZN(n92) );
  AOI21D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[235]), .B(n92), .ZN(n94)
         );
  ND2D1BWP30P140LVT U120 ( .A1(n2), .A2(i_data_bus[11]), .ZN(n93) );
  ND4D1BWP30P140LVT U121 ( .A1(n96), .A2(n95), .A3(n94), .A4(n93), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U122 ( .A1(n274), .A2(i_data_bus[74]), .B1(n283), .B2(
        i_data_bus[42]), .ZN(n103) );
  AOI22D1BWP30P140LVT U123 ( .A1(n267), .A2(i_data_bus[106]), .B1(n266), .B2(
        i_data_bus[138]), .ZN(n102) );
  INVD1BWP30P140LVT U124 ( .I(i_data_bus[202]), .ZN(n98) );
  INVD1BWP30P140LVT U125 ( .I(i_data_bus[170]), .ZN(n97) );
  OAI22D1BWP30P140LVT U126 ( .A1(n290), .A2(n98), .B1(n277), .B2(n97), .ZN(n99) );
  AOI21D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[234]), .B(n99), .ZN(n101)
         );
  ND2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[10]), .ZN(n100) );
  ND4D1BWP30P140LVT U129 ( .A1(n103), .A2(n102), .A3(n101), .A4(n100), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U130 ( .A1(n274), .A2(i_data_bus[73]), .B1(n283), .B2(
        i_data_bus[41]), .ZN(n110) );
  AOI22D1BWP30P140LVT U131 ( .A1(n267), .A2(i_data_bus[105]), .B1(n266), .B2(
        i_data_bus[137]), .ZN(n109) );
  INVD1BWP30P140LVT U132 ( .I(i_data_bus[201]), .ZN(n105) );
  INVD1BWP30P140LVT U133 ( .I(i_data_bus[169]), .ZN(n104) );
  OAI22D1BWP30P140LVT U134 ( .A1(n290), .A2(n105), .B1(n277), .B2(n104), .ZN(
        n106) );
  AOI21D1BWP30P140LVT U135 ( .A1(n1), .A2(i_data_bus[233]), .B(n106), .ZN(n108) );
  ND2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[9]), .ZN(n107) );
  ND4D1BWP30P140LVT U137 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U138 ( .A1(n274), .A2(i_data_bus[71]), .B1(n283), .B2(
        i_data_bus[39]), .ZN(n117) );
  AOI22D1BWP30P140LVT U139 ( .A1(n267), .A2(i_data_bus[103]), .B1(n266), .B2(
        i_data_bus[135]), .ZN(n116) );
  INVD1BWP30P140LVT U140 ( .I(i_data_bus[199]), .ZN(n112) );
  INVD1BWP30P140LVT U141 ( .I(i_data_bus[167]), .ZN(n111) );
  OAI22D1BWP30P140LVT U142 ( .A1(n290), .A2(n112), .B1(n277), .B2(n111), .ZN(
        n113) );
  AOI21D1BWP30P140LVT U143 ( .A1(n1), .A2(i_data_bus[231]), .B(n113), .ZN(n115) );
  ND2D1BWP30P140LVT U144 ( .A1(n2), .A2(i_data_bus[7]), .ZN(n114) );
  ND4D1BWP30P140LVT U145 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U146 ( .A1(n274), .A2(i_data_bus[70]), .B1(n283), .B2(
        i_data_bus[38]), .ZN(n124) );
  AOI22D1BWP30P140LVT U147 ( .A1(n267), .A2(i_data_bus[102]), .B1(n266), .B2(
        i_data_bus[134]), .ZN(n123) );
  INVD1BWP30P140LVT U148 ( .I(i_data_bus[198]), .ZN(n119) );
  INVD1BWP30P140LVT U149 ( .I(i_data_bus[166]), .ZN(n118) );
  OAI22D1BWP30P140LVT U150 ( .A1(n290), .A2(n119), .B1(n277), .B2(n118), .ZN(
        n120) );
  AOI21D1BWP30P140LVT U151 ( .A1(n1), .A2(i_data_bus[230]), .B(n120), .ZN(n122) );
  ND2D1BWP30P140LVT U152 ( .A1(n2), .A2(i_data_bus[6]), .ZN(n121) );
  ND4D1BWP30P140LVT U153 ( .A1(n124), .A2(n123), .A3(n122), .A4(n121), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U154 ( .A1(n274), .A2(i_data_bus[69]), .B1(n283), .B2(
        i_data_bus[37]), .ZN(n131) );
  AOI22D1BWP30P140LVT U155 ( .A1(n267), .A2(i_data_bus[101]), .B1(n266), .B2(
        i_data_bus[133]), .ZN(n130) );
  INVD1BWP30P140LVT U156 ( .I(i_data_bus[197]), .ZN(n126) );
  INVD1BWP30P140LVT U157 ( .I(i_data_bus[165]), .ZN(n125) );
  OAI22D1BWP30P140LVT U158 ( .A1(n290), .A2(n126), .B1(n288), .B2(n125), .ZN(
        n127) );
  AOI21D1BWP30P140LVT U159 ( .A1(n1), .A2(i_data_bus[229]), .B(n127), .ZN(n129) );
  ND2D1BWP30P140LVT U160 ( .A1(n2), .A2(i_data_bus[5]), .ZN(n128) );
  ND4D1BWP30P140LVT U161 ( .A1(n131), .A2(n130), .A3(n129), .A4(n128), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U162 ( .A1(n274), .A2(i_data_bus[68]), .B1(n283), .B2(
        i_data_bus[36]), .ZN(n137) );
  AOI22D1BWP30P140LVT U163 ( .A1(n267), .A2(i_data_bus[100]), .B1(n266), .B2(
        i_data_bus[132]), .ZN(n136) );
  INVD1BWP30P140LVT U164 ( .I(i_data_bus[164]), .ZN(n132) );
  MOAI22D1BWP30P140LVT U165 ( .A1(n277), .A2(n132), .B1(n275), .B2(
        i_data_bus[196]), .ZN(n133) );
  AOI21D1BWP30P140LVT U166 ( .A1(n1), .A2(i_data_bus[228]), .B(n133), .ZN(n135) );
  ND2D1BWP30P140LVT U167 ( .A1(n2), .A2(i_data_bus[4]), .ZN(n134) );
  ND4D1BWP30P140LVT U168 ( .A1(n137), .A2(n136), .A3(n135), .A4(n134), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U169 ( .A1(n274), .A2(i_data_bus[67]), .B1(n283), .B2(
        i_data_bus[35]), .ZN(n143) );
  AOI22D1BWP30P140LVT U170 ( .A1(n267), .A2(i_data_bus[99]), .B1(n266), .B2(
        i_data_bus[131]), .ZN(n142) );
  INVD1BWP30P140LVT U171 ( .I(i_data_bus[163]), .ZN(n138) );
  MOAI22D1BWP30P140LVT U172 ( .A1(n277), .A2(n138), .B1(n275), .B2(
        i_data_bus[195]), .ZN(n139) );
  AOI21D1BWP30P140LVT U173 ( .A1(n1), .A2(i_data_bus[227]), .B(n139), .ZN(n141) );
  ND2D1BWP30P140LVT U174 ( .A1(n2), .A2(i_data_bus[3]), .ZN(n140) );
  ND4D1BWP30P140LVT U175 ( .A1(n143), .A2(n142), .A3(n141), .A4(n140), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U176 ( .A1(n168), .A2(i_data_bus[93]), .B1(n283), .B2(
        i_data_bus[61]), .ZN(n151) );
  AOI22D1BWP30P140LVT U177 ( .A1(n169), .A2(i_data_bus[125]), .B1(n285), .B2(
        i_data_bus[157]), .ZN(n150) );
  INVD1BWP30P140LVT U178 ( .I(i_data_bus[221]), .ZN(n146) );
  INVD2BWP30P140LVT U179 ( .I(n153), .ZN(n144) );
  INVD3BWP30P140LVT U180 ( .I(n144), .ZN(n248) );
  INVD1BWP30P140LVT U181 ( .I(i_data_bus[189]), .ZN(n145) );
  OAI22D1BWP30P140LVT U182 ( .A1(n290), .A2(n146), .B1(n248), .B2(n145), .ZN(
        n147) );
  AOI21D1BWP30P140LVT U183 ( .A1(n1), .A2(i_data_bus[253]), .B(n147), .ZN(n149) );
  ND2D1BWP30P140LVT U184 ( .A1(n2), .A2(i_data_bus[29]), .ZN(n148) );
  ND4D1BWP30P140LVT U185 ( .A1(n151), .A2(n150), .A3(n149), .A4(n148), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U186 ( .A1(n168), .A2(i_data_bus[92]), .B1(n283), .B2(
        i_data_bus[60]), .ZN(n160) );
  AOI22D1BWP30P140LVT U187 ( .A1(n169), .A2(i_data_bus[124]), .B1(n285), .B2(
        i_data_bus[156]), .ZN(n159) );
  INVD1BWP30P140LVT U188 ( .I(i_data_bus[188]), .ZN(n152) );
  OR2D1BWP30P140LVT U189 ( .A1(n153), .A2(n152), .Z(n155) );
  ND2D1BWP30P140LVT U190 ( .A1(n275), .A2(i_data_bus[220]), .ZN(n154) );
  ND2D1BWP30P140LVT U191 ( .A1(n155), .A2(n154), .ZN(n156) );
  AOI21D1BWP30P140LVT U192 ( .A1(n1), .A2(i_data_bus[252]), .B(n156), .ZN(n158) );
  ND2D1BWP30P140LVT U193 ( .A1(n2), .A2(i_data_bus[28]), .ZN(n157) );
  ND4D1BWP30P140LVT U194 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U195 ( .A1(n168), .A2(i_data_bus[91]), .B1(n283), .B2(
        i_data_bus[59]), .ZN(n167) );
  AOI22D1BWP30P140LVT U196 ( .A1(n169), .A2(i_data_bus[123]), .B1(n285), .B2(
        i_data_bus[155]), .ZN(n166) );
  INVD1BWP30P140LVT U197 ( .I(i_data_bus[219]), .ZN(n162) );
  INVD1BWP30P140LVT U198 ( .I(i_data_bus[187]), .ZN(n161) );
  OAI22D1BWP30P140LVT U199 ( .A1(n290), .A2(n162), .B1(n248), .B2(n161), .ZN(
        n163) );
  AOI21D1BWP30P140LVT U200 ( .A1(n1), .A2(i_data_bus[251]), .B(n163), .ZN(n165) );
  ND2D1BWP30P140LVT U201 ( .A1(n2), .A2(i_data_bus[27]), .ZN(n164) );
  ND4D1BWP30P140LVT U202 ( .A1(n167), .A2(n166), .A3(n165), .A4(n164), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U203 ( .A1(n168), .A2(i_data_bus[90]), .B1(n283), .B2(
        i_data_bus[58]), .ZN(n176) );
  AOI22D1BWP30P140LVT U204 ( .A1(n169), .A2(i_data_bus[122]), .B1(n285), .B2(
        i_data_bus[154]), .ZN(n175) );
  INVD1BWP30P140LVT U205 ( .I(i_data_bus[218]), .ZN(n171) );
  INVD1BWP30P140LVT U206 ( .I(i_data_bus[186]), .ZN(n170) );
  OAI22D1BWP30P140LVT U207 ( .A1(n290), .A2(n171), .B1(n248), .B2(n170), .ZN(
        n172) );
  AOI21D1BWP30P140LVT U208 ( .A1(n1), .A2(i_data_bus[250]), .B(n172), .ZN(n174) );
  ND2D1BWP30P140LVT U209 ( .A1(n2), .A2(i_data_bus[26]), .ZN(n173) );
  ND4D1BWP30P140LVT U210 ( .A1(n176), .A2(n175), .A3(n174), .A4(n173), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U211 ( .A1(n274), .A2(i_data_bus[89]), .B1(n283), .B2(
        i_data_bus[57]), .ZN(n184) );
  INVD2BWP30P140LVT U212 ( .I(n177), .ZN(n286) );
  AOI22D1BWP30P140LVT U213 ( .A1(n286), .A2(i_data_bus[121]), .B1(n285), .B2(
        i_data_bus[153]), .ZN(n183) );
  INVD1BWP30P140LVT U214 ( .I(i_data_bus[217]), .ZN(n179) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[185]), .ZN(n178) );
  OAI22D1BWP30P140LVT U216 ( .A1(n207), .A2(n179), .B1(n288), .B2(n178), .ZN(
        n180) );
  AOI21D1BWP30P140LVT U217 ( .A1(n1), .A2(i_data_bus[249]), .B(n180), .ZN(n182) );
  ND2D1BWP30P140LVT U218 ( .A1(n2), .A2(i_data_bus[25]), .ZN(n181) );
  ND4D1BWP30P140LVT U219 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U220 ( .A1(n274), .A2(i_data_bus[88]), .B1(n283), .B2(
        i_data_bus[56]), .ZN(n191) );
  AOI22D1BWP30P140LVT U221 ( .A1(n286), .A2(i_data_bus[120]), .B1(n285), .B2(
        i_data_bus[152]), .ZN(n190) );
  INVD1BWP30P140LVT U222 ( .I(i_data_bus[216]), .ZN(n186) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[184]), .ZN(n185) );
  OAI22D1BWP30P140LVT U224 ( .A1(n207), .A2(n186), .B1(n248), .B2(n185), .ZN(
        n187) );
  AOI21D1BWP30P140LVT U225 ( .A1(n1), .A2(i_data_bus[248]), .B(n187), .ZN(n189) );
  ND2D1BWP30P140LVT U226 ( .A1(n2), .A2(i_data_bus[24]), .ZN(n188) );
  ND4D1BWP30P140LVT U227 ( .A1(n191), .A2(n190), .A3(n189), .A4(n188), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U228 ( .A1(n274), .A2(i_data_bus[87]), .B1(n283), .B2(
        i_data_bus[55]), .ZN(n198) );
  AOI22D1BWP30P140LVT U229 ( .A1(n286), .A2(i_data_bus[119]), .B1(n285), .B2(
        i_data_bus[151]), .ZN(n197) );
  INVD1BWP30P140LVT U230 ( .I(i_data_bus[215]), .ZN(n193) );
  INVD1BWP30P140LVT U231 ( .I(i_data_bus[183]), .ZN(n192) );
  OAI22D1BWP30P140LVT U232 ( .A1(n290), .A2(n193), .B1(n248), .B2(n192), .ZN(
        n194) );
  AOI21D1BWP30P140LVT U233 ( .A1(n1), .A2(i_data_bus[247]), .B(n194), .ZN(n196) );
  ND2D1BWP30P140LVT U234 ( .A1(n2), .A2(i_data_bus[23]), .ZN(n195) );
  ND4D1BWP30P140LVT U235 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U236 ( .A1(n274), .A2(i_data_bus[86]), .B1(n283), .B2(
        i_data_bus[54]), .ZN(n205) );
  AOI22D1BWP30P140LVT U237 ( .A1(n286), .A2(i_data_bus[118]), .B1(n285), .B2(
        i_data_bus[150]), .ZN(n204) );
  INVD1BWP30P140LVT U238 ( .I(i_data_bus[214]), .ZN(n200) );
  INVD1BWP30P140LVT U239 ( .I(i_data_bus[182]), .ZN(n199) );
  OAI22D1BWP30P140LVT U240 ( .A1(n207), .A2(n200), .B1(n248), .B2(n199), .ZN(
        n201) );
  AOI21D1BWP30P140LVT U241 ( .A1(n1), .A2(i_data_bus[246]), .B(n201), .ZN(n203) );
  ND2D1BWP30P140LVT U242 ( .A1(n2), .A2(i_data_bus[22]), .ZN(n202) );
  ND4D1BWP30P140LVT U243 ( .A1(n205), .A2(n204), .A3(n203), .A4(n202), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U244 ( .A1(n274), .A2(i_data_bus[85]), .B1(n283), .B2(
        i_data_bus[53]), .ZN(n215) );
  AOI22D1BWP30P140LVT U245 ( .A1(n286), .A2(i_data_bus[117]), .B1(n285), .B2(
        i_data_bus[149]), .ZN(n214) );
  INVD1BWP30P140LVT U246 ( .I(i_data_bus[245]), .ZN(n210) );
  INVD1BWP30P140LVT U247 ( .I(i_data_bus[181]), .ZN(n208) );
  INVD1BWP30P140LVT U248 ( .I(i_data_bus[213]), .ZN(n206) );
  OAI22D1BWP30P140LVT U249 ( .A1(n208), .A2(n248), .B1(n207), .B2(n206), .ZN(
        n209) );
  IAO21D1BWP30P140LVT U250 ( .A1(n211), .A2(n210), .B(n209), .ZN(n213) );
  ND2D1BWP30P140LVT U251 ( .A1(n2), .A2(i_data_bus[21]), .ZN(n212) );
  ND4D1BWP30P140LVT U252 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U253 ( .A1(n274), .A2(i_data_bus[84]), .B1(n283), .B2(
        i_data_bus[52]), .ZN(n222) );
  AOI22D1BWP30P140LVT U254 ( .A1(n286), .A2(i_data_bus[116]), .B1(n285), .B2(
        i_data_bus[148]), .ZN(n221) );
  INVD1BWP30P140LVT U255 ( .I(i_data_bus[212]), .ZN(n217) );
  INVD1BWP30P140LVT U256 ( .I(i_data_bus[180]), .ZN(n216) );
  OAI22D1BWP30P140LVT U257 ( .A1(n290), .A2(n217), .B1(n248), .B2(n216), .ZN(
        n218) );
  AOI21D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[244]), .B(n218), .ZN(n220) );
  ND2D1BWP30P140LVT U259 ( .A1(n2), .A2(i_data_bus[20]), .ZN(n219) );
  ND4D1BWP30P140LVT U260 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U261 ( .A1(n274), .A2(i_data_bus[83]), .B1(n283), .B2(
        i_data_bus[51]), .ZN(n228) );
  AOI22D1BWP30P140LVT U262 ( .A1(n286), .A2(i_data_bus[115]), .B1(n285), .B2(
        i_data_bus[147]), .ZN(n227) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[179]), .ZN(n223) );
  MOAI22D1BWP30P140LVT U264 ( .A1(n248), .A2(n223), .B1(n275), .B2(
        i_data_bus[211]), .ZN(n224) );
  AOI21D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[243]), .B(n224), .ZN(n226) );
  ND2D1BWP30P140LVT U266 ( .A1(n2), .A2(i_data_bus[19]), .ZN(n225) );
  ND4D1BWP30P140LVT U267 ( .A1(n228), .A2(n227), .A3(n226), .A4(n225), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U268 ( .A1(n274), .A2(i_data_bus[82]), .B1(n283), .B2(
        i_data_bus[50]), .ZN(n234) );
  AOI22D1BWP30P140LVT U269 ( .A1(n286), .A2(i_data_bus[114]), .B1(n285), .B2(
        i_data_bus[146]), .ZN(n233) );
  INVD1BWP30P140LVT U270 ( .I(i_data_bus[178]), .ZN(n229) );
  MOAI22D1BWP30P140LVT U271 ( .A1(n248), .A2(n229), .B1(n275), .B2(
        i_data_bus[210]), .ZN(n230) );
  AOI21D1BWP30P140LVT U272 ( .A1(n1), .A2(i_data_bus[242]), .B(n230), .ZN(n232) );
  ND2D1BWP30P140LVT U273 ( .A1(n2), .A2(i_data_bus[18]), .ZN(n231) );
  ND4D1BWP30P140LVT U274 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U275 ( .A1(n274), .A2(i_data_bus[81]), .B1(n283), .B2(
        i_data_bus[49]), .ZN(n240) );
  AOI22D1BWP30P140LVT U276 ( .A1(n286), .A2(i_data_bus[113]), .B1(n285), .B2(
        i_data_bus[145]), .ZN(n239) );
  INVD1BWP30P140LVT U277 ( .I(i_data_bus[177]), .ZN(n235) );
  MOAI22D1BWP30P140LVT U278 ( .A1(n248), .A2(n235), .B1(n275), .B2(
        i_data_bus[209]), .ZN(n236) );
  AOI21D1BWP30P140LVT U279 ( .A1(n1), .A2(i_data_bus[241]), .B(n236), .ZN(n238) );
  ND2D1BWP30P140LVT U280 ( .A1(n2), .A2(i_data_bus[17]), .ZN(n237) );
  ND4D1BWP30P140LVT U281 ( .A1(n240), .A2(n239), .A3(n238), .A4(n237), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U282 ( .A1(n274), .A2(i_data_bus[80]), .B1(n283), .B2(
        i_data_bus[48]), .ZN(n246) );
  AOI22D1BWP30P140LVT U283 ( .A1(n286), .A2(i_data_bus[112]), .B1(n285), .B2(
        i_data_bus[144]), .ZN(n245) );
  INVD1BWP30P140LVT U284 ( .I(i_data_bus[176]), .ZN(n241) );
  MOAI22D1BWP30P140LVT U285 ( .A1(n248), .A2(n241), .B1(n275), .B2(
        i_data_bus[208]), .ZN(n242) );
  AOI21D1BWP30P140LVT U286 ( .A1(n1), .A2(i_data_bus[240]), .B(n242), .ZN(n244) );
  ND2D1BWP30P140LVT U287 ( .A1(n2), .A2(i_data_bus[16]), .ZN(n243) );
  ND4D1BWP30P140LVT U288 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U289 ( .A1(n274), .A2(i_data_bus[79]), .B1(n283), .B2(
        i_data_bus[47]), .ZN(n253) );
  AOI22D1BWP30P140LVT U290 ( .A1(n286), .A2(i_data_bus[111]), .B1(n285), .B2(
        i_data_bus[143]), .ZN(n252) );
  INVD1BWP30P140LVT U291 ( .I(i_data_bus[175]), .ZN(n247) );
  MOAI22D1BWP30P140LVT U292 ( .A1(n248), .A2(n247), .B1(n275), .B2(
        i_data_bus[207]), .ZN(n249) );
  AOI21D1BWP30P140LVT U293 ( .A1(n1), .A2(i_data_bus[239]), .B(n249), .ZN(n251) );
  ND2D1BWP30P140LVT U294 ( .A1(n2), .A2(i_data_bus[15]), .ZN(n250) );
  ND4D1BWP30P140LVT U295 ( .A1(n253), .A2(n252), .A3(n251), .A4(n250), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U296 ( .A1(n274), .A2(i_data_bus[64]), .B1(n283), .B2(
        i_data_bus[32]), .ZN(n259) );
  AOI22D1BWP30P140LVT U297 ( .A1(n267), .A2(i_data_bus[96]), .B1(n266), .B2(
        i_data_bus[128]), .ZN(n258) );
  INR2D1BWP30P140LVT U298 ( .A1(i_data_bus[192]), .B1(n290), .ZN(n255) );
  INR2D1BWP30P140LVT U299 ( .A1(i_data_bus[160]), .B1(n277), .ZN(n254) );
  AOI211D1BWP30P140LVT U300 ( .A1(i_data_bus[224]), .A2(n1), .B(n255), .C(n254), .ZN(n257) );
  ND4D1BWP30P140LVT U301 ( .A1(n259), .A2(n258), .A3(n257), .A4(n256), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U302 ( .A1(n274), .A2(i_data_bus[66]), .B1(n283), .B2(
        i_data_bus[34]), .ZN(n265) );
  AOI22D1BWP30P140LVT U303 ( .A1(n267), .A2(i_data_bus[98]), .B1(n266), .B2(
        i_data_bus[130]), .ZN(n264) );
  INVD1BWP30P140LVT U304 ( .I(i_data_bus[162]), .ZN(n260) );
  MOAI22D1BWP30P140LVT U305 ( .A1(n277), .A2(n260), .B1(n275), .B2(
        i_data_bus[194]), .ZN(n261) );
  AOI21D1BWP30P140LVT U306 ( .A1(n1), .A2(i_data_bus[226]), .B(n261), .ZN(n263) );
  ND2D1BWP30P140LVT U307 ( .A1(n2), .A2(i_data_bus[2]), .ZN(n262) );
  ND4D1BWP30P140LVT U308 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U309 ( .A1(n274), .A2(i_data_bus[65]), .B1(n283), .B2(
        i_data_bus[33]), .ZN(n273) );
  AOI22D1BWP30P140LVT U310 ( .A1(n267), .A2(i_data_bus[97]), .B1(n266), .B2(
        i_data_bus[129]), .ZN(n272) );
  INVD1BWP30P140LVT U311 ( .I(i_data_bus[161]), .ZN(n268) );
  MOAI22D1BWP30P140LVT U312 ( .A1(n277), .A2(n268), .B1(n275), .B2(
        i_data_bus[193]), .ZN(n269) );
  AOI21D1BWP30P140LVT U313 ( .A1(n1), .A2(i_data_bus[225]), .B(n269), .ZN(n271) );
  ND2D1BWP30P140LVT U314 ( .A1(n2), .A2(i_data_bus[1]), .ZN(n270) );
  ND4D1BWP30P140LVT U315 ( .A1(n273), .A2(n272), .A3(n271), .A4(n270), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U316 ( .A1(n274), .A2(i_data_bus[78]), .B1(n283), .B2(
        i_data_bus[46]), .ZN(n282) );
  AOI22D1BWP30P140LVT U317 ( .A1(n286), .A2(i_data_bus[110]), .B1(n285), .B2(
        i_data_bus[142]), .ZN(n281) );
  INVD1BWP30P140LVT U318 ( .I(i_data_bus[174]), .ZN(n276) );
  MOAI22D1BWP30P140LVT U319 ( .A1(n277), .A2(n276), .B1(n275), .B2(
        i_data_bus[206]), .ZN(n278) );
  AOI21D1BWP30P140LVT U320 ( .A1(n1), .A2(i_data_bus[238]), .B(n278), .ZN(n280) );
  ND2D1BWP30P140LVT U321 ( .A1(n2), .A2(i_data_bus[14]), .ZN(n279) );
  ND4D1BWP30P140LVT U322 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U323 ( .A1(n284), .A2(i_data_bus[77]), .B1(n283), .B2(
        i_data_bus[45]), .ZN(n295) );
  AOI22D1BWP30P140LVT U324 ( .A1(n286), .A2(i_data_bus[109]), .B1(n285), .B2(
        i_data_bus[141]), .ZN(n294) );
  INVD1BWP30P140LVT U325 ( .I(i_data_bus[205]), .ZN(n289) );
  INVD1BWP30P140LVT U326 ( .I(i_data_bus[173]), .ZN(n287) );
  OAI22D1BWP30P140LVT U327 ( .A1(n290), .A2(n289), .B1(n288), .B2(n287), .ZN(
        n291) );
  AOI21D1BWP30P140LVT U328 ( .A1(n1), .A2(i_data_bus[237]), .B(n291), .ZN(n293) );
  ND2D1BWP30P140LVT U329 ( .A1(n2), .A2(i_data_bus[13]), .ZN(n292) );
  ND4D1BWP30P140LVT U330 ( .A1(n295), .A2(n294), .A3(n293), .A4(n292), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_10 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  OR2D1BWP30P140LVT U3 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n20) );
  INVD2BWP30P140LVT U4 ( .I(n22), .ZN(n279) );
  INVD2BWP30P140LVT U5 ( .I(n22), .ZN(n217) );
  INVD1BWP30P140LVT U6 ( .I(n22), .ZN(n159) );
  INVD2BWP30P140LVT U7 ( .I(n156), .ZN(n1) );
  INVD2BWP30P140LVT U8 ( .I(n157), .ZN(n2) );
  INVD4BWP30P140LVT U9 ( .I(n85), .ZN(n3) );
  INVD2BWP30P140LVT U10 ( .I(n267), .ZN(n281) );
  INVD1BWP30P140LVT U11 ( .I(n26), .ZN(n76) );
  INVD1BWP30P140LVT U12 ( .I(n34), .ZN(n158) );
  ND2D1BWP30P140LVT U13 ( .A1(n11), .A2(n10), .ZN(n13) );
  ND2D1BWP30P140LVT U14 ( .A1(n31), .A2(n6), .ZN(n37) );
  AOI21D1BWP30P140LVT U15 ( .A1(n283), .A2(i_data_bus[237]), .B(n282), .ZN(
        n286) );
  OR2D2BWP30P140LVT U16 ( .A1(n37), .A2(n36), .Z(n85) );
  INVD1BWP30P140LVT U17 ( .I(n8), .ZN(n163) );
  INR2D1BWP30P140LVT U18 ( .A1(n44), .B1(n43), .ZN(n157) );
  INVD1BWP30P140LVT U19 ( .I(i_cmd[0]), .ZN(n29) );
  INR3D0BWP30P140LVT U20 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n29), .ZN(n7)
         );
  INVD1BWP30P140LVT U21 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U22 ( .A1(n4), .A2(i_en), .ZN(n9) );
  NR2OPTPAD1BWP30P140LVT U23 ( .A1(i_cmd[5]), .A2(n9), .ZN(n5) );
  INR2D2BWP30P140LVT U24 ( .A1(n5), .B1(n20), .ZN(n31) );
  OR2D1BWP30P140LVT U25 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n42) );
  NR2D1BWP30P140LVT U26 ( .A1(n42), .A2(i_cmd[1]), .ZN(n6) );
  INR2D1BWP30P140LVT U27 ( .A1(n7), .B1(n37), .ZN(n8) );
  NR2D1BWP30P140LVT U28 ( .A1(i_cmd[3]), .A2(i_cmd[0]), .ZN(n11) );
  NR2D1BWP30P140LVT U29 ( .A1(i_cmd[4]), .A2(n9), .ZN(n10) );
  INVD1BWP30P140LVT U30 ( .I(i_cmd[2]), .ZN(n39) );
  INVD1BWP30P140LVT U31 ( .I(i_cmd[1]), .ZN(n12) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n39), .A2(n12), .ZN(n28) );
  OR2D2BWP30P140LVT U33 ( .A1(n13), .A2(n28), .Z(n24) );
  NR2D1BWP30P140LVT U34 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n15) );
  CKAN2D1BWP30P140LVT U35 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n14) );
  ND2D1BWP30P140LVT U36 ( .A1(n15), .A2(n14), .ZN(n16) );
  NR2OPTPAD1BWP30P140LVT U37 ( .A1(n24), .A2(n16), .ZN(n17) );
  INVD2BWP30P140LVT U38 ( .I(n17), .ZN(n18) );
  INVD3BWP30P140LVT U39 ( .I(n18), .ZN(n267) );
  ND2D1BWP30P140LVT U40 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n19) );
  NR2OPTPAD1BWP30P140LVT U41 ( .A1(n20), .A2(n19), .ZN(n21) );
  INR2D2BWP30P140LVT U42 ( .A1(n21), .B1(n24), .ZN(n22) );
  INVD1BWP30P140LVT U43 ( .I(i_cmd[7]), .ZN(n23) );
  INR4D0BWP30P140LVT U44 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n23), .ZN(n25) );
  INR2D1BWP30P140LVT U45 ( .A1(n25), .B1(n24), .ZN(n26) );
  INVD2BWP30P140LVT U46 ( .I(n76), .ZN(n283) );
  NR4D0BWP30P140LVT U47 ( .A1(n284), .A2(n267), .A3(n22), .A4(n283), .ZN(n46)
         );
  ND2D1BWP30P140LVT U48 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n27) );
  NR2D1BWP30P140LVT U49 ( .A1(n28), .A2(n27), .ZN(n33) );
  INVD1BWP30P140LVT U50 ( .I(i_cmd[4]), .ZN(n30) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n30), .A2(n29), .Z(n32) );
  ND2OPTIBD2BWP30P140LVT U52 ( .A1(n32), .A2(n31), .ZN(n43) );
  INR2D1BWP30P140LVT U53 ( .A1(n33), .B1(n43), .ZN(n34) );
  INVD1BWP30P140LVT U54 ( .I(n158), .ZN(n86) );
  ND2D1BWP30P140LVT U55 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n35) );
  OR2D1BWP30P140LVT U56 ( .A1(n35), .A2(i_cmd[0]), .Z(n36) );
  NR2D1BWP30P140LVT U57 ( .A1(n86), .A2(n3), .ZN(n45) );
  INVD1BWP30P140LVT U58 ( .I(i_valid[2]), .ZN(n38) );
  NR4D0BWP30P140LVT U59 ( .A1(n39), .A2(i_cmd[1]), .A3(i_cmd[3]), .A4(n38), 
        .ZN(n40) );
  INR2D2BWP30P140LVT U60 ( .A1(n40), .B1(n43), .ZN(n156) );
  ND2D1BWP30P140LVT U61 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n41) );
  NR2D1BWP30P140LVT U62 ( .A1(n42), .A2(n41), .ZN(n44) );
  ND4D1BWP30P140LVT U63 ( .A1(n46), .A2(n45), .A3(n1), .A4(n2), .ZN(N402) );
  INVD1BWP30P140LVT U64 ( .I(n2), .ZN(n84) );
  AOI22D1BWP30P140LVT U65 ( .A1(n276), .A2(i_data_bus[94]), .B1(n84), .B2(
        i_data_bus[62]), .ZN(n53) );
  AOI22D1BWP30P140LVT U66 ( .A1(n86), .A2(i_data_bus[126]), .B1(n3), .B2(
        i_data_bus[158]), .ZN(n52) );
  INVD1BWP30P140LVT U67 ( .I(n76), .ZN(n71) );
  INVD2BWP30P140LVT U68 ( .I(n267), .ZN(n250) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[222]), .ZN(n48) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[190]), .ZN(n47) );
  OAI22D1BWP30P140LVT U71 ( .A1(n250), .A2(n48), .B1(n159), .B2(n47), .ZN(n49)
         );
  AOI21D1BWP30P140LVT U72 ( .A1(n71), .A2(i_data_bus[254]), .B(n49), .ZN(n51)
         );
  ND2D1BWP30P140LVT U73 ( .A1(n262), .A2(i_data_bus[30]), .ZN(n50) );
  ND4D1BWP30P140LVT U74 ( .A1(n53), .A2(n52), .A3(n51), .A4(n50), .ZN(N399) );
  AOI22D1BWP30P140LVT U75 ( .A1(n258), .A2(i_data_bus[95]), .B1(n84), .B2(
        i_data_bus[63]), .ZN(n60) );
  AOI22D1BWP30P140LVT U76 ( .A1(n86), .A2(i_data_bus[127]), .B1(n3), .B2(
        i_data_bus[159]), .ZN(n59) );
  INVD1BWP30P140LVT U77 ( .I(i_data_bus[223]), .ZN(n55) );
  INVD1BWP30P140LVT U78 ( .I(i_data_bus[191]), .ZN(n54) );
  OAI22D1BWP30P140LVT U79 ( .A1(n250), .A2(n55), .B1(n159), .B2(n54), .ZN(n56)
         );
  AOI21D1BWP30P140LVT U80 ( .A1(n283), .A2(i_data_bus[255]), .B(n56), .ZN(n58)
         );
  ND2D1BWP30P140LVT U81 ( .A1(n284), .A2(i_data_bus[31]), .ZN(n57) );
  ND4D1BWP30P140LVT U82 ( .A1(n60), .A2(n59), .A3(n58), .A4(n57), .ZN(N400) );
  AOI22D1BWP30P140LVT U83 ( .A1(n156), .A2(i_data_bus[93]), .B1(n84), .B2(
        i_data_bus[61]), .ZN(n67) );
  AOI22D1BWP30P140LVT U84 ( .A1(n86), .A2(i_data_bus[125]), .B1(n3), .B2(
        i_data_bus[157]), .ZN(n66) );
  INVD1BWP30P140LVT U85 ( .I(i_data_bus[221]), .ZN(n62) );
  INVD1BWP30P140LVT U86 ( .I(i_data_bus[189]), .ZN(n61) );
  OAI22D1BWP30P140LVT U87 ( .A1(n250), .A2(n62), .B1(n217), .B2(n61), .ZN(n63)
         );
  AOI21D1BWP30P140LVT U88 ( .A1(n71), .A2(i_data_bus[253]), .B(n63), .ZN(n65)
         );
  ND2D1BWP30P140LVT U89 ( .A1(n262), .A2(i_data_bus[29]), .ZN(n64) );
  ND4D1BWP30P140LVT U90 ( .A1(n67), .A2(n66), .A3(n65), .A4(n64), .ZN(N398) );
  AOI22D1BWP30P140LVT U91 ( .A1(n156), .A2(i_data_bus[92]), .B1(n84), .B2(
        i_data_bus[60]), .ZN(n75) );
  AOI22D1BWP30P140LVT U92 ( .A1(n86), .A2(i_data_bus[124]), .B1(n3), .B2(
        i_data_bus[156]), .ZN(n74) );
  INVD1BWP30P140LVT U93 ( .I(i_data_bus[220]), .ZN(n69) );
  INVD1BWP30P140LVT U94 ( .I(i_data_bus[188]), .ZN(n68) );
  OAI22D1BWP30P140LVT U95 ( .A1(n250), .A2(n69), .B1(n217), .B2(n68), .ZN(n70)
         );
  AOI21D1BWP30P140LVT U96 ( .A1(n71), .A2(i_data_bus[252]), .B(n70), .ZN(n73)
         );
  ND2D1BWP30P140LVT U97 ( .A1(n284), .A2(i_data_bus[28]), .ZN(n72) );
  ND4D1BWP30P140LVT U98 ( .A1(n75), .A2(n74), .A3(n73), .A4(n72), .ZN(N397) );
  AOI22D1BWP30P140LVT U99 ( .A1(n156), .A2(i_data_bus[91]), .B1(n84), .B2(
        i_data_bus[59]), .ZN(n83) );
  AOI22D1BWP30P140LVT U100 ( .A1(n86), .A2(i_data_bus[123]), .B1(n3), .B2(
        i_data_bus[155]), .ZN(n82) );
  INVD2BWP30P140LVT U101 ( .I(n76), .ZN(n270) );
  INVD1BWP30P140LVT U102 ( .I(i_data_bus[219]), .ZN(n78) );
  INVD1BWP30P140LVT U103 ( .I(i_data_bus[187]), .ZN(n77) );
  OAI22D1BWP30P140LVT U104 ( .A1(n250), .A2(n78), .B1(n217), .B2(n77), .ZN(n79) );
  AOI21D1BWP30P140LVT U105 ( .A1(n270), .A2(i_data_bus[251]), .B(n79), .ZN(n81) );
  ND2D1BWP30P140LVT U106 ( .A1(n262), .A2(i_data_bus[27]), .ZN(n80) );
  ND4D1BWP30P140LVT U107 ( .A1(n83), .A2(n82), .A3(n81), .A4(n80), .ZN(N396)
         );
  AOI22D1BWP30P140LVT U108 ( .A1(n156), .A2(i_data_bus[90]), .B1(n84), .B2(
        i_data_bus[58]), .ZN(n93) );
  AOI22D1BWP30P140LVT U109 ( .A1(n86), .A2(i_data_bus[122]), .B1(n3), .B2(
        i_data_bus[154]), .ZN(n92) );
  INVD1BWP30P140LVT U110 ( .I(i_data_bus[218]), .ZN(n88) );
  INVD1BWP30P140LVT U111 ( .I(i_data_bus[186]), .ZN(n87) );
  OAI22D1BWP30P140LVT U112 ( .A1(n250), .A2(n88), .B1(n217), .B2(n87), .ZN(n89) );
  AOI21D1BWP30P140LVT U113 ( .A1(n270), .A2(i_data_bus[250]), .B(n89), .ZN(n91) );
  ND2D1BWP30P140LVT U114 ( .A1(n8), .A2(i_data_bus[26]), .ZN(n90) );
  ND4D1BWP30P140LVT U115 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(N395)
         );
  INVD2BWP30P140LVT U116 ( .I(n1), .ZN(n276) );
  INVD2BWP30P140LVT U117 ( .I(n2), .ZN(n275) );
  AOI22D1BWP30P140LVT U118 ( .A1(n276), .A2(i_data_bus[89]), .B1(n275), .B2(
        i_data_bus[57]), .ZN(n100) );
  INVD2BWP30P140LVT U119 ( .I(n158), .ZN(n277) );
  AOI22D1BWP30P140LVT U120 ( .A1(n277), .A2(i_data_bus[121]), .B1(n3), .B2(
        i_data_bus[153]), .ZN(n99) );
  INVD1BWP30P140LVT U121 ( .I(i_data_bus[217]), .ZN(n95) );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[185]), .ZN(n94) );
  OAI22D1BWP30P140LVT U123 ( .A1(n250), .A2(n95), .B1(n217), .B2(n94), .ZN(n96) );
  AOI21D1BWP30P140LVT U124 ( .A1(n270), .A2(i_data_bus[249]), .B(n96), .ZN(n98) );
  INVD2BWP30P140LVT U125 ( .I(n163), .ZN(n284) );
  ND2D1BWP30P140LVT U126 ( .A1(n284), .A2(i_data_bus[25]), .ZN(n97) );
  ND4D1BWP30P140LVT U127 ( .A1(n100), .A2(n99), .A3(n98), .A4(n97), .ZN(N394)
         );
  AOI22D1BWP30P140LVT U128 ( .A1(n276), .A2(i_data_bus[88]), .B1(n275), .B2(
        i_data_bus[56]), .ZN(n107) );
  AOI22D1BWP30P140LVT U129 ( .A1(n277), .A2(i_data_bus[120]), .B1(n3), .B2(
        i_data_bus[152]), .ZN(n106) );
  INVD1BWP30P140LVT U130 ( .I(i_data_bus[216]), .ZN(n102) );
  INVD1BWP30P140LVT U131 ( .I(i_data_bus[184]), .ZN(n101) );
  OAI22D1BWP30P140LVT U132 ( .A1(n281), .A2(n102), .B1(n217), .B2(n101), .ZN(
        n103) );
  AOI21D1BWP30P140LVT U133 ( .A1(n270), .A2(i_data_bus[248]), .B(n103), .ZN(
        n105) );
  ND2D1BWP30P140LVT U134 ( .A1(n284), .A2(i_data_bus[24]), .ZN(n104) );
  ND4D1BWP30P140LVT U135 ( .A1(n107), .A2(n106), .A3(n105), .A4(n104), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U136 ( .A1(n276), .A2(i_data_bus[87]), .B1(n275), .B2(
        i_data_bus[55]), .ZN(n114) );
  AOI22D1BWP30P140LVT U137 ( .A1(n277), .A2(i_data_bus[119]), .B1(n3), .B2(
        i_data_bus[151]), .ZN(n113) );
  INVD1BWP30P140LVT U138 ( .I(i_data_bus[215]), .ZN(n109) );
  INVD1BWP30P140LVT U139 ( .I(i_data_bus[183]), .ZN(n108) );
  OAI22D1BWP30P140LVT U140 ( .A1(n281), .A2(n109), .B1(n217), .B2(n108), .ZN(
        n110) );
  AOI21D1BWP30P140LVT U141 ( .A1(n270), .A2(i_data_bus[247]), .B(n110), .ZN(
        n112) );
  ND2D1BWP30P140LVT U142 ( .A1(n284), .A2(i_data_bus[23]), .ZN(n111) );
  ND4D1BWP30P140LVT U143 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U144 ( .A1(n276), .A2(i_data_bus[86]), .B1(n275), .B2(
        i_data_bus[54]), .ZN(n121) );
  AOI22D1BWP30P140LVT U145 ( .A1(n277), .A2(i_data_bus[118]), .B1(n3), .B2(
        i_data_bus[150]), .ZN(n120) );
  INVD1BWP30P140LVT U146 ( .I(i_data_bus[214]), .ZN(n116) );
  INVD1BWP30P140LVT U147 ( .I(i_data_bus[182]), .ZN(n115) );
  OAI22D1BWP30P140LVT U148 ( .A1(n281), .A2(n116), .B1(n217), .B2(n115), .ZN(
        n117) );
  AOI21D1BWP30P140LVT U149 ( .A1(n270), .A2(i_data_bus[246]), .B(n117), .ZN(
        n119) );
  ND2D1BWP30P140LVT U150 ( .A1(n284), .A2(i_data_bus[22]), .ZN(n118) );
  ND4D1BWP30P140LVT U151 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U152 ( .A1(n276), .A2(i_data_bus[85]), .B1(n275), .B2(
        i_data_bus[53]), .ZN(n128) );
  AOI22D1BWP30P140LVT U153 ( .A1(n277), .A2(i_data_bus[117]), .B1(n3), .B2(
        i_data_bus[149]), .ZN(n127) );
  INVD1BWP30P140LVT U154 ( .I(i_data_bus[213]), .ZN(n123) );
  INVD1BWP30P140LVT U155 ( .I(i_data_bus[181]), .ZN(n122) );
  OAI22D1BWP30P140LVT U156 ( .A1(n281), .A2(n123), .B1(n217), .B2(n122), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U157 ( .A1(n270), .A2(i_data_bus[245]), .B(n124), .ZN(
        n126) );
  ND2D1BWP30P140LVT U158 ( .A1(n284), .A2(i_data_bus[21]), .ZN(n125) );
  ND4D1BWP30P140LVT U159 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U160 ( .A1(n276), .A2(i_data_bus[84]), .B1(n275), .B2(
        i_data_bus[52]), .ZN(n135) );
  AOI22D1BWP30P140LVT U161 ( .A1(n277), .A2(i_data_bus[116]), .B1(n3), .B2(
        i_data_bus[148]), .ZN(n134) );
  INVD1BWP30P140LVT U162 ( .I(i_data_bus[212]), .ZN(n130) );
  INVD1BWP30P140LVT U163 ( .I(i_data_bus[180]), .ZN(n129) );
  OAI22D1BWP30P140LVT U164 ( .A1(n281), .A2(n130), .B1(n217), .B2(n129), .ZN(
        n131) );
  AOI21D1BWP30P140LVT U165 ( .A1(n270), .A2(i_data_bus[244]), .B(n131), .ZN(
        n133) );
  ND2D1BWP30P140LVT U166 ( .A1(n284), .A2(i_data_bus[20]), .ZN(n132) );
  ND4D1BWP30P140LVT U167 ( .A1(n135), .A2(n134), .A3(n133), .A4(n132), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U168 ( .A1(n276), .A2(i_data_bus[83]), .B1(n275), .B2(
        i_data_bus[51]), .ZN(n142) );
  AOI22D1BWP30P140LVT U169 ( .A1(n277), .A2(i_data_bus[115]), .B1(n3), .B2(
        i_data_bus[147]), .ZN(n141) );
  INVD1BWP30P140LVT U170 ( .I(i_data_bus[211]), .ZN(n137) );
  INVD1BWP30P140LVT U171 ( .I(i_data_bus[179]), .ZN(n136) );
  OAI22D1BWP30P140LVT U172 ( .A1(n281), .A2(n137), .B1(n217), .B2(n136), .ZN(
        n138) );
  AOI21D1BWP30P140LVT U173 ( .A1(n270), .A2(i_data_bus[243]), .B(n138), .ZN(
        n140) );
  ND2D1BWP30P140LVT U174 ( .A1(n284), .A2(i_data_bus[19]), .ZN(n139) );
  ND4D1BWP30P140LVT U175 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U176 ( .A1(n276), .A2(i_data_bus[82]), .B1(n275), .B2(
        i_data_bus[50]), .ZN(n149) );
  AOI22D1BWP30P140LVT U177 ( .A1(n277), .A2(i_data_bus[114]), .B1(n3), .B2(
        i_data_bus[146]), .ZN(n148) );
  INVD1BWP30P140LVT U178 ( .I(i_data_bus[210]), .ZN(n144) );
  INVD1BWP30P140LVT U179 ( .I(i_data_bus[178]), .ZN(n143) );
  OAI22D1BWP30P140LVT U180 ( .A1(n281), .A2(n144), .B1(n217), .B2(n143), .ZN(
        n145) );
  AOI21D1BWP30P140LVT U181 ( .A1(n270), .A2(i_data_bus[242]), .B(n145), .ZN(
        n147) );
  ND2D1BWP30P140LVT U182 ( .A1(n284), .A2(i_data_bus[18]), .ZN(n146) );
  ND4D1BWP30P140LVT U183 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U184 ( .A1(n276), .A2(i_data_bus[81]), .B1(n275), .B2(
        i_data_bus[49]), .ZN(n155) );
  AOI22D1BWP30P140LVT U185 ( .A1(n277), .A2(i_data_bus[113]), .B1(n3), .B2(
        i_data_bus[145]), .ZN(n154) );
  INVD1BWP30P140LVT U186 ( .I(i_data_bus[177]), .ZN(n150) );
  MOAI22D1BWP30P140LVT U187 ( .A1(n217), .A2(n150), .B1(n267), .B2(
        i_data_bus[209]), .ZN(n151) );
  AOI21D1BWP30P140LVT U188 ( .A1(n270), .A2(i_data_bus[241]), .B(n151), .ZN(
        n153) );
  ND2D1BWP30P140LVT U189 ( .A1(n284), .A2(i_data_bus[17]), .ZN(n152) );
  ND4D1BWP30P140LVT U190 ( .A1(n155), .A2(n154), .A3(n153), .A4(n152), .ZN(
        N386) );
  INVD2BWP30P140LVT U191 ( .I(n1), .ZN(n258) );
  INVD2BWP30P140LVT U192 ( .I(n2), .ZN(n257) );
  AOI22D1BWP30P140LVT U193 ( .A1(n258), .A2(i_data_bus[76]), .B1(n257), .B2(
        i_data_bus[44]), .ZN(n167) );
  INVD2BWP30P140LVT U194 ( .I(n158), .ZN(n259) );
  AOI22D1BWP30P140LVT U195 ( .A1(n259), .A2(i_data_bus[108]), .B1(n3), .B2(
        i_data_bus[140]), .ZN(n166) );
  INVD1BWP30P140LVT U196 ( .I(i_data_bus[204]), .ZN(n161) );
  INVD1BWP30P140LVT U197 ( .I(i_data_bus[172]), .ZN(n160) );
  OAI22D1BWP30P140LVT U198 ( .A1(n281), .A2(n161), .B1(n279), .B2(n160), .ZN(
        n162) );
  AOI21D1BWP30P140LVT U199 ( .A1(n283), .A2(i_data_bus[236]), .B(n162), .ZN(
        n165) );
  INVD2BWP30P140LVT U200 ( .I(n163), .ZN(n262) );
  ND2D1BWP30P140LVT U201 ( .A1(n262), .A2(i_data_bus[12]), .ZN(n164) );
  ND4D1BWP30P140LVT U202 ( .A1(n167), .A2(n166), .A3(n165), .A4(n164), .ZN(
        N381) );
  AOI22D1BWP30P140LVT U203 ( .A1(n258), .A2(i_data_bus[75]), .B1(n257), .B2(
        i_data_bus[43]), .ZN(n174) );
  AOI22D1BWP30P140LVT U204 ( .A1(n259), .A2(i_data_bus[107]), .B1(n3), .B2(
        i_data_bus[139]), .ZN(n173) );
  INVD1BWP30P140LVT U205 ( .I(i_data_bus[203]), .ZN(n169) );
  INVD1BWP30P140LVT U206 ( .I(i_data_bus[171]), .ZN(n168) );
  OAI22D1BWP30P140LVT U207 ( .A1(n281), .A2(n169), .B1(n279), .B2(n168), .ZN(
        n170) );
  AOI21D1BWP30P140LVT U208 ( .A1(n283), .A2(i_data_bus[235]), .B(n170), .ZN(
        n172) );
  ND2D1BWP30P140LVT U209 ( .A1(n262), .A2(i_data_bus[11]), .ZN(n171) );
  ND4D1BWP30P140LVT U210 ( .A1(n174), .A2(n173), .A3(n172), .A4(n171), .ZN(
        N380) );
  AOI22D1BWP30P140LVT U211 ( .A1(n258), .A2(i_data_bus[74]), .B1(n257), .B2(
        i_data_bus[42]), .ZN(n181) );
  AOI22D1BWP30P140LVT U212 ( .A1(n259), .A2(i_data_bus[106]), .B1(n3), .B2(
        i_data_bus[138]), .ZN(n180) );
  INVD1BWP30P140LVT U213 ( .I(i_data_bus[202]), .ZN(n176) );
  INVD1BWP30P140LVT U214 ( .I(i_data_bus[170]), .ZN(n175) );
  OAI22D1BWP30P140LVT U215 ( .A1(n281), .A2(n176), .B1(n279), .B2(n175), .ZN(
        n177) );
  AOI21D1BWP30P140LVT U216 ( .A1(n283), .A2(i_data_bus[234]), .B(n177), .ZN(
        n179) );
  ND2D1BWP30P140LVT U217 ( .A1(n262), .A2(i_data_bus[10]), .ZN(n178) );
  ND4D1BWP30P140LVT U218 ( .A1(n181), .A2(n180), .A3(n179), .A4(n178), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U219 ( .A1(n258), .A2(i_data_bus[73]), .B1(n257), .B2(
        i_data_bus[41]), .ZN(n188) );
  AOI22D1BWP30P140LVT U220 ( .A1(n259), .A2(i_data_bus[105]), .B1(n3), .B2(
        i_data_bus[137]), .ZN(n187) );
  INVD1BWP30P140LVT U221 ( .I(i_data_bus[201]), .ZN(n183) );
  INVD1BWP30P140LVT U222 ( .I(i_data_bus[169]), .ZN(n182) );
  OAI22D1BWP30P140LVT U223 ( .A1(n281), .A2(n183), .B1(n279), .B2(n182), .ZN(
        n184) );
  AOI21D1BWP30P140LVT U224 ( .A1(n283), .A2(i_data_bus[233]), .B(n184), .ZN(
        n186) );
  ND2D1BWP30P140LVT U225 ( .A1(n262), .A2(i_data_bus[9]), .ZN(n185) );
  ND4D1BWP30P140LVT U226 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U227 ( .A1(n258), .A2(i_data_bus[71]), .B1(n257), .B2(
        i_data_bus[39]), .ZN(n195) );
  AOI22D1BWP30P140LVT U228 ( .A1(n259), .A2(i_data_bus[103]), .B1(n3), .B2(
        i_data_bus[135]), .ZN(n194) );
  INVD1BWP30P140LVT U229 ( .I(i_data_bus[199]), .ZN(n190) );
  INVD1BWP30P140LVT U230 ( .I(i_data_bus[167]), .ZN(n189) );
  OAI22D1BWP30P140LVT U231 ( .A1(n281), .A2(n190), .B1(n279), .B2(n189), .ZN(
        n191) );
  AOI21D1BWP30P140LVT U232 ( .A1(n283), .A2(i_data_bus[231]), .B(n191), .ZN(
        n193) );
  ND2D1BWP30P140LVT U233 ( .A1(n262), .A2(i_data_bus[7]), .ZN(n192) );
  ND4D1BWP30P140LVT U234 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U235 ( .A1(n258), .A2(i_data_bus[70]), .B1(n257), .B2(
        i_data_bus[38]), .ZN(n202) );
  AOI22D1BWP30P140LVT U236 ( .A1(n259), .A2(i_data_bus[102]), .B1(n3), .B2(
        i_data_bus[134]), .ZN(n201) );
  INVD1BWP30P140LVT U237 ( .I(i_data_bus[198]), .ZN(n197) );
  INVD1BWP30P140LVT U238 ( .I(i_data_bus[166]), .ZN(n196) );
  OAI22D1BWP30P140LVT U239 ( .A1(n281), .A2(n197), .B1(n279), .B2(n196), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U240 ( .A1(n283), .A2(i_data_bus[230]), .B(n198), .ZN(
        n200) );
  ND2D1BWP30P140LVT U241 ( .A1(n262), .A2(i_data_bus[6]), .ZN(n199) );
  ND4D1BWP30P140LVT U242 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U243 ( .A1(n258), .A2(i_data_bus[69]), .B1(n257), .B2(
        i_data_bus[37]), .ZN(n209) );
  AOI22D1BWP30P140LVT U244 ( .A1(n259), .A2(i_data_bus[101]), .B1(n3), .B2(
        i_data_bus[133]), .ZN(n208) );
  INVD1BWP30P140LVT U245 ( .I(i_data_bus[197]), .ZN(n204) );
  INVD1BWP30P140LVT U246 ( .I(i_data_bus[165]), .ZN(n203) );
  OAI22D1BWP30P140LVT U247 ( .A1(n281), .A2(n204), .B1(n279), .B2(n203), .ZN(
        n205) );
  AOI21D1BWP30P140LVT U248 ( .A1(n283), .A2(i_data_bus[229]), .B(n205), .ZN(
        n207) );
  ND2D1BWP30P140LVT U249 ( .A1(n262), .A2(i_data_bus[5]), .ZN(n206) );
  ND4D1BWP30P140LVT U250 ( .A1(n209), .A2(n208), .A3(n207), .A4(n206), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U251 ( .A1(n276), .A2(i_data_bus[80]), .B1(n275), .B2(
        i_data_bus[48]), .ZN(n215) );
  AOI22D1BWP30P140LVT U252 ( .A1(n277), .A2(i_data_bus[112]), .B1(n3), .B2(
        i_data_bus[144]), .ZN(n214) );
  INVD1BWP30P140LVT U253 ( .I(i_data_bus[176]), .ZN(n210) );
  MOAI22D1BWP30P140LVT U254 ( .A1(n217), .A2(n210), .B1(n267), .B2(
        i_data_bus[208]), .ZN(n211) );
  AOI21D1BWP30P140LVT U255 ( .A1(n270), .A2(i_data_bus[240]), .B(n211), .ZN(
        n213) );
  ND2D1BWP30P140LVT U256 ( .A1(n284), .A2(i_data_bus[16]), .ZN(n212) );
  ND4D1BWP30P140LVT U257 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U258 ( .A1(n276), .A2(i_data_bus[79]), .B1(n275), .B2(
        i_data_bus[47]), .ZN(n222) );
  AOI22D1BWP30P140LVT U259 ( .A1(n277), .A2(i_data_bus[111]), .B1(n3), .B2(
        i_data_bus[143]), .ZN(n221) );
  INVD1BWP30P140LVT U260 ( .I(i_data_bus[175]), .ZN(n216) );
  MOAI22D1BWP30P140LVT U261 ( .A1(n217), .A2(n216), .B1(n267), .B2(
        i_data_bus[207]), .ZN(n218) );
  AOI21D1BWP30P140LVT U262 ( .A1(n270), .A2(i_data_bus[239]), .B(n218), .ZN(
        n220) );
  ND2D1BWP30P140LVT U263 ( .A1(n284), .A2(i_data_bus[15]), .ZN(n219) );
  ND4D1BWP30P140LVT U264 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U265 ( .A1(n258), .A2(i_data_bus[68]), .B1(n257), .B2(
        i_data_bus[36]), .ZN(n229) );
  AOI22D1BWP30P140LVT U266 ( .A1(n259), .A2(i_data_bus[100]), .B1(n3), .B2(
        i_data_bus[132]), .ZN(n228) );
  INVD1BWP30P140LVT U267 ( .I(i_data_bus[196]), .ZN(n224) );
  INVD1BWP30P140LVT U268 ( .I(i_data_bus[164]), .ZN(n223) );
  OAI22D1BWP30P140LVT U269 ( .A1(n281), .A2(n224), .B1(n279), .B2(n223), .ZN(
        n225) );
  AOI21D1BWP30P140LVT U270 ( .A1(n283), .A2(i_data_bus[228]), .B(n225), .ZN(
        n227) );
  ND2D1BWP30P140LVT U271 ( .A1(n262), .A2(i_data_bus[4]), .ZN(n226) );
  ND4D1BWP30P140LVT U272 ( .A1(n229), .A2(n228), .A3(n227), .A4(n226), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U273 ( .A1(n258), .A2(i_data_bus[67]), .B1(n257), .B2(
        i_data_bus[35]), .ZN(n236) );
  AOI22D1BWP30P140LVT U274 ( .A1(n259), .A2(i_data_bus[99]), .B1(n3), .B2(
        i_data_bus[131]), .ZN(n235) );
  INVD1BWP30P140LVT U275 ( .I(i_data_bus[195]), .ZN(n231) );
  INVD1BWP30P140LVT U276 ( .I(i_data_bus[163]), .ZN(n230) );
  OAI22D1BWP30P140LVT U277 ( .A1(n281), .A2(n231), .B1(n279), .B2(n230), .ZN(
        n232) );
  AOI21D1BWP30P140LVT U278 ( .A1(n283), .A2(i_data_bus[227]), .B(n232), .ZN(
        n234) );
  ND2D1BWP30P140LVT U279 ( .A1(n262), .A2(i_data_bus[3]), .ZN(n233) );
  ND4D1BWP30P140LVT U280 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U281 ( .A1(n258), .A2(i_data_bus[66]), .B1(n257), .B2(
        i_data_bus[34]), .ZN(n242) );
  AOI22D1BWP30P140LVT U282 ( .A1(n259), .A2(i_data_bus[98]), .B1(n3), .B2(
        i_data_bus[130]), .ZN(n241) );
  INVD1BWP30P140LVT U283 ( .I(i_data_bus[162]), .ZN(n237) );
  MOAI22D1BWP30P140LVT U284 ( .A1(n279), .A2(n237), .B1(n267), .B2(
        i_data_bus[194]), .ZN(n238) );
  AOI21D1BWP30P140LVT U285 ( .A1(n283), .A2(i_data_bus[226]), .B(n238), .ZN(
        n240) );
  ND2D1BWP30P140LVT U286 ( .A1(n262), .A2(i_data_bus[2]), .ZN(n239) );
  ND4D1BWP30P140LVT U287 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U288 ( .A1(n258), .A2(i_data_bus[65]), .B1(n257), .B2(
        i_data_bus[33]), .ZN(n248) );
  AOI22D1BWP30P140LVT U289 ( .A1(n259), .A2(i_data_bus[97]), .B1(n3), .B2(
        i_data_bus[129]), .ZN(n247) );
  INVD1BWP30P140LVT U290 ( .I(i_data_bus[161]), .ZN(n243) );
  MOAI22D1BWP30P140LVT U291 ( .A1(n279), .A2(n243), .B1(n267), .B2(
        i_data_bus[193]), .ZN(n244) );
  AOI21D1BWP30P140LVT U292 ( .A1(n283), .A2(i_data_bus[225]), .B(n244), .ZN(
        n246) );
  ND2D1BWP30P140LVT U293 ( .A1(n262), .A2(i_data_bus[1]), .ZN(n245) );
  ND4D1BWP30P140LVT U294 ( .A1(n248), .A2(n247), .A3(n246), .A4(n245), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U295 ( .A1(n258), .A2(i_data_bus[72]), .B1(n257), .B2(
        i_data_bus[40]), .ZN(n256) );
  AOI22D1BWP30P140LVT U296 ( .A1(n259), .A2(i_data_bus[104]), .B1(n3), .B2(
        i_data_bus[136]), .ZN(n255) );
  INVD1BWP30P140LVT U297 ( .I(i_data_bus[168]), .ZN(n251) );
  INVD1BWP30P140LVT U298 ( .I(i_data_bus[200]), .ZN(n249) );
  OAI22D1BWP30P140LVT U299 ( .A1(n279), .A2(n251), .B1(n250), .B2(n249), .ZN(
        n252) );
  AOI21D1BWP30P140LVT U300 ( .A1(n270), .A2(i_data_bus[232]), .B(n252), .ZN(
        n254) );
  ND2D1BWP30P140LVT U301 ( .A1(n262), .A2(i_data_bus[8]), .ZN(n253) );
  ND4D1BWP30P140LVT U302 ( .A1(n256), .A2(n255), .A3(n254), .A4(n253), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U303 ( .A1(n258), .A2(i_data_bus[64]), .B1(n257), .B2(
        i_data_bus[32]), .ZN(n266) );
  AOI22D1BWP30P140LVT U304 ( .A1(n259), .A2(i_data_bus[96]), .B1(n3), .B2(
        i_data_bus[128]), .ZN(n265) );
  INR2D1BWP30P140LVT U305 ( .A1(i_data_bus[192]), .B1(n281), .ZN(n261) );
  INR2D1BWP30P140LVT U306 ( .A1(i_data_bus[160]), .B1(n279), .ZN(n260) );
  AOI211D1BWP30P140LVT U307 ( .A1(i_data_bus[224]), .A2(n283), .B(n261), .C(
        n260), .ZN(n264) );
  ND2D1BWP30P140LVT U308 ( .A1(n262), .A2(i_data_bus[0]), .ZN(n263) );
  ND4D1BWP30P140LVT U309 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U310 ( .A1(n276), .A2(i_data_bus[78]), .B1(n275), .B2(
        i_data_bus[46]), .ZN(n274) );
  AOI22D1BWP30P140LVT U311 ( .A1(n277), .A2(i_data_bus[110]), .B1(n3), .B2(
        i_data_bus[142]), .ZN(n273) );
  INVD1BWP30P140LVT U312 ( .I(i_data_bus[174]), .ZN(n268) );
  MOAI22D1BWP30P140LVT U313 ( .A1(n279), .A2(n268), .B1(n267), .B2(
        i_data_bus[206]), .ZN(n269) );
  AOI21D1BWP30P140LVT U314 ( .A1(n270), .A2(i_data_bus[238]), .B(n269), .ZN(
        n272) );
  ND2D1BWP30P140LVT U315 ( .A1(n284), .A2(i_data_bus[14]), .ZN(n271) );
  ND4D1BWP30P140LVT U316 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U317 ( .A1(n276), .A2(i_data_bus[77]), .B1(n275), .B2(
        i_data_bus[45]), .ZN(n288) );
  AOI22D1BWP30P140LVT U318 ( .A1(n277), .A2(i_data_bus[109]), .B1(n3), .B2(
        i_data_bus[141]), .ZN(n287) );
  INVD1BWP30P140LVT U319 ( .I(i_data_bus[205]), .ZN(n280) );
  INVD1BWP30P140LVT U320 ( .I(i_data_bus[173]), .ZN(n278) );
  OAI22D1BWP30P140LVT U321 ( .A1(n281), .A2(n280), .B1(n279), .B2(n278), .ZN(
        n282) );
  ND2D1BWP30P140LVT U322 ( .A1(n284), .A2(i_data_bus[13]), .ZN(n285) );
  ND4D1BWP30P140LVT U323 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_11 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n47), .ZN(n2) );
  ND2OPTIBD1BWP30P140LVT U4 ( .A1(n36), .A2(n5), .ZN(n47) );
  INVD4BWP30P140LVT U5 ( .I(n145), .ZN(n1) );
  INVD3BWP30P140LVT U6 ( .I(n183), .ZN(n3) );
  INR2D1BWP30P140LVT U7 ( .A1(n35), .B1(n32), .ZN(n10) );
  NR2OPTPAD1BWP30P140LVT U8 ( .A1(n16), .A2(n15), .ZN(n20) );
  AOI21D1BWP30P140LVT U9 ( .A1(n268), .A2(i_data_bus[239]), .B(n195), .ZN(n197) );
  IND3D2BWP30P140LVT U10 ( .A1(n14), .B1(n13), .B2(n21), .ZN(n48) );
  NR2D3BWP30P140LVT U11 ( .A1(n15), .A2(n18), .ZN(n21) );
  INVD1BWP30P140LVT U12 ( .I(n4), .ZN(n274) );
  INVD1BWP30P140LVT U13 ( .I(n4), .ZN(n281) );
  ND2D1BWP30P140LVT U14 ( .A1(n27), .A2(n7), .ZN(n32) );
  ND2D1BWP30P140LVT U15 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n17) );
  INVD1BWP30P140LVT U16 ( .I(n129), .ZN(n244) );
  INVD1BWP30P140LVT U17 ( .I(n48), .ZN(n129) );
  ND2D1BWP30P140LVT U18 ( .A1(n287), .A2(i_data_bus[1]), .ZN(n111) );
  ND2D1BWP30P140LVT U19 ( .A1(n287), .A2(i_data_bus[2]), .ZN(n97) );
  ND2D1BWP30P140LVT U20 ( .A1(n287), .A2(i_data_bus[3]), .ZN(n125) );
  ND2D1BWP30P140LVT U21 ( .A1(n287), .A2(i_data_bus[4]), .ZN(n118) );
  ND2D1BWP30P140LVT U22 ( .A1(n287), .A2(i_data_bus[5]), .ZN(n76) );
  ND2D1BWP30P140LVT U23 ( .A1(n287), .A2(i_data_bus[6]), .ZN(n62) );
  ND2D1BWP30P140LVT U24 ( .A1(n287), .A2(i_data_bus[7]), .ZN(n104) );
  AOI21D1BWP30P140LVT U25 ( .A1(n268), .A2(i_data_bus[232]), .B(n169), .ZN(
        n171) );
  ND2D1BWP30P140LVT U26 ( .A1(n287), .A2(i_data_bus[8]), .ZN(n170) );
  ND2D1BWP30P140LVT U27 ( .A1(n287), .A2(i_data_bus[9]), .ZN(n69) );
  ND2D1BWP30P140LVT U28 ( .A1(n287), .A2(i_data_bus[10]), .ZN(n83) );
  ND2D1BWP30P140LVT U29 ( .A1(n287), .A2(i_data_bus[11]), .ZN(n90) );
  ND2D1BWP30P140LVT U30 ( .A1(n287), .A2(i_data_bus[12]), .ZN(n55) );
  AOI21D1BWP30P140LVT U31 ( .A1(n268), .A2(i_data_bus[238]), .B(n267), .ZN(
        n270) );
  INR2D1BWP30P140LVT U32 ( .A1(n43), .B1(n40), .ZN(n184) );
  INVD1BWP30P140LVT U33 ( .I(n184), .ZN(n46) );
  ND2OPTIBD1BWP30P140LVT U34 ( .A1(n21), .A2(n24), .ZN(n137) );
  OR2D1BWP30P140LVT U35 ( .A1(n40), .A2(n31), .Z(n4) );
  OR2D1BWP30P140LVT U36 ( .A1(n40), .A2(n39), .Z(n183) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n35), .A2(n34), .Z(n5) );
  OR2D1BWP30P140LVT U38 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n42) );
  NR2D1BWP30P140LVT U39 ( .A1(n42), .A2(i_cmd[1]), .ZN(n35) );
  OR2D2BWP30P140LVT U40 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n16) );
  NR2OPTPAD1BWP30P140LVT U41 ( .A1(i_cmd[5]), .A2(n16), .ZN(n27) );
  INVD1BWP30P140LVT U42 ( .I(rst), .ZN(n6) );
  ND2D1BWP30P140LVT U43 ( .A1(n6), .A2(i_en), .ZN(n11) );
  INVD1BWP30P140LVT U44 ( .I(n11), .ZN(n7) );
  INVD1BWP30P140LVT U45 ( .I(i_cmd[0]), .ZN(n8) );
  INR3D0BWP30P140LVT U46 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n8), .ZN(n9) );
  ND2OPTIBD2BWP30P140LVT U47 ( .A1(n10), .A2(n9), .ZN(n188) );
  ND2D1BWP30P140LVT U48 ( .A1(i_cmd[6]), .A2(i_valid[6]), .ZN(n14) );
  NR2D1BWP30P140LVT U49 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n13) );
  OR2D4BWP30P140LVT U50 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .Z(n30) );
  OR2D4BWP30P140LVT U51 ( .A1(n30), .A2(i_cmd[4]), .Z(n15) );
  NR2D1BWP30P140LVT U52 ( .A1(i_cmd[0]), .A2(n11), .ZN(n26) );
  INVD1BWP30P140LVT U53 ( .I(i_cmd[3]), .ZN(n12) );
  ND2OPTIBD2BWP30P140LVT U54 ( .A1(n26), .A2(n12), .ZN(n18) );
  NR2D1BWP30P140LVT U55 ( .A1(n18), .A2(n17), .ZN(n19) );
  ND2OPTPAD2BWP30P140LVT U56 ( .A1(n20), .A2(n19), .ZN(n49) );
  BUFFD4BWP30P140LVT U57 ( .I(n49), .Z(n145) );
  INVD1BWP30P140LVT U58 ( .I(i_cmd[7]), .ZN(n23) );
  INVD1BWP30P140LVT U59 ( .I(i_valid[7]), .ZN(n22) );
  NR4D0BWP30P140LVT U60 ( .A1(n23), .A2(n22), .A3(i_cmd[6]), .A4(i_cmd[5]), 
        .ZN(n24) );
  NR4D0BWP30P140LVT U61 ( .A1(n287), .A2(n129), .A3(n1), .A4(n268), .ZN(n45)
         );
  INVD1BWP30P140LVT U62 ( .I(i_cmd[4]), .ZN(n25) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n26), .A2(n25), .Z(n28) );
  ND2OPTIBD1BWP30P140LVT U64 ( .A1(n28), .A2(n27), .ZN(n40) );
  ND2D1BWP30P140LVT U65 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n29) );
  OR2D1BWP30P140LVT U66 ( .A1(n30), .A2(n29), .Z(n31) );
  INVD1BWP30P140LVT U67 ( .I(n4), .ZN(n175) );
  INVD1BWP30P140LVT U68 ( .I(n32), .ZN(n36) );
  ND2D1BWP30P140LVT U69 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n33) );
  NR2D1BWP30P140LVT U70 ( .A1(n33), .A2(i_cmd[0]), .ZN(n34) );
  NR2D1BWP30P140LVT U71 ( .A1(n175), .A2(n2), .ZN(n44) );
  INVD1BWP30P140LVT U72 ( .I(i_cmd[2]), .ZN(n37) );
  INR4D0BWP30P140LVT U73 ( .A1(i_valid[2]), .B1(i_cmd[1]), .B2(i_cmd[3]), .B3(
        n37), .ZN(n38) );
  INVD1BWP30P140LVT U74 ( .I(n38), .ZN(n39) );
  ND2D1BWP30P140LVT U75 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n41) );
  NR2D1BWP30P140LVT U76 ( .A1(n42), .A2(n41), .ZN(n43) );
  ND4D1BWP30P140LVT U77 ( .A1(n45), .A2(n44), .A3(n183), .A4(n46), .ZN(N402)
         );
  INVD2BWP30P140LVT U78 ( .I(n46), .ZN(n273) );
  AOI22D1BWP30P140LVT U79 ( .A1(n3), .A2(i_data_bus[76]), .B1(n273), .B2(
        i_data_bus[44]), .ZN(n58) );
  AOI22D1BWP30P140LVT U80 ( .A1(n274), .A2(i_data_bus[108]), .B1(n2), .B2(
        i_data_bus[140]), .ZN(n57) );
  INVD1BWP30P140LVT U81 ( .I(i_data_bus[236]), .ZN(n54) );
  BUFFD4BWP30P140LVT U82 ( .I(n48), .Z(n285) );
  INVD1BWP30P140LVT U83 ( .I(i_data_bus[204]), .ZN(n52) );
  INVD1BWP30P140LVT U84 ( .I(n49), .ZN(n50) );
  INVD2BWP30P140LVT U85 ( .I(n50), .ZN(n283) );
  INVD1BWP30P140LVT U86 ( .I(i_data_bus[172]), .ZN(n51) );
  OAI22D1BWP30P140LVT U87 ( .A1(n285), .A2(n52), .B1(n283), .B2(n51), .ZN(n53)
         );
  IAO21D1BWP30P140LVT U88 ( .A1(n137), .A2(n54), .B(n53), .ZN(n56) );
  ND4D1BWP30P140LVT U89 ( .A1(n58), .A2(n57), .A3(n56), .A4(n55), .ZN(N381) );
  AOI22D1BWP30P140LVT U90 ( .A1(n3), .A2(i_data_bus[70]), .B1(n273), .B2(
        i_data_bus[38]), .ZN(n65) );
  AOI22D1BWP30P140LVT U91 ( .A1(n274), .A2(i_data_bus[102]), .B1(n2), .B2(
        i_data_bus[134]), .ZN(n64) );
  INVD1BWP30P140LVT U92 ( .I(i_data_bus[198]), .ZN(n60) );
  INVD1BWP30P140LVT U93 ( .I(i_data_bus[166]), .ZN(n59) );
  OAI22D1BWP30P140LVT U94 ( .A1(n285), .A2(n60), .B1(n283), .B2(n59), .ZN(n61)
         );
  AOI21D1BWP30P140LVT U95 ( .A1(n268), .A2(i_data_bus[230]), .B(n61), .ZN(n63)
         );
  ND4D1BWP30P140LVT U96 ( .A1(n65), .A2(n64), .A3(n63), .A4(n62), .ZN(N375) );
  AOI22D1BWP30P140LVT U97 ( .A1(n3), .A2(i_data_bus[73]), .B1(n273), .B2(
        i_data_bus[41]), .ZN(n72) );
  AOI22D1BWP30P140LVT U98 ( .A1(n274), .A2(i_data_bus[105]), .B1(n2), .B2(
        i_data_bus[137]), .ZN(n71) );
  INVD1BWP30P140LVT U99 ( .I(i_data_bus[201]), .ZN(n67) );
  INVD1BWP30P140LVT U100 ( .I(i_data_bus[169]), .ZN(n66) );
  OAI22D1BWP30P140LVT U101 ( .A1(n285), .A2(n67), .B1(n283), .B2(n66), .ZN(n68) );
  AOI21D1BWP30P140LVT U102 ( .A1(n268), .A2(i_data_bus[233]), .B(n68), .ZN(n70) );
  ND4D1BWP30P140LVT U103 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(N378)
         );
  AOI22D1BWP30P140LVT U104 ( .A1(n3), .A2(i_data_bus[69]), .B1(n273), .B2(
        i_data_bus[37]), .ZN(n79) );
  AOI22D1BWP30P140LVT U105 ( .A1(n274), .A2(i_data_bus[101]), .B1(n2), .B2(
        i_data_bus[133]), .ZN(n78) );
  INVD1BWP30P140LVT U106 ( .I(i_data_bus[197]), .ZN(n74) );
  INVD1BWP30P140LVT U107 ( .I(i_data_bus[165]), .ZN(n73) );
  OAI22D1BWP30P140LVT U108 ( .A1(n285), .A2(n74), .B1(n283), .B2(n73), .ZN(n75) );
  AOI21D1BWP30P140LVT U109 ( .A1(n268), .A2(i_data_bus[229]), .B(n75), .ZN(n77) );
  ND4D1BWP30P140LVT U110 ( .A1(n79), .A2(n78), .A3(n77), .A4(n76), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U111 ( .A1(n3), .A2(i_data_bus[74]), .B1(n273), .B2(
        i_data_bus[42]), .ZN(n86) );
  AOI22D1BWP30P140LVT U112 ( .A1(n274), .A2(i_data_bus[106]), .B1(n2), .B2(
        i_data_bus[138]), .ZN(n85) );
  INVD1BWP30P140LVT U113 ( .I(i_data_bus[202]), .ZN(n81) );
  INVD1BWP30P140LVT U114 ( .I(i_data_bus[170]), .ZN(n80) );
  OAI22D1BWP30P140LVT U115 ( .A1(n285), .A2(n81), .B1(n283), .B2(n80), .ZN(n82) );
  AOI21D1BWP30P140LVT U116 ( .A1(n268), .A2(i_data_bus[234]), .B(n82), .ZN(n84) );
  ND4D1BWP30P140LVT U117 ( .A1(n86), .A2(n85), .A3(n84), .A4(n83), .ZN(N379)
         );
  AOI22D1BWP30P140LVT U118 ( .A1(n3), .A2(i_data_bus[75]), .B1(n273), .B2(
        i_data_bus[43]), .ZN(n93) );
  AOI22D1BWP30P140LVT U119 ( .A1(n274), .A2(i_data_bus[107]), .B1(n2), .B2(
        i_data_bus[139]), .ZN(n92) );
  INVD1BWP30P140LVT U120 ( .I(i_data_bus[203]), .ZN(n88) );
  INVD1BWP30P140LVT U121 ( .I(i_data_bus[171]), .ZN(n87) );
  OAI22D1BWP30P140LVT U122 ( .A1(n285), .A2(n88), .B1(n283), .B2(n87), .ZN(n89) );
  AOI21D1BWP30P140LVT U123 ( .A1(n268), .A2(i_data_bus[235]), .B(n89), .ZN(n91) );
  ND4D1BWP30P140LVT U124 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U125 ( .A1(n3), .A2(i_data_bus[66]), .B1(n273), .B2(
        i_data_bus[34]), .ZN(n100) );
  AOI22D1BWP30P140LVT U126 ( .A1(n274), .A2(i_data_bus[98]), .B1(n2), .B2(
        i_data_bus[130]), .ZN(n99) );
  INVD1BWP30P140LVT U127 ( .I(i_data_bus[194]), .ZN(n95) );
  INVD1BWP30P140LVT U128 ( .I(i_data_bus[162]), .ZN(n94) );
  OAI22D1BWP30P140LVT U129 ( .A1(n285), .A2(n95), .B1(n283), .B2(n94), .ZN(n96) );
  AOI21D1BWP30P140LVT U130 ( .A1(n268), .A2(i_data_bus[226]), .B(n96), .ZN(n98) );
  ND4D1BWP30P140LVT U131 ( .A1(n100), .A2(n99), .A3(n98), .A4(n97), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U132 ( .A1(n3), .A2(i_data_bus[71]), .B1(n273), .B2(
        i_data_bus[39]), .ZN(n107) );
  AOI22D1BWP30P140LVT U133 ( .A1(n274), .A2(i_data_bus[103]), .B1(n2), .B2(
        i_data_bus[135]), .ZN(n106) );
  INVD1BWP30P140LVT U134 ( .I(i_data_bus[199]), .ZN(n102) );
  INVD1BWP30P140LVT U135 ( .I(i_data_bus[167]), .ZN(n101) );
  OAI22D1BWP30P140LVT U136 ( .A1(n285), .A2(n102), .B1(n283), .B2(n101), .ZN(
        n103) );
  AOI21D1BWP30P140LVT U137 ( .A1(n268), .A2(i_data_bus[231]), .B(n103), .ZN(
        n105) );
  ND4D1BWP30P140LVT U138 ( .A1(n107), .A2(n106), .A3(n105), .A4(n104), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U139 ( .A1(n3), .A2(i_data_bus[65]), .B1(n273), .B2(
        i_data_bus[33]), .ZN(n114) );
  AOI22D1BWP30P140LVT U140 ( .A1(n274), .A2(i_data_bus[97]), .B1(n2), .B2(
        i_data_bus[129]), .ZN(n113) );
  INVD1BWP30P140LVT U141 ( .I(i_data_bus[193]), .ZN(n109) );
  INVD1BWP30P140LVT U142 ( .I(i_data_bus[161]), .ZN(n108) );
  OAI22D1BWP30P140LVT U143 ( .A1(n285), .A2(n109), .B1(n283), .B2(n108), .ZN(
        n110) );
  AOI21D1BWP30P140LVT U144 ( .A1(n268), .A2(i_data_bus[225]), .B(n110), .ZN(
        n112) );
  ND4D1BWP30P140LVT U145 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U146 ( .A1(n3), .A2(i_data_bus[68]), .B1(n273), .B2(
        i_data_bus[36]), .ZN(n121) );
  AOI22D1BWP30P140LVT U147 ( .A1(n274), .A2(i_data_bus[100]), .B1(n2), .B2(
        i_data_bus[132]), .ZN(n120) );
  INVD1BWP30P140LVT U148 ( .I(i_data_bus[196]), .ZN(n116) );
  INVD1BWP30P140LVT U149 ( .I(i_data_bus[164]), .ZN(n115) );
  OAI22D1BWP30P140LVT U150 ( .A1(n285), .A2(n116), .B1(n283), .B2(n115), .ZN(
        n117) );
  AOI21D1BWP30P140LVT U151 ( .A1(n268), .A2(i_data_bus[228]), .B(n117), .ZN(
        n119) );
  ND4D1BWP30P140LVT U152 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U153 ( .A1(n3), .A2(i_data_bus[67]), .B1(n273), .B2(
        i_data_bus[35]), .ZN(n128) );
  AOI22D1BWP30P140LVT U154 ( .A1(n274), .A2(i_data_bus[99]), .B1(n2), .B2(
        i_data_bus[131]), .ZN(n127) );
  INVD1BWP30P140LVT U155 ( .I(i_data_bus[195]), .ZN(n123) );
  INVD1BWP30P140LVT U156 ( .I(i_data_bus[163]), .ZN(n122) );
  OAI22D1BWP30P140LVT U157 ( .A1(n285), .A2(n123), .B1(n283), .B2(n122), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U158 ( .A1(n268), .A2(i_data_bus[227]), .B(n124), .ZN(
        n126) );
  ND4D1BWP30P140LVT U159 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(
        N372) );
  INVD2BWP30P140LVT U160 ( .I(n46), .ZN(n174) );
  AOI22D1BWP30P140LVT U161 ( .A1(n3), .A2(i_data_bus[95]), .B1(n174), .B2(
        i_data_bus[63]), .ZN(n136) );
  AOI22D1BWP30P140LVT U162 ( .A1(n175), .A2(i_data_bus[127]), .B1(n2), .B2(
        i_data_bus[159]), .ZN(n135) );
  INVD1BWP30P140LVT U163 ( .I(i_data_bus[223]), .ZN(n131) );
  INVD1BWP30P140LVT U164 ( .I(i_data_bus[191]), .ZN(n130) );
  OAI22D1BWP30P140LVT U165 ( .A1(n244), .A2(n131), .B1(n145), .B2(n130), .ZN(
        n132) );
  AOI21D1BWP30P140LVT U166 ( .A1(n268), .A2(i_data_bus[255]), .B(n132), .ZN(
        n134) );
  ND2D1BWP30P140LVT U167 ( .A1(n287), .A2(i_data_bus[31]), .ZN(n133) );
  ND4D1BWP30P140LVT U168 ( .A1(n136), .A2(n135), .A3(n134), .A4(n133), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U169 ( .A1(n3), .A2(i_data_bus[94]), .B1(n174), .B2(
        i_data_bus[62]), .ZN(n144) );
  AOI22D1BWP30P140LVT U170 ( .A1(n175), .A2(i_data_bus[126]), .B1(n2), .B2(
        i_data_bus[158]), .ZN(n143) );
  INVD2BWP30P140LVT U171 ( .I(n137), .ZN(n268) );
  INVD1BWP30P140LVT U172 ( .I(i_data_bus[222]), .ZN(n139) );
  INVD1BWP30P140LVT U173 ( .I(i_data_bus[190]), .ZN(n138) );
  OAI22D1BWP30P140LVT U174 ( .A1(n244), .A2(n139), .B1(n145), .B2(n138), .ZN(
        n140) );
  AOI21D1BWP30P140LVT U175 ( .A1(n268), .A2(i_data_bus[254]), .B(n140), .ZN(
        n142) );
  ND2D1BWP30P140LVT U176 ( .A1(n287), .A2(i_data_bus[30]), .ZN(n141) );
  ND4D1BWP30P140LVT U177 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U178 ( .A1(n3), .A2(i_data_bus[90]), .B1(n174), .B2(
        i_data_bus[58]), .ZN(n152) );
  AOI22D1BWP30P140LVT U179 ( .A1(n175), .A2(i_data_bus[122]), .B1(n2), .B2(
        i_data_bus[154]), .ZN(n151) );
  INVD1BWP30P140LVT U180 ( .I(i_data_bus[218]), .ZN(n147) );
  INVD4BWP30P140LVT U181 ( .I(n1), .ZN(n258) );
  INVD1BWP30P140LVT U182 ( .I(i_data_bus[186]), .ZN(n146) );
  OAI22D1BWP30P140LVT U183 ( .A1(n244), .A2(n147), .B1(n258), .B2(n146), .ZN(
        n148) );
  AOI21D1BWP30P140LVT U184 ( .A1(n268), .A2(i_data_bus[250]), .B(n148), .ZN(
        n150) );
  ND2D1BWP30P140LVT U185 ( .A1(n287), .A2(i_data_bus[26]), .ZN(n149) );
  ND4D1BWP30P140LVT U186 ( .A1(n152), .A2(n151), .A3(n150), .A4(n149), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U187 ( .A1(n3), .A2(i_data_bus[91]), .B1(n174), .B2(
        i_data_bus[59]), .ZN(n159) );
  AOI22D1BWP30P140LVT U188 ( .A1(n175), .A2(i_data_bus[123]), .B1(n2), .B2(
        i_data_bus[155]), .ZN(n158) );
  INVD1BWP30P140LVT U189 ( .I(i_data_bus[219]), .ZN(n154) );
  INVD1BWP30P140LVT U190 ( .I(i_data_bus[187]), .ZN(n153) );
  OAI22D1BWP30P140LVT U191 ( .A1(n244), .A2(n154), .B1(n258), .B2(n153), .ZN(
        n155) );
  AOI21D1BWP30P140LVT U192 ( .A1(n268), .A2(i_data_bus[251]), .B(n155), .ZN(
        n157) );
  ND2D1BWP30P140LVT U193 ( .A1(n287), .A2(i_data_bus[27]), .ZN(n156) );
  ND4D1BWP30P140LVT U194 ( .A1(n159), .A2(n158), .A3(n157), .A4(n156), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U195 ( .A1(n3), .A2(i_data_bus[93]), .B1(n174), .B2(
        i_data_bus[61]), .ZN(n166) );
  AOI22D1BWP30P140LVT U196 ( .A1(n175), .A2(i_data_bus[125]), .B1(n2), .B2(
        i_data_bus[157]), .ZN(n165) );
  INVD1BWP30P140LVT U197 ( .I(i_data_bus[221]), .ZN(n161) );
  INVD1BWP30P140LVT U198 ( .I(i_data_bus[189]), .ZN(n160) );
  OAI22D1BWP30P140LVT U199 ( .A1(n244), .A2(n161), .B1(n258), .B2(n160), .ZN(
        n162) );
  AOI21D1BWP30P140LVT U200 ( .A1(n268), .A2(i_data_bus[253]), .B(n162), .ZN(
        n164) );
  ND2D1BWP30P140LVT U201 ( .A1(n287), .A2(i_data_bus[29]), .ZN(n163) );
  ND4D1BWP30P140LVT U202 ( .A1(n166), .A2(n165), .A3(n164), .A4(n163), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U203 ( .A1(n3), .A2(i_data_bus[72]), .B1(n273), .B2(
        i_data_bus[40]), .ZN(n173) );
  AOI22D1BWP30P140LVT U204 ( .A1(n274), .A2(i_data_bus[104]), .B1(n2), .B2(
        i_data_bus[136]), .ZN(n172) );
  INVD1BWP30P140LVT U205 ( .I(i_data_bus[200]), .ZN(n168) );
  INVD1BWP30P140LVT U206 ( .I(i_data_bus[168]), .ZN(n167) );
  OAI22D1BWP30P140LVT U207 ( .A1(n285), .A2(n168), .B1(n283), .B2(n167), .ZN(
        n169) );
  ND4D1BWP30P140LVT U208 ( .A1(n173), .A2(n172), .A3(n171), .A4(n170), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U209 ( .A1(n3), .A2(i_data_bus[92]), .B1(n174), .B2(
        i_data_bus[60]), .ZN(n182) );
  AOI22D1BWP30P140LVT U210 ( .A1(n175), .A2(i_data_bus[124]), .B1(n2), .B2(
        i_data_bus[156]), .ZN(n181) );
  INVD1BWP30P140LVT U211 ( .I(i_data_bus[220]), .ZN(n177) );
  INVD1BWP30P140LVT U212 ( .I(i_data_bus[188]), .ZN(n176) );
  OAI22D1BWP30P140LVT U213 ( .A1(n244), .A2(n177), .B1(n258), .B2(n176), .ZN(
        n178) );
  AOI21D1BWP30P140LVT U214 ( .A1(n268), .A2(i_data_bus[252]), .B(n178), .ZN(
        n180) );
  ND2D1BWP30P140LVT U215 ( .A1(n287), .A2(i_data_bus[28]), .ZN(n179) );
  ND4D1BWP30P140LVT U216 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U217 ( .A1(n3), .A2(i_data_bus[81]), .B1(n174), .B2(
        i_data_bus[49]), .ZN(n192) );
  AOI22D1BWP30P140LVT U218 ( .A1(n281), .A2(i_data_bus[113]), .B1(n2), .B2(
        i_data_bus[145]), .ZN(n191) );
  INVD1BWP30P140LVT U219 ( .I(i_data_bus[209]), .ZN(n186) );
  INVD1BWP30P140LVT U220 ( .I(i_data_bus[177]), .ZN(n185) );
  OAI22D1BWP30P140LVT U221 ( .A1(n285), .A2(n186), .B1(n258), .B2(n185), .ZN(
        n187) );
  AOI21D1BWP30P140LVT U222 ( .A1(n268), .A2(i_data_bus[241]), .B(n187), .ZN(
        n190) );
  INVD2BWP30P140LVT U223 ( .I(n188), .ZN(n287) );
  ND2D1BWP30P140LVT U224 ( .A1(n287), .A2(i_data_bus[17]), .ZN(n189) );
  ND4D1BWP30P140LVT U225 ( .A1(n192), .A2(n191), .A3(n190), .A4(n189), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U226 ( .A1(n3), .A2(i_data_bus[79]), .B1(n174), .B2(
        i_data_bus[47]), .ZN(n199) );
  AOI22D1BWP30P140LVT U227 ( .A1(n281), .A2(i_data_bus[111]), .B1(n2), .B2(
        i_data_bus[143]), .ZN(n198) );
  INVD1BWP30P140LVT U228 ( .I(i_data_bus[207]), .ZN(n194) );
  INVD1BWP30P140LVT U229 ( .I(i_data_bus[175]), .ZN(n193) );
  OAI22D1BWP30P140LVT U230 ( .A1(n285), .A2(n194), .B1(n258), .B2(n193), .ZN(
        n195) );
  ND2D1BWP30P140LVT U231 ( .A1(n287), .A2(i_data_bus[15]), .ZN(n196) );
  ND4D1BWP30P140LVT U232 ( .A1(n199), .A2(n198), .A3(n197), .A4(n196), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U233 ( .A1(n3), .A2(i_data_bus[84]), .B1(n273), .B2(
        i_data_bus[52]), .ZN(n206) );
  AOI22D1BWP30P140LVT U234 ( .A1(n281), .A2(i_data_bus[116]), .B1(n2), .B2(
        i_data_bus[148]), .ZN(n205) );
  INVD1BWP30P140LVT U235 ( .I(i_data_bus[212]), .ZN(n201) );
  INVD1BWP30P140LVT U236 ( .I(i_data_bus[180]), .ZN(n200) );
  OAI22D1BWP30P140LVT U237 ( .A1(n285), .A2(n201), .B1(n258), .B2(n200), .ZN(
        n202) );
  AOI21D1BWP30P140LVT U238 ( .A1(n268), .A2(i_data_bus[244]), .B(n202), .ZN(
        n204) );
  ND2D1BWP30P140LVT U239 ( .A1(n287), .A2(i_data_bus[20]), .ZN(n203) );
  ND4D1BWP30P140LVT U240 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U241 ( .A1(n3), .A2(i_data_bus[82]), .B1(n174), .B2(
        i_data_bus[50]), .ZN(n213) );
  AOI22D1BWP30P140LVT U242 ( .A1(n281), .A2(i_data_bus[114]), .B1(n2), .B2(
        i_data_bus[146]), .ZN(n212) );
  INVD1BWP30P140LVT U243 ( .I(i_data_bus[210]), .ZN(n208) );
  INVD1BWP30P140LVT U244 ( .I(i_data_bus[178]), .ZN(n207) );
  OAI22D1BWP30P140LVT U245 ( .A1(n285), .A2(n208), .B1(n258), .B2(n207), .ZN(
        n209) );
  AOI21D1BWP30P140LVT U246 ( .A1(n268), .A2(i_data_bus[242]), .B(n209), .ZN(
        n211) );
  ND2D1BWP30P140LVT U247 ( .A1(n287), .A2(i_data_bus[18]), .ZN(n210) );
  ND4D1BWP30P140LVT U248 ( .A1(n213), .A2(n212), .A3(n211), .A4(n210), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U249 ( .A1(n3), .A2(i_data_bus[86]), .B1(n174), .B2(
        i_data_bus[54]), .ZN(n220) );
  AOI22D1BWP30P140LVT U250 ( .A1(n281), .A2(i_data_bus[118]), .B1(n2), .B2(
        i_data_bus[150]), .ZN(n219) );
  INVD1BWP30P140LVT U251 ( .I(i_data_bus[214]), .ZN(n215) );
  INVD1BWP30P140LVT U252 ( .I(i_data_bus[182]), .ZN(n214) );
  OAI22D1BWP30P140LVT U253 ( .A1(n285), .A2(n215), .B1(n258), .B2(n214), .ZN(
        n216) );
  AOI21D1BWP30P140LVT U254 ( .A1(n268), .A2(i_data_bus[246]), .B(n216), .ZN(
        n218) );
  ND2D1BWP30P140LVT U255 ( .A1(n287), .A2(i_data_bus[22]), .ZN(n217) );
  ND4D1BWP30P140LVT U256 ( .A1(n220), .A2(n219), .A3(n218), .A4(n217), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U257 ( .A1(n3), .A2(i_data_bus[85]), .B1(n174), .B2(
        i_data_bus[53]), .ZN(n227) );
  AOI22D1BWP30P140LVT U258 ( .A1(n281), .A2(i_data_bus[117]), .B1(n2), .B2(
        i_data_bus[149]), .ZN(n226) );
  INVD1BWP30P140LVT U259 ( .I(i_data_bus[213]), .ZN(n222) );
  INVD1BWP30P140LVT U260 ( .I(i_data_bus[181]), .ZN(n221) );
  OAI22D1BWP30P140LVT U261 ( .A1(n285), .A2(n222), .B1(n258), .B2(n221), .ZN(
        n223) );
  AOI21D1BWP30P140LVT U262 ( .A1(n268), .A2(i_data_bus[245]), .B(n223), .ZN(
        n225) );
  ND2D1BWP30P140LVT U263 ( .A1(n287), .A2(i_data_bus[21]), .ZN(n224) );
  ND4D1BWP30P140LVT U264 ( .A1(n227), .A2(n226), .A3(n225), .A4(n224), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U265 ( .A1(n3), .A2(i_data_bus[83]), .B1(n174), .B2(
        i_data_bus[51]), .ZN(n234) );
  AOI22D1BWP30P140LVT U266 ( .A1(n281), .A2(i_data_bus[115]), .B1(n2), .B2(
        i_data_bus[147]), .ZN(n233) );
  INVD1BWP30P140LVT U267 ( .I(i_data_bus[211]), .ZN(n229) );
  INVD1BWP30P140LVT U268 ( .I(i_data_bus[179]), .ZN(n228) );
  OAI22D1BWP30P140LVT U269 ( .A1(n285), .A2(n229), .B1(n258), .B2(n228), .ZN(
        n230) );
  AOI21D1BWP30P140LVT U270 ( .A1(n268), .A2(i_data_bus[243]), .B(n230), .ZN(
        n232) );
  ND2D1BWP30P140LVT U271 ( .A1(n287), .A2(i_data_bus[19]), .ZN(n231) );
  ND4D1BWP30P140LVT U272 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U273 ( .A1(n3), .A2(i_data_bus[87]), .B1(n174), .B2(
        i_data_bus[55]), .ZN(n241) );
  AOI22D1BWP30P140LVT U274 ( .A1(n281), .A2(i_data_bus[119]), .B1(n2), .B2(
        i_data_bus[151]), .ZN(n240) );
  INVD1BWP30P140LVT U275 ( .I(i_data_bus[215]), .ZN(n236) );
  INVD1BWP30P140LVT U276 ( .I(i_data_bus[183]), .ZN(n235) );
  OAI22D1BWP30P140LVT U277 ( .A1(n285), .A2(n236), .B1(n258), .B2(n235), .ZN(
        n237) );
  AOI21D1BWP30P140LVT U278 ( .A1(n268), .A2(i_data_bus[247]), .B(n237), .ZN(
        n239) );
  ND2D1BWP30P140LVT U279 ( .A1(n287), .A2(i_data_bus[23]), .ZN(n238) );
  ND4D1BWP30P140LVT U280 ( .A1(n241), .A2(n240), .A3(n239), .A4(n238), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U281 ( .A1(n3), .A2(i_data_bus[89]), .B1(n273), .B2(
        i_data_bus[57]), .ZN(n249) );
  AOI22D1BWP30P140LVT U282 ( .A1(n281), .A2(i_data_bus[121]), .B1(n2), .B2(
        i_data_bus[153]), .ZN(n248) );
  INVD1BWP30P140LVT U283 ( .I(i_data_bus[217]), .ZN(n243) );
  INVD1BWP30P140LVT U284 ( .I(i_data_bus[185]), .ZN(n242) );
  OAI22D1BWP30P140LVT U285 ( .A1(n244), .A2(n243), .B1(n258), .B2(n242), .ZN(
        n245) );
  AOI21D1BWP30P140LVT U286 ( .A1(n268), .A2(i_data_bus[249]), .B(n245), .ZN(
        n247) );
  ND2D1BWP30P140LVT U287 ( .A1(n287), .A2(i_data_bus[25]), .ZN(n246) );
  ND4D1BWP30P140LVT U288 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U289 ( .A1(n3), .A2(i_data_bus[88]), .B1(n174), .B2(
        i_data_bus[56]), .ZN(n256) );
  AOI22D1BWP30P140LVT U290 ( .A1(n281), .A2(i_data_bus[120]), .B1(n2), .B2(
        i_data_bus[152]), .ZN(n255) );
  INVD1BWP30P140LVT U291 ( .I(i_data_bus[216]), .ZN(n251) );
  INVD1BWP30P140LVT U292 ( .I(i_data_bus[184]), .ZN(n250) );
  OAI22D1BWP30P140LVT U293 ( .A1(n285), .A2(n251), .B1(n258), .B2(n250), .ZN(
        n252) );
  AOI21D1BWP30P140LVT U294 ( .A1(n268), .A2(i_data_bus[248]), .B(n252), .ZN(
        n254) );
  ND2D1BWP30P140LVT U295 ( .A1(n287), .A2(i_data_bus[24]), .ZN(n253) );
  ND4D1BWP30P140LVT U296 ( .A1(n256), .A2(n255), .A3(n254), .A4(n253), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U297 ( .A1(n3), .A2(i_data_bus[80]), .B1(n174), .B2(
        i_data_bus[48]), .ZN(n264) );
  AOI22D1BWP30P140LVT U298 ( .A1(n281), .A2(i_data_bus[112]), .B1(n2), .B2(
        i_data_bus[144]), .ZN(n263) );
  INVD1BWP30P140LVT U299 ( .I(i_data_bus[208]), .ZN(n259) );
  INVD1BWP30P140LVT U300 ( .I(i_data_bus[176]), .ZN(n257) );
  OAI22D1BWP30P140LVT U301 ( .A1(n285), .A2(n259), .B1(n258), .B2(n257), .ZN(
        n260) );
  AOI21D1BWP30P140LVT U302 ( .A1(n268), .A2(i_data_bus[240]), .B(n260), .ZN(
        n262) );
  ND2D1BWP30P140LVT U303 ( .A1(n287), .A2(i_data_bus[16]), .ZN(n261) );
  ND4D1BWP30P140LVT U304 ( .A1(n264), .A2(n263), .A3(n262), .A4(n261), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U305 ( .A1(n3), .A2(i_data_bus[78]), .B1(n174), .B2(
        i_data_bus[46]), .ZN(n272) );
  AOI22D1BWP30P140LVT U306 ( .A1(n281), .A2(i_data_bus[110]), .B1(n2), .B2(
        i_data_bus[142]), .ZN(n271) );
  INVD1BWP30P140LVT U307 ( .I(i_data_bus[206]), .ZN(n266) );
  INVD1BWP30P140LVT U308 ( .I(i_data_bus[174]), .ZN(n265) );
  OAI22D1BWP30P140LVT U309 ( .A1(n285), .A2(n266), .B1(n283), .B2(n265), .ZN(
        n267) );
  ND2D1BWP30P140LVT U310 ( .A1(n287), .A2(i_data_bus[14]), .ZN(n269) );
  ND4D1BWP30P140LVT U311 ( .A1(n272), .A2(n271), .A3(n270), .A4(n269), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U312 ( .A1(n3), .A2(i_data_bus[64]), .B1(n273), .B2(
        i_data_bus[32]), .ZN(n280) );
  AOI22D1BWP30P140LVT U313 ( .A1(n274), .A2(i_data_bus[96]), .B1(n2), .B2(
        i_data_bus[128]), .ZN(n279) );
  INR2D1BWP30P140LVT U314 ( .A1(i_data_bus[192]), .B1(n285), .ZN(n276) );
  INR2D1BWP30P140LVT U315 ( .A1(i_data_bus[160]), .B1(n283), .ZN(n275) );
  AOI211D1BWP30P140LVT U316 ( .A1(i_data_bus[224]), .A2(n268), .B(n276), .C(
        n275), .ZN(n278) );
  ND2D1BWP30P140LVT U317 ( .A1(n287), .A2(i_data_bus[0]), .ZN(n277) );
  ND4D1BWP30P140LVT U318 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U319 ( .A1(n3), .A2(i_data_bus[77]), .B1(n174), .B2(
        i_data_bus[45]), .ZN(n291) );
  AOI22D1BWP30P140LVT U320 ( .A1(n281), .A2(i_data_bus[109]), .B1(n2), .B2(
        i_data_bus[141]), .ZN(n290) );
  INVD1BWP30P140LVT U321 ( .I(i_data_bus[205]), .ZN(n284) );
  INVD1BWP30P140LVT U322 ( .I(i_data_bus[173]), .ZN(n282) );
  OAI22D1BWP30P140LVT U323 ( .A1(n285), .A2(n284), .B1(n283), .B2(n282), .ZN(
        n286) );
  AOI21D1BWP30P140LVT U324 ( .A1(n268), .A2(i_data_bus[237]), .B(n286), .ZN(
        n289) );
  ND2D1BWP30P140LVT U325 ( .A1(n287), .A2(i_data_bus[13]), .ZN(n288) );
  ND4D1BWP30P140LVT U326 ( .A1(n291), .A2(n290), .A3(n289), .A4(n288), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_12 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  DFD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  AOI22D1BWP30P140LVT U3 ( .A1(n4), .A2(i_data_bus[127]), .B1(n274), .B2(
        i_data_bus[159]), .ZN(n71) );
  INVD3BWP30P140LVT U4 ( .I(n73), .ZN(n1) );
  INR2D6BWP30P140LVT U5 ( .A1(n25), .B1(n19), .ZN(n242) );
  CKND2D3BWP30P140LVT U6 ( .A1(n23), .A2(n25), .ZN(n116) );
  INVD4BWP30P140LVT U7 ( .I(n56), .ZN(n2) );
  NR2OPTPAD2BWP30P140LVT U8 ( .A1(n20), .A2(i_cmd[5]), .ZN(n31) );
  OR2D4BWP30P140LVT U9 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n20) );
  ND2OPTIBD2BWP30P140LVT U10 ( .A1(n5), .A2(n9), .ZN(n36) );
  NR2D1BWP30P140LVT U11 ( .A1(n42), .A2(i_cmd[1]), .ZN(n9) );
  ND2OPTIBD2BWP30P140LVT U12 ( .A1(n6), .A2(n31), .ZN(n43) );
  INVD1BWP30P140LVT U13 ( .I(n38), .ZN(n48) );
  INR2D1BWP30P140LVT U14 ( .A1(n37), .B1(n36), .ZN(n38) );
  ND2D1BWP30P140LVT U15 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n35) );
  INVD1BWP30P140LVT U16 ( .I(n11), .ZN(n68) );
  INR2D1BWP30P140LVT U17 ( .A1(n10), .B1(n36), .ZN(n11) );
  ND2D1BWP30P140LVT U18 ( .A1(n242), .A2(i_data_bus[194]), .ZN(n243) );
  ND2D1BWP30P140LVT U19 ( .A1(n242), .A2(i_data_bus[195]), .ZN(n235) );
  INVD2BWP30P140LVT U20 ( .I(n48), .ZN(n257) );
  ND2D1BWP30P140LVT U21 ( .A1(n242), .A2(i_data_bus[207]), .ZN(n214) );
  AOI21D1BWP30P140LVT U22 ( .A1(n1), .A2(i_data_bus[245]), .B(n176), .ZN(n178)
         );
  INVD3BWP30P140LVT U23 ( .I(n48), .ZN(n274) );
  ND2D1BWP30P140LVT U24 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n32) );
  INR2D4BWP30P140LVT U25 ( .A1(n44), .B1(n43), .ZN(n273) );
  NR2D3BWP30P140LVT U26 ( .A1(n43), .A2(n34), .ZN(n4) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n31), .A2(n13), .Z(n5) );
  INVD1BWP30P140LVT U28 ( .I(n28), .ZN(n73) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n30), .A2(n29), .Z(n6) );
  INR2D1BWP30P140LVT U30 ( .A1(n40), .B1(n43), .ZN(n145) );
  INVD1BWP30P140LVT U31 ( .I(i_cmd[0]), .ZN(n7) );
  INR3D0BWP30P140LVT U32 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n7), .ZN(n10)
         );
  INVD1BWP30P140LVT U33 ( .I(rst), .ZN(n8) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n8), .A2(i_en), .Z(n13) );
  OR2D1BWP30P140LVT U35 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n42) );
  INVD2BWP30P140LVT U36 ( .I(n68), .ZN(n230) );
  INVD1BWP30P140LVT U37 ( .I(i_cmd[4]), .ZN(n30) );
  INVD1BWP30P140LVT U38 ( .I(i_cmd[3]), .ZN(n12) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(n30), .A2(n12), .ZN(n16) );
  INVD1BWP30P140LVT U40 ( .I(n13), .ZN(n14) );
  NR2D1BWP30P140LVT U41 ( .A1(i_cmd[0]), .A2(n14), .ZN(n29) );
  INVD1BWP30P140LVT U42 ( .I(n29), .ZN(n15) );
  OR2D2BWP30P140LVT U43 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n33) );
  NR3D3BWP30P140LVT U44 ( .A1(n16), .A2(n15), .A3(n33), .ZN(n25) );
  ND2D1BWP30P140LVT U45 ( .A1(i_cmd[6]), .A2(i_valid[6]), .ZN(n18) );
  NR2D1BWP30P140LVT U46 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n17) );
  IND2D1BWP30P140LVT U47 ( .A1(n18), .B1(n17), .ZN(n19) );
  INVD1BWP30P140LVT U48 ( .I(n20), .ZN(n22) );
  ND2D1BWP30P140LVT U49 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n21) );
  INR2D1BWP30P140LVT U50 ( .A1(n22), .B1(n21), .ZN(n23) );
  INVD1BWP30P140LVT U51 ( .I(n116), .ZN(n57) );
  INVD1BWP30P140LVT U52 ( .I(i_cmd[7]), .ZN(n24) );
  INR4D0BWP30P140LVT U53 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n24), .ZN(n27) );
  INVD1BWP30P140LVT U54 ( .I(n25), .ZN(n26) );
  INR2D1BWP30P140LVT U55 ( .A1(n27), .B1(n26), .ZN(n28) );
  NR4D0BWP30P140LVT U56 ( .A1(n230), .A2(n242), .A3(n57), .A4(n1), .ZN(n47) );
  OR2D1BWP30P140LVT U57 ( .A1(n33), .A2(n32), .Z(n34) );
  NR2D1BWP30P140LVT U58 ( .A1(n35), .A2(i_cmd[0]), .ZN(n37) );
  NR2D1BWP30P140LVT U59 ( .A1(n4), .A2(n274), .ZN(n46) );
  INVD1BWP30P140LVT U60 ( .I(i_cmd[2]), .ZN(n39) );
  INR4D0BWP30P140LVT U61 ( .A1(i_valid[2]), .B1(i_cmd[1]), .B2(i_cmd[3]), .B3(
        n39), .ZN(n40) );
  INVD1BWP30P140LVT U62 ( .I(n145), .ZN(n56) );
  ND2D1BWP30P140LVT U63 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n41) );
  NR2D1BWP30P140LVT U64 ( .A1(n42), .A2(n41), .ZN(n44) );
  INVD1BWP30P140LVT U65 ( .I(n273), .ZN(n45) );
  ND4D1BWP30P140LVT U66 ( .A1(n47), .A2(n46), .A3(n56), .A4(n45), .ZN(N402) );
  AOI22D1BWP30P140LVT U67 ( .A1(n2), .A2(i_data_bus[70]), .B1(n273), .B2(
        i_data_bus[38]), .ZN(n55) );
  AOI22D1BWP30P140LVT U68 ( .A1(n4), .A2(i_data_bus[102]), .B1(n257), .B2(
        i_data_bus[134]), .ZN(n54) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[166]), .ZN(n50) );
  INVD3BWP30P140LVT U70 ( .I(n242), .ZN(n259) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[198]), .ZN(n49) );
  OAI22D1BWP30P140LVT U72 ( .A1(n215), .A2(n50), .B1(n259), .B2(n49), .ZN(n51)
         );
  AOI21D1BWP30P140LVT U73 ( .A1(n1), .A2(i_data_bus[230]), .B(n51), .ZN(n53)
         );
  INVD2BWP30P140LVT U74 ( .I(n68), .ZN(n252) );
  ND2D1BWP30P140LVT U75 ( .A1(n252), .A2(i_data_bus[6]), .ZN(n52) );
  ND4D1BWP30P140LVT U76 ( .A1(n55), .A2(n54), .A3(n53), .A4(n52), .ZN(N375) );
  AOI22D1BWP30P140LVT U77 ( .A1(n2), .A2(i_data_bus[94]), .B1(n273), .B2(
        i_data_bus[62]), .ZN(n64) );
  AOI22D1BWP30P140LVT U78 ( .A1(n4), .A2(i_data_bus[126]), .B1(n274), .B2(
        i_data_bus[158]), .ZN(n63) );
  INVD1BWP30P140LVT U79 ( .I(i_data_bus[222]), .ZN(n59) );
  INVD1BWP30P140LVT U80 ( .I(n57), .ZN(n189) );
  INVD1BWP30P140LVT U81 ( .I(i_data_bus[190]), .ZN(n58) );
  OAI22D1BWP30P140LVT U82 ( .A1(n259), .A2(n59), .B1(n189), .B2(n58), .ZN(n60)
         );
  AOI21D1BWP30P140LVT U83 ( .A1(n1), .A2(i_data_bus[254]), .B(n60), .ZN(n62)
         );
  ND2D1BWP30P140LVT U84 ( .A1(n252), .A2(i_data_bus[30]), .ZN(n61) );
  ND4D1BWP30P140LVT U85 ( .A1(n63), .A2(n64), .A3(n62), .A4(n61), .ZN(N399) );
  AOI22D1BWP30P140LVT U86 ( .A1(n2), .A2(i_data_bus[95]), .B1(n273), .B2(
        i_data_bus[63]), .ZN(n72) );
  INVD1BWP30P140LVT U87 ( .I(i_data_bus[223]), .ZN(n66) );
  INVD1BWP30P140LVT U88 ( .I(i_data_bus[191]), .ZN(n65) );
  OAI22D1BWP30P140LVT U89 ( .A1(n259), .A2(n66), .B1(n189), .B2(n65), .ZN(n67)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n1), .A2(i_data_bus[255]), .B(n67), .ZN(n70)
         );
  INVD2BWP30P140LVT U91 ( .I(n68), .ZN(n279) );
  ND2D1BWP30P140LVT U92 ( .A1(n279), .A2(i_data_bus[31]), .ZN(n69) );
  ND4D1BWP30P140LVT U93 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(N400) );
  AOI22D1BWP30P140LVT U94 ( .A1(n2), .A2(i_data_bus[72]), .B1(n273), .B2(
        i_data_bus[40]), .ZN(n80) );
  AOI22D1BWP30P140LVT U95 ( .A1(n4), .A2(i_data_bus[104]), .B1(n257), .B2(
        i_data_bus[136]), .ZN(n79) );
  INVD3BWP30P140LVT U96 ( .I(n242), .ZN(n277) );
  INVD1BWP30P140LVT U97 ( .I(i_data_bus[200]), .ZN(n75) );
  INVD1BWP30P140LVT U98 ( .I(i_data_bus[168]), .ZN(n74) );
  OAI22D1BWP30P140LVT U99 ( .A1(n277), .A2(n75), .B1(n215), .B2(n74), .ZN(n76)
         );
  AOI21D1BWP30P140LVT U100 ( .A1(n1), .A2(i_data_bus[232]), .B(n76), .ZN(n78)
         );
  ND2D1BWP30P140LVT U101 ( .A1(n252), .A2(i_data_bus[8]), .ZN(n77) );
  ND4D1BWP30P140LVT U102 ( .A1(n80), .A2(n79), .A3(n78), .A4(n77), .ZN(N377)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n2), .A2(i_data_bus[76]), .B1(n273), .B2(
        i_data_bus[44]), .ZN(n87) );
  AOI22D1BWP30P140LVT U104 ( .A1(n4), .A2(i_data_bus[108]), .B1(n257), .B2(
        i_data_bus[140]), .ZN(n86) );
  INVD1BWP30P140LVT U105 ( .I(i_data_bus[204]), .ZN(n82) );
  INVD1BWP30P140LVT U106 ( .I(i_data_bus[172]), .ZN(n81) );
  OAI22D1BWP30P140LVT U107 ( .A1(n277), .A2(n82), .B1(n215), .B2(n81), .ZN(n83) );
  AOI21D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[236]), .B(n83), .ZN(n85)
         );
  ND2D1BWP30P140LVT U109 ( .A1(n279), .A2(i_data_bus[12]), .ZN(n84) );
  ND4D1BWP30P140LVT U110 ( .A1(n87), .A2(n86), .A3(n85), .A4(n84), .ZN(N381)
         );
  AOI22D1BWP30P140LVT U111 ( .A1(n2), .A2(i_data_bus[75]), .B1(n273), .B2(
        i_data_bus[43]), .ZN(n94) );
  AOI22D1BWP30P140LVT U112 ( .A1(n4), .A2(i_data_bus[107]), .B1(n257), .B2(
        i_data_bus[139]), .ZN(n93) );
  INVD1BWP30P140LVT U113 ( .I(i_data_bus[203]), .ZN(n89) );
  INVD1BWP30P140LVT U114 ( .I(i_data_bus[171]), .ZN(n88) );
  OAI22D1BWP30P140LVT U115 ( .A1(n277), .A2(n89), .B1(n215), .B2(n88), .ZN(n90) );
  AOI21D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[235]), .B(n90), .ZN(n92)
         );
  ND2D1BWP30P140LVT U117 ( .A1(n252), .A2(i_data_bus[11]), .ZN(n91) );
  ND4D1BWP30P140LVT U118 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U119 ( .A1(n2), .A2(i_data_bus[74]), .B1(n273), .B2(
        i_data_bus[42]), .ZN(n101) );
  AOI22D1BWP30P140LVT U120 ( .A1(n4), .A2(i_data_bus[106]), .B1(n257), .B2(
        i_data_bus[138]), .ZN(n100) );
  INVD1BWP30P140LVT U121 ( .I(i_data_bus[202]), .ZN(n96) );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[170]), .ZN(n95) );
  OAI22D1BWP30P140LVT U123 ( .A1(n277), .A2(n96), .B1(n215), .B2(n95), .ZN(n97) );
  AOI21D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[234]), .B(n97), .ZN(n99)
         );
  ND2D1BWP30P140LVT U125 ( .A1(n230), .A2(i_data_bus[10]), .ZN(n98) );
  ND4D1BWP30P140LVT U126 ( .A1(n101), .A2(n100), .A3(n99), .A4(n98), .ZN(N379)
         );
  AOI22D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[73]), .B1(n273), .B2(
        i_data_bus[41]), .ZN(n108) );
  AOI22D1BWP30P140LVT U128 ( .A1(n4), .A2(i_data_bus[105]), .B1(n257), .B2(
        i_data_bus[137]), .ZN(n107) );
  INVD1BWP30P140LVT U129 ( .I(i_data_bus[201]), .ZN(n103) );
  INVD1BWP30P140LVT U130 ( .I(i_data_bus[169]), .ZN(n102) );
  OAI22D1BWP30P140LVT U131 ( .A1(n277), .A2(n103), .B1(n215), .B2(n102), .ZN(
        n104) );
  AOI21D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[233]), .B(n104), .ZN(n106) );
  ND2D1BWP30P140LVT U133 ( .A1(n230), .A2(i_data_bus[9]), .ZN(n105) );
  ND4D1BWP30P140LVT U134 ( .A1(n108), .A2(n107), .A3(n106), .A4(n105), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[71]), .B1(n273), .B2(
        i_data_bus[39]), .ZN(n115) );
  AOI22D1BWP30P140LVT U136 ( .A1(n4), .A2(i_data_bus[103]), .B1(n257), .B2(
        i_data_bus[135]), .ZN(n114) );
  INVD1BWP30P140LVT U137 ( .I(i_data_bus[199]), .ZN(n110) );
  INVD1BWP30P140LVT U138 ( .I(i_data_bus[167]), .ZN(n109) );
  OAI22D1BWP30P140LVT U139 ( .A1(n277), .A2(n110), .B1(n215), .B2(n109), .ZN(
        n111) );
  AOI21D1BWP30P140LVT U140 ( .A1(n1), .A2(i_data_bus[231]), .B(n111), .ZN(n113) );
  ND2D1BWP30P140LVT U141 ( .A1(n230), .A2(i_data_bus[7]), .ZN(n112) );
  ND4D1BWP30P140LVT U142 ( .A1(n115), .A2(n114), .A3(n113), .A4(n112), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U143 ( .A1(n2), .A2(i_data_bus[93]), .B1(n273), .B2(
        i_data_bus[61]), .ZN(n123) );
  AOI22D1BWP30P140LVT U144 ( .A1(n4), .A2(i_data_bus[125]), .B1(n274), .B2(
        i_data_bus[157]), .ZN(n122) );
  INVD1BWP30P140LVT U145 ( .I(i_data_bus[221]), .ZN(n118) );
  BUFFD4BWP30P140LVT U146 ( .I(n116), .Z(n215) );
  INVD1BWP30P140LVT U147 ( .I(i_data_bus[189]), .ZN(n117) );
  OAI22D1BWP30P140LVT U148 ( .A1(n259), .A2(n118), .B1(n215), .B2(n117), .ZN(
        n119) );
  AOI21D1BWP30P140LVT U149 ( .A1(n1), .A2(i_data_bus[253]), .B(n119), .ZN(n121) );
  ND2D1BWP30P140LVT U150 ( .A1(n252), .A2(i_data_bus[29]), .ZN(n120) );
  ND4D1BWP30P140LVT U151 ( .A1(n122), .A2(n123), .A3(n121), .A4(n120), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U152 ( .A1(n2), .A2(i_data_bus[92]), .B1(n273), .B2(
        i_data_bus[60]), .ZN(n130) );
  AOI22D1BWP30P140LVT U153 ( .A1(n4), .A2(i_data_bus[124]), .B1(n274), .B2(
        i_data_bus[156]), .ZN(n129) );
  INVD1BWP30P140LVT U154 ( .I(i_data_bus[220]), .ZN(n125) );
  INVD1BWP30P140LVT U155 ( .I(i_data_bus[188]), .ZN(n124) );
  OAI22D1BWP30P140LVT U156 ( .A1(n259), .A2(n125), .B1(n215), .B2(n124), .ZN(
        n126) );
  AOI21D1BWP30P140LVT U157 ( .A1(n1), .A2(i_data_bus[252]), .B(n126), .ZN(n128) );
  ND2D1BWP30P140LVT U158 ( .A1(n230), .A2(i_data_bus[28]), .ZN(n127) );
  ND4D1BWP30P140LVT U159 ( .A1(n129), .A2(n130), .A3(n128), .A4(n127), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U160 ( .A1(n2), .A2(i_data_bus[91]), .B1(n273), .B2(
        i_data_bus[59]), .ZN(n137) );
  AOI22D1BWP30P140LVT U161 ( .A1(n4), .A2(i_data_bus[123]), .B1(n274), .B2(
        i_data_bus[155]), .ZN(n136) );
  INVD1BWP30P140LVT U162 ( .I(i_data_bus[219]), .ZN(n132) );
  INVD1BWP30P140LVT U163 ( .I(i_data_bus[187]), .ZN(n131) );
  OAI22D1BWP30P140LVT U164 ( .A1(n259), .A2(n132), .B1(n215), .B2(n131), .ZN(
        n133) );
  AOI21D1BWP30P140LVT U165 ( .A1(n1), .A2(i_data_bus[251]), .B(n133), .ZN(n135) );
  ND2D1BWP30P140LVT U166 ( .A1(n230), .A2(i_data_bus[27]), .ZN(n134) );
  ND4D1BWP30P140LVT U167 ( .A1(n136), .A2(n137), .A3(n135), .A4(n134), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U168 ( .A1(n2), .A2(i_data_bus[90]), .B1(n273), .B2(
        i_data_bus[58]), .ZN(n144) );
  AOI22D1BWP30P140LVT U169 ( .A1(n4), .A2(i_data_bus[122]), .B1(n274), .B2(
        i_data_bus[154]), .ZN(n143) );
  INVD1BWP30P140LVT U170 ( .I(i_data_bus[218]), .ZN(n139) );
  INVD1BWP30P140LVT U171 ( .I(i_data_bus[186]), .ZN(n138) );
  OAI22D1BWP30P140LVT U172 ( .A1(n259), .A2(n139), .B1(n215), .B2(n138), .ZN(
        n140) );
  AOI21D1BWP30P140LVT U173 ( .A1(n1), .A2(i_data_bus[250]), .B(n140), .ZN(n142) );
  ND2D1BWP30P140LVT U174 ( .A1(n279), .A2(i_data_bus[26]), .ZN(n141) );
  ND4D1BWP30P140LVT U175 ( .A1(n143), .A2(n144), .A3(n142), .A4(n141), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U176 ( .A1(n2), .A2(i_data_bus[89]), .B1(n273), .B2(
        i_data_bus[57]), .ZN(n152) );
  AOI22D1BWP30P140LVT U177 ( .A1(n4), .A2(i_data_bus[121]), .B1(n274), .B2(
        i_data_bus[153]), .ZN(n151) );
  INVD1BWP30P140LVT U178 ( .I(i_data_bus[217]), .ZN(n147) );
  INVD1BWP30P140LVT U179 ( .I(i_data_bus[185]), .ZN(n146) );
  OAI22D1BWP30P140LVT U180 ( .A1(n259), .A2(n147), .B1(n215), .B2(n146), .ZN(
        n148) );
  AOI21D1BWP30P140LVT U181 ( .A1(n1), .A2(i_data_bus[249]), .B(n148), .ZN(n150) );
  ND2D1BWP30P140LVT U182 ( .A1(n279), .A2(i_data_bus[25]), .ZN(n149) );
  ND4D1BWP30P140LVT U183 ( .A1(n151), .A2(n152), .A3(n150), .A4(n149), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U184 ( .A1(n2), .A2(i_data_bus[88]), .B1(n273), .B2(
        i_data_bus[56]), .ZN(n159) );
  AOI22D1BWP30P140LVT U185 ( .A1(n4), .A2(i_data_bus[120]), .B1(n274), .B2(
        i_data_bus[152]), .ZN(n158) );
  INVD1BWP30P140LVT U186 ( .I(i_data_bus[216]), .ZN(n154) );
  INVD1BWP30P140LVT U187 ( .I(i_data_bus[184]), .ZN(n153) );
  OAI22D1BWP30P140LVT U188 ( .A1(n277), .A2(n154), .B1(n215), .B2(n153), .ZN(
        n155) );
  AOI21D1BWP30P140LVT U189 ( .A1(n1), .A2(i_data_bus[248]), .B(n155), .ZN(n157) );
  ND2D1BWP30P140LVT U190 ( .A1(n230), .A2(i_data_bus[24]), .ZN(n156) );
  ND4D1BWP30P140LVT U191 ( .A1(n158), .A2(n159), .A3(n157), .A4(n156), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U192 ( .A1(n2), .A2(i_data_bus[87]), .B1(n273), .B2(
        i_data_bus[55]), .ZN(n166) );
  AOI22D1BWP30P140LVT U193 ( .A1(n4), .A2(i_data_bus[119]), .B1(n274), .B2(
        i_data_bus[151]), .ZN(n165) );
  INVD1BWP30P140LVT U194 ( .I(i_data_bus[215]), .ZN(n161) );
  INVD1BWP30P140LVT U195 ( .I(i_data_bus[183]), .ZN(n160) );
  OAI22D1BWP30P140LVT U196 ( .A1(n277), .A2(n161), .B1(n215), .B2(n160), .ZN(
        n162) );
  AOI21D1BWP30P140LVT U197 ( .A1(n1), .A2(i_data_bus[247]), .B(n162), .ZN(n164) );
  ND2D1BWP30P140LVT U198 ( .A1(n230), .A2(i_data_bus[23]), .ZN(n163) );
  ND4D1BWP30P140LVT U199 ( .A1(n165), .A2(n166), .A3(n164), .A4(n163), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U200 ( .A1(n2), .A2(i_data_bus[86]), .B1(n273), .B2(
        i_data_bus[54]), .ZN(n173) );
  AOI22D1BWP30P140LVT U201 ( .A1(n4), .A2(i_data_bus[118]), .B1(n274), .B2(
        i_data_bus[150]), .ZN(n172) );
  INVD1BWP30P140LVT U202 ( .I(i_data_bus[214]), .ZN(n168) );
  INVD1BWP30P140LVT U203 ( .I(i_data_bus[182]), .ZN(n167) );
  OAI22D1BWP30P140LVT U204 ( .A1(n277), .A2(n168), .B1(n215), .B2(n167), .ZN(
        n169) );
  AOI21D1BWP30P140LVT U205 ( .A1(n1), .A2(i_data_bus[246]), .B(n169), .ZN(n171) );
  ND2D1BWP30P140LVT U206 ( .A1(n252), .A2(i_data_bus[22]), .ZN(n170) );
  ND4D1BWP30P140LVT U207 ( .A1(n172), .A2(n173), .A3(n171), .A4(n170), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U208 ( .A1(n2), .A2(i_data_bus[85]), .B1(n273), .B2(
        i_data_bus[53]), .ZN(n180) );
  AOI22D1BWP30P140LVT U209 ( .A1(n4), .A2(i_data_bus[117]), .B1(n274), .B2(
        i_data_bus[149]), .ZN(n179) );
  INVD1BWP30P140LVT U210 ( .I(i_data_bus[213]), .ZN(n175) );
  INVD1BWP30P140LVT U211 ( .I(i_data_bus[181]), .ZN(n174) );
  OAI22D1BWP30P140LVT U212 ( .A1(n277), .A2(n175), .B1(n215), .B2(n174), .ZN(
        n176) );
  ND2D1BWP30P140LVT U213 ( .A1(n279), .A2(i_data_bus[21]), .ZN(n177) );
  ND4D1BWP30P140LVT U214 ( .A1(n179), .A2(n180), .A3(n178), .A4(n177), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U215 ( .A1(n2), .A2(i_data_bus[84]), .B1(n273), .B2(
        i_data_bus[52]), .ZN(n187) );
  AOI22D1BWP30P140LVT U216 ( .A1(n4), .A2(i_data_bus[116]), .B1(n274), .B2(
        i_data_bus[148]), .ZN(n186) );
  INVD1BWP30P140LVT U217 ( .I(i_data_bus[212]), .ZN(n182) );
  INVD1BWP30P140LVT U218 ( .I(i_data_bus[180]), .ZN(n181) );
  OAI22D1BWP30P140LVT U219 ( .A1(n277), .A2(n182), .B1(n189), .B2(n181), .ZN(
        n183) );
  AOI21D1BWP30P140LVT U220 ( .A1(n1), .A2(i_data_bus[244]), .B(n183), .ZN(n185) );
  ND2D1BWP30P140LVT U221 ( .A1(n279), .A2(i_data_bus[20]), .ZN(n184) );
  ND4D1BWP30P140LVT U222 ( .A1(n186), .A2(n187), .A3(n185), .A4(n184), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U223 ( .A1(n2), .A2(i_data_bus[83]), .B1(n273), .B2(
        i_data_bus[51]), .ZN(n195) );
  AOI22D1BWP30P140LVT U224 ( .A1(n4), .A2(i_data_bus[115]), .B1(n274), .B2(
        i_data_bus[147]), .ZN(n194) );
  INVD1BWP30P140LVT U225 ( .I(i_data_bus[211]), .ZN(n190) );
  INVD1BWP30P140LVT U226 ( .I(i_data_bus[179]), .ZN(n188) );
  OAI22D1BWP30P140LVT U227 ( .A1(n277), .A2(n190), .B1(n189), .B2(n188), .ZN(
        n191) );
  AOI21D1BWP30P140LVT U228 ( .A1(n1), .A2(i_data_bus[243]), .B(n191), .ZN(n193) );
  ND2D1BWP30P140LVT U229 ( .A1(n252), .A2(i_data_bus[19]), .ZN(n192) );
  ND4D1BWP30P140LVT U230 ( .A1(n194), .A2(n195), .A3(n193), .A4(n192), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U231 ( .A1(n2), .A2(i_data_bus[82]), .B1(n273), .B2(
        i_data_bus[50]), .ZN(n201) );
  AOI22D1BWP30P140LVT U232 ( .A1(n4), .A2(i_data_bus[114]), .B1(n274), .B2(
        i_data_bus[146]), .ZN(n200) );
  INVD1BWP30P140LVT U233 ( .I(i_data_bus[178]), .ZN(n196) );
  MOAI22D1BWP30P140LVT U234 ( .A1(n215), .A2(n196), .B1(n242), .B2(
        i_data_bus[210]), .ZN(n197) );
  AOI21D1BWP30P140LVT U235 ( .A1(n1), .A2(i_data_bus[242]), .B(n197), .ZN(n199) );
  ND2D1BWP30P140LVT U236 ( .A1(n252), .A2(i_data_bus[18]), .ZN(n198) );
  ND4D1BWP30P140LVT U237 ( .A1(n200), .A2(n201), .A3(n199), .A4(n198), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U238 ( .A1(n2), .A2(i_data_bus[81]), .B1(n273), .B2(
        i_data_bus[49]), .ZN(n207) );
  AOI22D1BWP30P140LVT U239 ( .A1(n4), .A2(i_data_bus[113]), .B1(n274), .B2(
        i_data_bus[145]), .ZN(n206) );
  INVD1BWP30P140LVT U240 ( .I(i_data_bus[177]), .ZN(n202) );
  MOAI22D1BWP30P140LVT U241 ( .A1(n215), .A2(n202), .B1(n242), .B2(
        i_data_bus[209]), .ZN(n203) );
  AOI21D1BWP30P140LVT U242 ( .A1(n1), .A2(i_data_bus[241]), .B(n203), .ZN(n205) );
  ND2D1BWP30P140LVT U243 ( .A1(n230), .A2(i_data_bus[17]), .ZN(n204) );
  ND4D1BWP30P140LVT U244 ( .A1(n206), .A2(n207), .A3(n205), .A4(n204), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U245 ( .A1(n2), .A2(i_data_bus[80]), .B1(n273), .B2(
        i_data_bus[48]), .ZN(n213) );
  AOI22D1BWP30P140LVT U246 ( .A1(n4), .A2(i_data_bus[112]), .B1(n274), .B2(
        i_data_bus[144]), .ZN(n212) );
  INVD1BWP30P140LVT U247 ( .I(i_data_bus[176]), .ZN(n208) );
  MOAI22D1BWP30P140LVT U248 ( .A1(n215), .A2(n208), .B1(n242), .B2(
        i_data_bus[208]), .ZN(n209) );
  AOI21D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[240]), .B(n209), .ZN(n211) );
  ND2D1BWP30P140LVT U250 ( .A1(n230), .A2(i_data_bus[16]), .ZN(n210) );
  ND4D1BWP30P140LVT U251 ( .A1(n212), .A2(n213), .A3(n211), .A4(n210), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U252 ( .A1(n2), .A2(i_data_bus[79]), .B1(n273), .B2(
        i_data_bus[47]), .ZN(n221) );
  AOI22D1BWP30P140LVT U253 ( .A1(n4), .A2(i_data_bus[111]), .B1(n274), .B2(
        i_data_bus[143]), .ZN(n220) );
  INVD1BWP30P140LVT U254 ( .I(i_data_bus[175]), .ZN(n216) );
  OAI21D1BWP30P140LVT U255 ( .A1(n216), .A2(n215), .B(n214), .ZN(n217) );
  AOI21D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[239]), .B(n217), .ZN(n219) );
  ND2D1BWP30P140LVT U257 ( .A1(n252), .A2(i_data_bus[15]), .ZN(n218) );
  ND4D1BWP30P140LVT U258 ( .A1(n221), .A2(n220), .A3(n219), .A4(n218), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U259 ( .A1(n2), .A2(i_data_bus[69]), .B1(n273), .B2(
        i_data_bus[37]), .ZN(n227) );
  AOI22D1BWP30P140LVT U260 ( .A1(n4), .A2(i_data_bus[101]), .B1(n257), .B2(
        i_data_bus[133]), .ZN(n226) );
  INVD1BWP30P140LVT U261 ( .I(i_data_bus[165]), .ZN(n222) );
  MOAI22D1BWP30P140LVT U262 ( .A1(n215), .A2(n222), .B1(n242), .B2(
        i_data_bus[197]), .ZN(n223) );
  AOI21D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[229]), .B(n223), .ZN(n225) );
  ND2D1BWP30P140LVT U264 ( .A1(n279), .A2(i_data_bus[5]), .ZN(n224) );
  ND4D1BWP30P140LVT U265 ( .A1(n227), .A2(n226), .A3(n225), .A4(n224), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U266 ( .A1(n2), .A2(i_data_bus[68]), .B1(n273), .B2(
        i_data_bus[36]), .ZN(n234) );
  AOI22D1BWP30P140LVT U267 ( .A1(n4), .A2(i_data_bus[100]), .B1(n257), .B2(
        i_data_bus[132]), .ZN(n233) );
  INVD1BWP30P140LVT U268 ( .I(i_data_bus[164]), .ZN(n228) );
  MOAI22D1BWP30P140LVT U269 ( .A1(n215), .A2(n228), .B1(n242), .B2(
        i_data_bus[196]), .ZN(n229) );
  AOI21D1BWP30P140LVT U270 ( .A1(n1), .A2(i_data_bus[228]), .B(n229), .ZN(n232) );
  ND2D1BWP30P140LVT U271 ( .A1(n230), .A2(i_data_bus[4]), .ZN(n231) );
  ND4D1BWP30P140LVT U272 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U273 ( .A1(n2), .A2(i_data_bus[67]), .B1(n273), .B2(
        i_data_bus[35]), .ZN(n241) );
  AOI22D1BWP30P140LVT U274 ( .A1(n4), .A2(i_data_bus[99]), .B1(n257), .B2(
        i_data_bus[131]), .ZN(n240) );
  INVD1BWP30P140LVT U275 ( .I(i_data_bus[163]), .ZN(n236) );
  OAI21D1BWP30P140LVT U276 ( .A1(n215), .A2(n236), .B(n235), .ZN(n237) );
  AOI21D1BWP30P140LVT U277 ( .A1(n1), .A2(i_data_bus[227]), .B(n237), .ZN(n239) );
  ND2D1BWP30P140LVT U278 ( .A1(n279), .A2(i_data_bus[3]), .ZN(n238) );
  ND4D1BWP30P140LVT U279 ( .A1(n241), .A2(n240), .A3(n239), .A4(n238), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U280 ( .A1(n2), .A2(i_data_bus[66]), .B1(n273), .B2(
        i_data_bus[34]), .ZN(n249) );
  AOI22D1BWP30P140LVT U281 ( .A1(n4), .A2(i_data_bus[98]), .B1(n257), .B2(
        i_data_bus[130]), .ZN(n248) );
  INVD1BWP30P140LVT U282 ( .I(i_data_bus[162]), .ZN(n244) );
  OAI21D1BWP30P140LVT U283 ( .A1(n215), .A2(n244), .B(n243), .ZN(n245) );
  AOI21D1BWP30P140LVT U284 ( .A1(n1), .A2(i_data_bus[226]), .B(n245), .ZN(n247) );
  ND2D1BWP30P140LVT U285 ( .A1(n252), .A2(i_data_bus[2]), .ZN(n246) );
  ND4D1BWP30P140LVT U286 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U287 ( .A1(n2), .A2(i_data_bus[64]), .B1(n273), .B2(
        i_data_bus[32]), .ZN(n256) );
  AOI22D1BWP30P140LVT U288 ( .A1(n4), .A2(i_data_bus[96]), .B1(n257), .B2(
        i_data_bus[128]), .ZN(n255) );
  INR2D1BWP30P140LVT U289 ( .A1(i_data_bus[192]), .B1(n277), .ZN(n251) );
  INR2D1BWP30P140LVT U290 ( .A1(i_data_bus[160]), .B1(n215), .ZN(n250) );
  AOI211D1BWP30P140LVT U291 ( .A1(i_data_bus[224]), .A2(n1), .B(n251), .C(n250), .ZN(n254) );
  ND2D1BWP30P140LVT U292 ( .A1(n252), .A2(i_data_bus[0]), .ZN(n253) );
  ND4D1BWP30P140LVT U293 ( .A1(n256), .A2(n255), .A3(n254), .A4(n253), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U294 ( .A1(n2), .A2(i_data_bus[65]), .B1(n273), .B2(
        i_data_bus[33]), .ZN(n265) );
  AOI22D1BWP30P140LVT U295 ( .A1(n4), .A2(i_data_bus[97]), .B1(n257), .B2(
        i_data_bus[129]), .ZN(n264) );
  INVD1BWP30P140LVT U296 ( .I(i_data_bus[161]), .ZN(n260) );
  INVD1BWP30P140LVT U297 ( .I(i_data_bus[193]), .ZN(n258) );
  OAI22D1BWP30P140LVT U298 ( .A1(n215), .A2(n260), .B1(n259), .B2(n258), .ZN(
        n261) );
  AOI21D1BWP30P140LVT U299 ( .A1(n1), .A2(i_data_bus[225]), .B(n261), .ZN(n263) );
  ND2D1BWP30P140LVT U300 ( .A1(n279), .A2(i_data_bus[1]), .ZN(n262) );
  ND4D1BWP30P140LVT U301 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U302 ( .A1(n2), .A2(i_data_bus[78]), .B1(n273), .B2(
        i_data_bus[46]), .ZN(n272) );
  AOI22D1BWP30P140LVT U303 ( .A1(n4), .A2(i_data_bus[110]), .B1(n274), .B2(
        i_data_bus[142]), .ZN(n271) );
  INVD1BWP30P140LVT U304 ( .I(i_data_bus[206]), .ZN(n267) );
  INVD1BWP30P140LVT U305 ( .I(i_data_bus[174]), .ZN(n266) );
  OAI22D1BWP30P140LVT U306 ( .A1(n277), .A2(n267), .B1(n215), .B2(n266), .ZN(
        n268) );
  AOI21D1BWP30P140LVT U307 ( .A1(n1), .A2(i_data_bus[238]), .B(n268), .ZN(n270) );
  ND2D1BWP30P140LVT U308 ( .A1(n279), .A2(i_data_bus[14]), .ZN(n269) );
  ND4D1BWP30P140LVT U309 ( .A1(n271), .A2(n272), .A3(n270), .A4(n269), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U310 ( .A1(n2), .A2(i_data_bus[77]), .B1(n273), .B2(
        i_data_bus[45]), .ZN(n283) );
  AOI22D1BWP30P140LVT U311 ( .A1(n4), .A2(i_data_bus[109]), .B1(n274), .B2(
        i_data_bus[141]), .ZN(n282) );
  INVD1BWP30P140LVT U312 ( .I(i_data_bus[205]), .ZN(n276) );
  INVD1BWP30P140LVT U313 ( .I(i_data_bus[173]), .ZN(n275) );
  OAI22D1BWP30P140LVT U314 ( .A1(n277), .A2(n276), .B1(n215), .B2(n275), .ZN(
        n278) );
  AOI21D1BWP30P140LVT U315 ( .A1(n1), .A2(i_data_bus[237]), .B(n278), .ZN(n281) );
  ND2D1BWP30P140LVT U316 ( .A1(n279), .A2(i_data_bus[13]), .ZN(n280) );
  ND4D1BWP30P140LVT U317 ( .A1(n282), .A2(n283), .A3(n281), .A4(n280), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_13 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n171), .ZN(n274) );
  INVD3BWP30P140LVT U4 ( .I(n173), .ZN(n277) );
  NR2D1BWP30P140LVT U5 ( .A1(n47), .A2(n43), .ZN(n44) );
  CKND2D3BWP30P140LVT U6 ( .A1(n25), .A2(n28), .ZN(n172) );
  NR2OPTPAD1BWP30P140LVT U7 ( .A1(n22), .A2(i_cmd[5]), .ZN(n32) );
  AN2D2BWP30P140LVT U8 ( .A1(n29), .A2(n28), .Z(n1) );
  INVD4BWP30P140LVT U9 ( .I(n266), .ZN(n2) );
  INVD2BWP30P140LVT U10 ( .I(n172), .ZN(n3) );
  NR2OPTPAD2BWP30P140LVT U11 ( .A1(n19), .A2(n18), .ZN(n28) );
  CKND2D2BWP30P140LVT U12 ( .A1(n5), .A2(n27), .ZN(n22) );
  INVD2BWP30P140LVT U13 ( .I(n171), .ZN(n257) );
  INVD2BWP30P140LVT U14 ( .I(n168), .ZN(n256) );
  INVD2BWP30P140LVT U15 ( .I(n40), .ZN(n171) );
  NR2D1BWP30P140LVT U16 ( .A1(n31), .A2(i_cmd[4]), .ZN(n33) );
  AOI22D1BWP30P140LVT U17 ( .A1(n258), .A2(i_data_bus[122]), .B1(n274), .B2(
        i_data_bus[154]), .ZN(n92) );
  ND2OPTIBD2BWP30P140LVT U18 ( .A1(n15), .A2(n14), .ZN(n19) );
  INR2D4BWP30P140LVT U19 ( .A1(n48), .B1(n47), .ZN(n169) );
  OR2D1BWP30P140LVT U20 ( .A1(n47), .A2(n36), .Z(n170) );
  INVD1BWP30P140LVT U21 ( .I(n11), .ZN(n177) );
  INVD1BWP30P140LVT U22 ( .I(i_cmd[0]), .ZN(n4) );
  INR3D0BWP30P140LVT U23 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n4), .ZN(n10)
         );
  INVD1BWP30P140LVT U24 ( .I(i_cmd[6]), .ZN(n5) );
  INVD2BWP30P140LVT U25 ( .I(i_cmd[7]), .ZN(n27) );
  INVD1BWP30P140LVT U26 ( .I(rst), .ZN(n6) );
  ND2D1BWP30P140LVT U27 ( .A1(n6), .A2(i_en), .ZN(n30) );
  INVD1BWP30P140LVT U28 ( .I(n30), .ZN(n7) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n32), .A2(n7), .Z(n9) );
  OR2D1BWP30P140LVT U30 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n46) );
  NR2D1BWP30P140LVT U31 ( .A1(n46), .A2(i_cmd[1]), .ZN(n8) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n9), .A2(n8), .ZN(n38) );
  INR2D1BWP30P140LVT U33 ( .A1(n10), .B1(n38), .ZN(n11) );
  NR2D1BWP30P140LVT U34 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n13) );
  CKAN2D1BWP30P140LVT U35 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n12) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n13), .A2(n12), .Z(n20) );
  OR2D4BWP30P140LVT U37 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n35) );
  INVD1BWP30P140LVT U38 ( .I(n35), .ZN(n15) );
  NR2D1BWP30P140LVT U39 ( .A1(i_cmd[0]), .A2(n30), .ZN(n14) );
  INVD1BWP30P140LVT U40 ( .I(i_cmd[3]), .ZN(n17) );
  INVD1BWP30P140LVT U41 ( .I(i_cmd[4]), .ZN(n16) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n17), .A2(n16), .ZN(n18) );
  ND2OPTIBD2BWP30P140LVT U43 ( .A1(n20), .A2(n28), .ZN(n21) );
  INVD3BWP30P140LVT U44 ( .I(n21), .ZN(n266) );
  INVD1BWP30P140LVT U45 ( .I(n22), .ZN(n24) );
  ND2D1BWP30P140LVT U46 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n23) );
  INR2D1BWP30P140LVT U47 ( .A1(n24), .B1(n23), .ZN(n25) );
  INVD1BWP30P140LVT U48 ( .I(i_valid[7]), .ZN(n26) );
  NR4D0BWP30P140LVT U49 ( .A1(n27), .A2(n26), .A3(i_cmd[6]), .A4(i_cmd[5]), 
        .ZN(n29) );
  NR4D0BWP30P140LVT U50 ( .A1(n261), .A2(n266), .A3(n3), .A4(n1), .ZN(n51) );
  OR2D1BWP30P140LVT U51 ( .A1(i_cmd[0]), .A2(n30), .Z(n31) );
  ND2OPTIBD2BWP30P140LVT U52 ( .A1(n33), .A2(n32), .ZN(n47) );
  ND2D1BWP30P140LVT U53 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n34) );
  OR2D1BWP30P140LVT U54 ( .A1(n35), .A2(n34), .Z(n36) );
  ND2OPTIBD1BWP30P140LVT U55 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n37) );
  NR2D1BWP30P140LVT U56 ( .A1(n37), .A2(i_cmd[0]), .ZN(n39) );
  INR2D1BWP30P140LVT U57 ( .A1(n39), .B1(n38), .ZN(n40) );
  NR2D1BWP30P140LVT U58 ( .A1(n275), .A2(n274), .ZN(n50) );
  INVD1BWP30P140LVT U59 ( .I(i_cmd[2]), .ZN(n42) );
  NR2D1BWP30P140LVT U60 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .ZN(n41) );
  IND3D1BWP30P140LVT U61 ( .A1(n42), .B1(i_valid[2]), .B2(n41), .ZN(n43) );
  INVD2BWP30P140LVT U62 ( .I(n44), .ZN(n168) );
  ND2D1BWP30P140LVT U63 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n45) );
  NR2D1BWP30P140LVT U64 ( .A1(n46), .A2(n45), .ZN(n48) );
  INVD1BWP30P140LVT U65 ( .I(n169), .ZN(n49) );
  ND4D1BWP30P140LVT U66 ( .A1(n51), .A2(n50), .A3(n168), .A4(n49), .ZN(N402)
         );
  INVD2BWP30P140LVT U67 ( .I(n168), .ZN(n273) );
  AOI22D1BWP30P140LVT U68 ( .A1(n273), .A2(i_data_bus[95]), .B1(n169), .B2(
        i_data_bus[63]), .ZN(n58) );
  AOI22D1BWP30P140LVT U69 ( .A1(n275), .A2(i_data_bus[127]), .B1(n274), .B2(
        i_data_bus[159]), .ZN(n57) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[223]), .ZN(n53) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[191]), .ZN(n52) );
  OAI22D1BWP30P140LVT U72 ( .A1(n2), .A2(n53), .B1(n172), .B2(n52), .ZN(n54)
         );
  AOI21D1BWP30P140LVT U73 ( .A1(n1), .A2(i_data_bus[255]), .B(n54), .ZN(n56)
         );
  ND2D1BWP30P140LVT U74 ( .A1(n280), .A2(i_data_bus[31]), .ZN(n55) );
  ND4D1BWP30P140LVT U75 ( .A1(n58), .A2(n57), .A3(n56), .A4(n55), .ZN(N400) );
  AOI22D1BWP30P140LVT U76 ( .A1(n273), .A2(i_data_bus[94]), .B1(n169), .B2(
        i_data_bus[62]), .ZN(n65) );
  AOI22D1BWP30P140LVT U77 ( .A1(n258), .A2(i_data_bus[126]), .B1(n274), .B2(
        i_data_bus[158]), .ZN(n64) );
  INVD1BWP30P140LVT U78 ( .I(i_data_bus[222]), .ZN(n60) );
  INVD1BWP30P140LVT U79 ( .I(i_data_bus[190]), .ZN(n59) );
  OAI22D1BWP30P140LVT U80 ( .A1(n2), .A2(n60), .B1(n172), .B2(n59), .ZN(n61)
         );
  AOI21D1BWP30P140LVT U81 ( .A1(n1), .A2(i_data_bus[254]), .B(n61), .ZN(n63)
         );
  ND2D1BWP30P140LVT U82 ( .A1(n261), .A2(i_data_bus[30]), .ZN(n62) );
  ND4D1BWP30P140LVT U83 ( .A1(n65), .A2(n64), .A3(n63), .A4(n62), .ZN(N399) );
  AOI22D1BWP30P140LVT U84 ( .A1(n273), .A2(i_data_bus[93]), .B1(n169), .B2(
        i_data_bus[61]), .ZN(n72) );
  AOI22D1BWP30P140LVT U85 ( .A1(n275), .A2(i_data_bus[125]), .B1(n274), .B2(
        i_data_bus[157]), .ZN(n71) );
  INVD1BWP30P140LVT U86 ( .I(i_data_bus[221]), .ZN(n67) );
  INVD3BWP30P140LVT U87 ( .I(n3), .ZN(n162) );
  INVD1BWP30P140LVT U88 ( .I(i_data_bus[189]), .ZN(n66) );
  OAI22D1BWP30P140LVT U89 ( .A1(n2), .A2(n67), .B1(n162), .B2(n66), .ZN(n68)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n1), .A2(i_data_bus[253]), .B(n68), .ZN(n70)
         );
  ND2D1BWP30P140LVT U91 ( .A1(n280), .A2(i_data_bus[29]), .ZN(n69) );
  ND4D1BWP30P140LVT U92 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(N398) );
  AOI22D1BWP30P140LVT U93 ( .A1(n273), .A2(i_data_bus[92]), .B1(n169), .B2(
        i_data_bus[60]), .ZN(n79) );
  AOI22D1BWP30P140LVT U94 ( .A1(n258), .A2(i_data_bus[124]), .B1(n274), .B2(
        i_data_bus[156]), .ZN(n78) );
  INVD1BWP30P140LVT U95 ( .I(i_data_bus[220]), .ZN(n74) );
  INVD1BWP30P140LVT U96 ( .I(i_data_bus[188]), .ZN(n73) );
  OAI22D1BWP30P140LVT U97 ( .A1(n2), .A2(n74), .B1(n162), .B2(n73), .ZN(n75)
         );
  AOI21D1BWP30P140LVT U98 ( .A1(n1), .A2(i_data_bus[252]), .B(n75), .ZN(n77)
         );
  ND2D1BWP30P140LVT U99 ( .A1(n261), .A2(i_data_bus[28]), .ZN(n76) );
  ND4D1BWP30P140LVT U100 ( .A1(n79), .A2(n78), .A3(n77), .A4(n76), .ZN(N397)
         );
  AOI22D1BWP30P140LVT U101 ( .A1(n273), .A2(i_data_bus[91]), .B1(n169), .B2(
        i_data_bus[59]), .ZN(n86) );
  AOI22D1BWP30P140LVT U102 ( .A1(n275), .A2(i_data_bus[123]), .B1(n274), .B2(
        i_data_bus[155]), .ZN(n85) );
  INVD1BWP30P140LVT U103 ( .I(i_data_bus[219]), .ZN(n81) );
  INVD1BWP30P140LVT U104 ( .I(i_data_bus[187]), .ZN(n80) );
  OAI22D1BWP30P140LVT U105 ( .A1(n2), .A2(n81), .B1(n162), .B2(n80), .ZN(n82)
         );
  AOI21D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[251]), .B(n82), .ZN(n84)
         );
  ND2D1BWP30P140LVT U107 ( .A1(n280), .A2(i_data_bus[27]), .ZN(n83) );
  ND4D1BWP30P140LVT U108 ( .A1(n86), .A2(n85), .A3(n84), .A4(n83), .ZN(N396)
         );
  AOI22D1BWP30P140LVT U109 ( .A1(n273), .A2(i_data_bus[90]), .B1(n169), .B2(
        i_data_bus[58]), .ZN(n93) );
  INVD1BWP30P140LVT U110 ( .I(i_data_bus[218]), .ZN(n88) );
  INVD1BWP30P140LVT U111 ( .I(i_data_bus[186]), .ZN(n87) );
  OAI22D1BWP30P140LVT U112 ( .A1(n2), .A2(n88), .B1(n162), .B2(n87), .ZN(n89)
         );
  AOI21D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[250]), .B(n89), .ZN(n91)
         );
  ND2D1BWP30P140LVT U114 ( .A1(n11), .A2(i_data_bus[26]), .ZN(n90) );
  ND4D1BWP30P140LVT U115 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(N395)
         );
  AOI22D1BWP30P140LVT U116 ( .A1(n273), .A2(i_data_bus[89]), .B1(n169), .B2(
        i_data_bus[57]), .ZN(n100) );
  INVD2BWP30P140LVT U117 ( .I(n170), .ZN(n275) );
  AOI22D1BWP30P140LVT U118 ( .A1(n275), .A2(i_data_bus[121]), .B1(n274), .B2(
        i_data_bus[153]), .ZN(n99) );
  INVD1BWP30P140LVT U119 ( .I(i_data_bus[217]), .ZN(n95) );
  INVD1BWP30P140LVT U120 ( .I(i_data_bus[185]), .ZN(n94) );
  OAI22D1BWP30P140LVT U121 ( .A1(n2), .A2(n95), .B1(n162), .B2(n94), .ZN(n96)
         );
  AOI21D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[249]), .B(n96), .ZN(n98)
         );
  INVD2BWP30P140LVT U123 ( .I(n177), .ZN(n280) );
  ND2D1BWP30P140LVT U124 ( .A1(n280), .A2(i_data_bus[25]), .ZN(n97) );
  ND4D1BWP30P140LVT U125 ( .A1(n100), .A2(n99), .A3(n98), .A4(n97), .ZN(N394)
         );
  AOI22D1BWP30P140LVT U126 ( .A1(n273), .A2(i_data_bus[88]), .B1(n169), .B2(
        i_data_bus[56]), .ZN(n107) );
  AOI22D1BWP30P140LVT U127 ( .A1(n275), .A2(i_data_bus[120]), .B1(n274), .B2(
        i_data_bus[152]), .ZN(n106) );
  INVD1BWP30P140LVT U128 ( .I(i_data_bus[216]), .ZN(n102) );
  INVD1BWP30P140LVT U129 ( .I(i_data_bus[184]), .ZN(n101) );
  OAI22D1BWP30P140LVT U130 ( .A1(n2), .A2(n102), .B1(n162), .B2(n101), .ZN(
        n103) );
  AOI21D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[248]), .B(n103), .ZN(n105) );
  ND2D1BWP30P140LVT U132 ( .A1(n280), .A2(i_data_bus[24]), .ZN(n104) );
  ND4D1BWP30P140LVT U133 ( .A1(n107), .A2(n106), .A3(n105), .A4(n104), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U134 ( .A1(n273), .A2(i_data_bus[87]), .B1(n169), .B2(
        i_data_bus[55]), .ZN(n114) );
  AOI22D1BWP30P140LVT U135 ( .A1(n275), .A2(i_data_bus[119]), .B1(n274), .B2(
        i_data_bus[151]), .ZN(n113) );
  INVD1BWP30P140LVT U136 ( .I(i_data_bus[215]), .ZN(n109) );
  INVD1BWP30P140LVT U137 ( .I(i_data_bus[183]), .ZN(n108) );
  OAI22D1BWP30P140LVT U138 ( .A1(n2), .A2(n109), .B1(n162), .B2(n108), .ZN(
        n110) );
  AOI21D1BWP30P140LVT U139 ( .A1(n1), .A2(i_data_bus[247]), .B(n110), .ZN(n112) );
  ND2D1BWP30P140LVT U140 ( .A1(n280), .A2(i_data_bus[23]), .ZN(n111) );
  ND4D1BWP30P140LVT U141 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U142 ( .A1(n273), .A2(i_data_bus[86]), .B1(n169), .B2(
        i_data_bus[54]), .ZN(n121) );
  AOI22D1BWP30P140LVT U143 ( .A1(n275), .A2(i_data_bus[118]), .B1(n274), .B2(
        i_data_bus[150]), .ZN(n120) );
  INVD1BWP30P140LVT U144 ( .I(i_data_bus[214]), .ZN(n116) );
  INVD1BWP30P140LVT U145 ( .I(i_data_bus[182]), .ZN(n115) );
  OAI22D1BWP30P140LVT U146 ( .A1(n2), .A2(n116), .B1(n162), .B2(n115), .ZN(
        n117) );
  AOI21D1BWP30P140LVT U147 ( .A1(n1), .A2(i_data_bus[246]), .B(n117), .ZN(n119) );
  ND2D1BWP30P140LVT U148 ( .A1(n280), .A2(i_data_bus[22]), .ZN(n118) );
  ND4D1BWP30P140LVT U149 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U150 ( .A1(n273), .A2(i_data_bus[85]), .B1(n169), .B2(
        i_data_bus[53]), .ZN(n128) );
  AOI22D1BWP30P140LVT U151 ( .A1(n275), .A2(i_data_bus[117]), .B1(n274), .B2(
        i_data_bus[149]), .ZN(n127) );
  INVD1BWP30P140LVT U152 ( .I(i_data_bus[213]), .ZN(n123) );
  INVD1BWP30P140LVT U153 ( .I(i_data_bus[181]), .ZN(n122) );
  OAI22D1BWP30P140LVT U154 ( .A1(n2), .A2(n123), .B1(n162), .B2(n122), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U155 ( .A1(n1), .A2(i_data_bus[245]), .B(n124), .ZN(n126) );
  ND2D1BWP30P140LVT U156 ( .A1(n280), .A2(i_data_bus[21]), .ZN(n125) );
  ND4D1BWP30P140LVT U157 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U158 ( .A1(n273), .A2(i_data_bus[84]), .B1(n169), .B2(
        i_data_bus[52]), .ZN(n135) );
  AOI22D1BWP30P140LVT U159 ( .A1(n275), .A2(i_data_bus[116]), .B1(n274), .B2(
        i_data_bus[148]), .ZN(n134) );
  INVD1BWP30P140LVT U160 ( .I(i_data_bus[212]), .ZN(n130) );
  INVD1BWP30P140LVT U161 ( .I(i_data_bus[180]), .ZN(n129) );
  OAI22D1BWP30P140LVT U162 ( .A1(n2), .A2(n130), .B1(n162), .B2(n129), .ZN(
        n131) );
  AOI21D1BWP30P140LVT U163 ( .A1(n1), .A2(i_data_bus[244]), .B(n131), .ZN(n133) );
  ND2D1BWP30P140LVT U164 ( .A1(n280), .A2(i_data_bus[20]), .ZN(n132) );
  ND4D1BWP30P140LVT U165 ( .A1(n135), .A2(n134), .A3(n133), .A4(n132), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U166 ( .A1(n273), .A2(i_data_bus[83]), .B1(n169), .B2(
        i_data_bus[51]), .ZN(n142) );
  AOI22D1BWP30P140LVT U167 ( .A1(n275), .A2(i_data_bus[115]), .B1(n274), .B2(
        i_data_bus[147]), .ZN(n141) );
  INVD1BWP30P140LVT U168 ( .I(i_data_bus[211]), .ZN(n137) );
  INVD1BWP30P140LVT U169 ( .I(i_data_bus[179]), .ZN(n136) );
  OAI22D1BWP30P140LVT U170 ( .A1(n2), .A2(n137), .B1(n162), .B2(n136), .ZN(
        n138) );
  AOI21D1BWP30P140LVT U171 ( .A1(n1), .A2(i_data_bus[243]), .B(n138), .ZN(n140) );
  ND2D1BWP30P140LVT U172 ( .A1(n280), .A2(i_data_bus[19]), .ZN(n139) );
  ND4D1BWP30P140LVT U173 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U174 ( .A1(n273), .A2(i_data_bus[82]), .B1(n169), .B2(
        i_data_bus[50]), .ZN(n148) );
  AOI22D1BWP30P140LVT U175 ( .A1(n275), .A2(i_data_bus[114]), .B1(n274), .B2(
        i_data_bus[146]), .ZN(n147) );
  INVD1BWP30P140LVT U176 ( .I(i_data_bus[178]), .ZN(n143) );
  MOAI22D1BWP30P140LVT U177 ( .A1(n162), .A2(n143), .B1(n266), .B2(
        i_data_bus[210]), .ZN(n144) );
  AOI21D1BWP30P140LVT U178 ( .A1(n1), .A2(i_data_bus[242]), .B(n144), .ZN(n146) );
  ND2D1BWP30P140LVT U179 ( .A1(n280), .A2(i_data_bus[18]), .ZN(n145) );
  ND4D1BWP30P140LVT U180 ( .A1(n148), .A2(n147), .A3(n146), .A4(n145), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U181 ( .A1(n273), .A2(i_data_bus[81]), .B1(n169), .B2(
        i_data_bus[49]), .ZN(n154) );
  AOI22D1BWP30P140LVT U182 ( .A1(n275), .A2(i_data_bus[113]), .B1(n274), .B2(
        i_data_bus[145]), .ZN(n153) );
  INVD1BWP30P140LVT U183 ( .I(i_data_bus[177]), .ZN(n149) );
  MOAI22D1BWP30P140LVT U184 ( .A1(n162), .A2(n149), .B1(n266), .B2(
        i_data_bus[209]), .ZN(n150) );
  AOI21D1BWP30P140LVT U185 ( .A1(n1), .A2(i_data_bus[241]), .B(n150), .ZN(n152) );
  ND2D1BWP30P140LVT U186 ( .A1(n280), .A2(i_data_bus[17]), .ZN(n151) );
  ND4D1BWP30P140LVT U187 ( .A1(n154), .A2(n153), .A3(n152), .A4(n151), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U188 ( .A1(n273), .A2(i_data_bus[80]), .B1(n169), .B2(
        i_data_bus[48]), .ZN(n160) );
  AOI22D1BWP30P140LVT U189 ( .A1(n275), .A2(i_data_bus[112]), .B1(n274), .B2(
        i_data_bus[144]), .ZN(n159) );
  INVD1BWP30P140LVT U190 ( .I(i_data_bus[176]), .ZN(n155) );
  MOAI22D1BWP30P140LVT U191 ( .A1(n162), .A2(n155), .B1(n266), .B2(
        i_data_bus[208]), .ZN(n156) );
  AOI21D1BWP30P140LVT U192 ( .A1(n1), .A2(i_data_bus[240]), .B(n156), .ZN(n158) );
  ND2D1BWP30P140LVT U193 ( .A1(n280), .A2(i_data_bus[16]), .ZN(n157) );
  ND4D1BWP30P140LVT U194 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U195 ( .A1(n273), .A2(i_data_bus[79]), .B1(n169), .B2(
        i_data_bus[47]), .ZN(n167) );
  AOI22D1BWP30P140LVT U196 ( .A1(n275), .A2(i_data_bus[111]), .B1(n274), .B2(
        i_data_bus[143]), .ZN(n166) );
  INVD1BWP30P140LVT U197 ( .I(i_data_bus[175]), .ZN(n161) );
  MOAI22D1BWP30P140LVT U198 ( .A1(n162), .A2(n161), .B1(n266), .B2(
        i_data_bus[207]), .ZN(n163) );
  AOI21D1BWP30P140LVT U199 ( .A1(n1), .A2(i_data_bus[239]), .B(n163), .ZN(n165) );
  ND2D1BWP30P140LVT U200 ( .A1(n280), .A2(i_data_bus[15]), .ZN(n164) );
  ND4D1BWP30P140LVT U201 ( .A1(n167), .A2(n166), .A3(n165), .A4(n164), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U202 ( .A1(n256), .A2(i_data_bus[76]), .B1(n169), .B2(
        i_data_bus[44]), .ZN(n181) );
  INVD2BWP30P140LVT U203 ( .I(n170), .ZN(n258) );
  AOI22D1BWP30P140LVT U204 ( .A1(n258), .A2(i_data_bus[108]), .B1(n257), .B2(
        i_data_bus[140]), .ZN(n180) );
  INVD1BWP30P140LVT U205 ( .I(i_data_bus[204]), .ZN(n175) );
  INVD1BWP30P140LVT U206 ( .I(n172), .ZN(n173) );
  INVD1BWP30P140LVT U207 ( .I(i_data_bus[172]), .ZN(n174) );
  OAI22D1BWP30P140LVT U208 ( .A1(n2), .A2(n175), .B1(n277), .B2(n174), .ZN(
        n176) );
  AOI21D1BWP30P140LVT U209 ( .A1(n1), .A2(i_data_bus[236]), .B(n176), .ZN(n179) );
  INVD2BWP30P140LVT U210 ( .I(n177), .ZN(n261) );
  ND2D1BWP30P140LVT U211 ( .A1(n261), .A2(i_data_bus[12]), .ZN(n178) );
  ND4D1BWP30P140LVT U212 ( .A1(n181), .A2(n180), .A3(n179), .A4(n178), .ZN(
        N381) );
  AOI22D1BWP30P140LVT U213 ( .A1(n256), .A2(i_data_bus[75]), .B1(n169), .B2(
        i_data_bus[43]), .ZN(n188) );
  AOI22D1BWP30P140LVT U214 ( .A1(n258), .A2(i_data_bus[107]), .B1(n257), .B2(
        i_data_bus[139]), .ZN(n187) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[203]), .ZN(n183) );
  INVD1BWP30P140LVT U216 ( .I(i_data_bus[171]), .ZN(n182) );
  OAI22D1BWP30P140LVT U217 ( .A1(n2), .A2(n183), .B1(n277), .B2(n182), .ZN(
        n184) );
  AOI21D1BWP30P140LVT U218 ( .A1(n1), .A2(i_data_bus[235]), .B(n184), .ZN(n186) );
  ND2D1BWP30P140LVT U219 ( .A1(n261), .A2(i_data_bus[11]), .ZN(n185) );
  ND4D1BWP30P140LVT U220 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .ZN(
        N380) );
  AOI22D1BWP30P140LVT U221 ( .A1(n256), .A2(i_data_bus[74]), .B1(n169), .B2(
        i_data_bus[42]), .ZN(n195) );
  AOI22D1BWP30P140LVT U222 ( .A1(n258), .A2(i_data_bus[106]), .B1(n257), .B2(
        i_data_bus[138]), .ZN(n194) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[202]), .ZN(n190) );
  INVD1BWP30P140LVT U224 ( .I(i_data_bus[170]), .ZN(n189) );
  OAI22D1BWP30P140LVT U225 ( .A1(n2), .A2(n190), .B1(n277), .B2(n189), .ZN(
        n191) );
  AOI21D1BWP30P140LVT U226 ( .A1(n1), .A2(i_data_bus[234]), .B(n191), .ZN(n193) );
  ND2D1BWP30P140LVT U227 ( .A1(n261), .A2(i_data_bus[10]), .ZN(n192) );
  ND4D1BWP30P140LVT U228 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U229 ( .A1(n256), .A2(i_data_bus[73]), .B1(n169), .B2(
        i_data_bus[41]), .ZN(n202) );
  AOI22D1BWP30P140LVT U230 ( .A1(n258), .A2(i_data_bus[105]), .B1(n257), .B2(
        i_data_bus[137]), .ZN(n201) );
  INVD1BWP30P140LVT U231 ( .I(i_data_bus[201]), .ZN(n197) );
  INVD1BWP30P140LVT U232 ( .I(i_data_bus[169]), .ZN(n196) );
  OAI22D1BWP30P140LVT U233 ( .A1(n2), .A2(n197), .B1(n277), .B2(n196), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U234 ( .A1(n1), .A2(i_data_bus[233]), .B(n198), .ZN(n200) );
  ND2D1BWP30P140LVT U235 ( .A1(n261), .A2(i_data_bus[9]), .ZN(n199) );
  ND4D1BWP30P140LVT U236 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U237 ( .A1(n256), .A2(i_data_bus[71]), .B1(n169), .B2(
        i_data_bus[39]), .ZN(n209) );
  AOI22D1BWP30P140LVT U238 ( .A1(n258), .A2(i_data_bus[103]), .B1(n257), .B2(
        i_data_bus[135]), .ZN(n208) );
  INVD1BWP30P140LVT U239 ( .I(i_data_bus[199]), .ZN(n204) );
  INVD1BWP30P140LVT U240 ( .I(i_data_bus[167]), .ZN(n203) );
  OAI22D1BWP30P140LVT U241 ( .A1(n2), .A2(n204), .B1(n277), .B2(n203), .ZN(
        n205) );
  AOI21D1BWP30P140LVT U242 ( .A1(n1), .A2(i_data_bus[231]), .B(n205), .ZN(n207) );
  ND2D1BWP30P140LVT U243 ( .A1(n261), .A2(i_data_bus[7]), .ZN(n206) );
  ND4D1BWP30P140LVT U244 ( .A1(n209), .A2(n208), .A3(n207), .A4(n206), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U245 ( .A1(n256), .A2(i_data_bus[70]), .B1(n169), .B2(
        i_data_bus[38]), .ZN(n216) );
  AOI22D1BWP30P140LVT U246 ( .A1(n258), .A2(i_data_bus[102]), .B1(n257), .B2(
        i_data_bus[134]), .ZN(n215) );
  INVD1BWP30P140LVT U247 ( .I(i_data_bus[198]), .ZN(n211) );
  INVD1BWP30P140LVT U248 ( .I(i_data_bus[166]), .ZN(n210) );
  OAI22D1BWP30P140LVT U249 ( .A1(n2), .A2(n211), .B1(n277), .B2(n210), .ZN(
        n212) );
  AOI21D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[230]), .B(n212), .ZN(n214) );
  ND2D1BWP30P140LVT U251 ( .A1(n261), .A2(i_data_bus[6]), .ZN(n213) );
  ND4D1BWP30P140LVT U252 ( .A1(n216), .A2(n215), .A3(n214), .A4(n213), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U253 ( .A1(n256), .A2(i_data_bus[69]), .B1(n169), .B2(
        i_data_bus[37]), .ZN(n223) );
  AOI22D1BWP30P140LVT U254 ( .A1(n258), .A2(i_data_bus[101]), .B1(n257), .B2(
        i_data_bus[133]), .ZN(n222) );
  INVD1BWP30P140LVT U255 ( .I(i_data_bus[197]), .ZN(n218) );
  INVD1BWP30P140LVT U256 ( .I(i_data_bus[165]), .ZN(n217) );
  OAI22D1BWP30P140LVT U257 ( .A1(n2), .A2(n218), .B1(n277), .B2(n217), .ZN(
        n219) );
  AOI21D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[229]), .B(n219), .ZN(n221) );
  ND2D1BWP30P140LVT U259 ( .A1(n261), .A2(i_data_bus[5]), .ZN(n220) );
  ND4D1BWP30P140LVT U260 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U261 ( .A1(n256), .A2(i_data_bus[72]), .B1(n169), .B2(
        i_data_bus[40]), .ZN(n230) );
  AOI22D1BWP30P140LVT U262 ( .A1(n258), .A2(i_data_bus[104]), .B1(n257), .B2(
        i_data_bus[136]), .ZN(n229) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[168]), .ZN(n225) );
  INVD1BWP30P140LVT U264 ( .I(i_data_bus[200]), .ZN(n224) );
  OAI22D1BWP30P140LVT U265 ( .A1(n277), .A2(n225), .B1(n2), .B2(n224), .ZN(
        n226) );
  AOI21OPTREPBD1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[232]), .B(n226), 
        .ZN(n228) );
  ND2D1BWP30P140LVT U267 ( .A1(n261), .A2(i_data_bus[8]), .ZN(n227) );
  ND4D1BWP30P140LVT U268 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U269 ( .A1(n256), .A2(i_data_bus[64]), .B1(n169), .B2(
        i_data_bus[32]), .ZN(n236) );
  AOI22D1BWP30P140LVT U270 ( .A1(n258), .A2(i_data_bus[96]), .B1(n257), .B2(
        i_data_bus[128]), .ZN(n235) );
  INR2D1BWP30P140LVT U271 ( .A1(i_data_bus[192]), .B1(n2), .ZN(n232) );
  INR2D1BWP30P140LVT U272 ( .A1(i_data_bus[160]), .B1(n277), .ZN(n231) );
  AOI211D1BWP30P140LVT U273 ( .A1(i_data_bus[224]), .A2(n1), .B(n232), .C(n231), .ZN(n234) );
  ND2D1BWP30P140LVT U274 ( .A1(n261), .A2(i_data_bus[0]), .ZN(n233) );
  ND4D1BWP30P140LVT U275 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U276 ( .A1(n256), .A2(i_data_bus[68]), .B1(n169), .B2(
        i_data_bus[36]), .ZN(n243) );
  AOI22D1BWP30P140LVT U277 ( .A1(n258), .A2(i_data_bus[100]), .B1(n257), .B2(
        i_data_bus[132]), .ZN(n242) );
  INVD1BWP30P140LVT U278 ( .I(i_data_bus[196]), .ZN(n238) );
  INVD1BWP30P140LVT U279 ( .I(i_data_bus[164]), .ZN(n237) );
  OAI22D1BWP30P140LVT U280 ( .A1(n2), .A2(n238), .B1(n277), .B2(n237), .ZN(
        n239) );
  AOI21D1BWP30P140LVT U281 ( .A1(n1), .A2(i_data_bus[228]), .B(n239), .ZN(n241) );
  ND2D1BWP30P140LVT U282 ( .A1(n261), .A2(i_data_bus[4]), .ZN(n240) );
  ND4D1BWP30P140LVT U283 ( .A1(n243), .A2(n242), .A3(n241), .A4(n240), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U284 ( .A1(n256), .A2(i_data_bus[67]), .B1(n169), .B2(
        i_data_bus[35]), .ZN(n249) );
  AOI22D1BWP30P140LVT U285 ( .A1(n258), .A2(i_data_bus[99]), .B1(n257), .B2(
        i_data_bus[131]), .ZN(n248) );
  INVD1BWP30P140LVT U286 ( .I(i_data_bus[163]), .ZN(n244) );
  MOAI22D1BWP30P140LVT U287 ( .A1(n277), .A2(n244), .B1(n266), .B2(
        i_data_bus[195]), .ZN(n245) );
  AOI21D1BWP30P140LVT U288 ( .A1(n1), .A2(i_data_bus[227]), .B(n245), .ZN(n247) );
  ND2D1BWP30P140LVT U289 ( .A1(n261), .A2(i_data_bus[3]), .ZN(n246) );
  ND4D1BWP30P140LVT U290 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U291 ( .A1(n256), .A2(i_data_bus[66]), .B1(n169), .B2(
        i_data_bus[34]), .ZN(n255) );
  AOI22D1BWP30P140LVT U292 ( .A1(n258), .A2(i_data_bus[98]), .B1(n257), .B2(
        i_data_bus[130]), .ZN(n254) );
  INVD1BWP30P140LVT U293 ( .I(i_data_bus[162]), .ZN(n250) );
  MOAI22D1BWP30P140LVT U294 ( .A1(n277), .A2(n250), .B1(n266), .B2(
        i_data_bus[194]), .ZN(n251) );
  AOI21D1BWP30P140LVT U295 ( .A1(n1), .A2(i_data_bus[226]), .B(n251), .ZN(n253) );
  ND2D1BWP30P140LVT U296 ( .A1(n261), .A2(i_data_bus[2]), .ZN(n252) );
  ND4D1BWP30P140LVT U297 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U298 ( .A1(n256), .A2(i_data_bus[65]), .B1(n169), .B2(
        i_data_bus[33]), .ZN(n265) );
  AOI22D1BWP30P140LVT U299 ( .A1(n258), .A2(i_data_bus[97]), .B1(n257), .B2(
        i_data_bus[129]), .ZN(n264) );
  INVD1BWP30P140LVT U300 ( .I(i_data_bus[161]), .ZN(n259) );
  MOAI22D1BWP30P140LVT U301 ( .A1(n277), .A2(n259), .B1(n266), .B2(
        i_data_bus[193]), .ZN(n260) );
  AOI21D1BWP30P140LVT U302 ( .A1(n1), .A2(i_data_bus[225]), .B(n260), .ZN(n263) );
  ND2D1BWP30P140LVT U303 ( .A1(n261), .A2(i_data_bus[1]), .ZN(n262) );
  ND4D1BWP30P140LVT U304 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U305 ( .A1(n273), .A2(i_data_bus[78]), .B1(n169), .B2(
        i_data_bus[46]), .ZN(n272) );
  AOI22D1BWP30P140LVT U306 ( .A1(n275), .A2(i_data_bus[110]), .B1(n274), .B2(
        i_data_bus[142]), .ZN(n271) );
  INVD1BWP30P140LVT U307 ( .I(i_data_bus[174]), .ZN(n267) );
  MOAI22D1BWP30P140LVT U308 ( .A1(n277), .A2(n267), .B1(n266), .B2(
        i_data_bus[206]), .ZN(n268) );
  AOI21D1BWP30P140LVT U309 ( .A1(n1), .A2(i_data_bus[238]), .B(n268), .ZN(n270) );
  ND2D1BWP30P140LVT U310 ( .A1(n280), .A2(i_data_bus[14]), .ZN(n269) );
  ND4D1BWP30P140LVT U311 ( .A1(n272), .A2(n271), .A3(n270), .A4(n269), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U312 ( .A1(n273), .A2(i_data_bus[77]), .B1(n169), .B2(
        i_data_bus[45]), .ZN(n284) );
  AOI22D1BWP30P140LVT U313 ( .A1(n275), .A2(i_data_bus[109]), .B1(n274), .B2(
        i_data_bus[141]), .ZN(n283) );
  INVD1BWP30P140LVT U314 ( .I(i_data_bus[205]), .ZN(n278) );
  INVD1BWP30P140LVT U315 ( .I(i_data_bus[173]), .ZN(n276) );
  OAI22D1BWP30P140LVT U316 ( .A1(n2), .A2(n278), .B1(n277), .B2(n276), .ZN(
        n279) );
  AOI21D1BWP30P140LVT U317 ( .A1(n1), .A2(i_data_bus[237]), .B(n279), .ZN(n282) );
  ND2D1BWP30P140LVT U318 ( .A1(n280), .A2(i_data_bus[13]), .ZN(n281) );
  ND4D1BWP30P140LVT U319 ( .A1(n284), .A2(n283), .A3(n282), .A4(n281), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_14 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n172), .ZN(n276) );
  INR2D4BWP30P140LVT U4 ( .A1(n24), .B1(n19), .ZN(n266) );
  CKBD1BWP30P140LVT U5 ( .I(n42), .Z(n45) );
  CKND2D3BWP30P140LVT U6 ( .A1(n22), .A2(n24), .ZN(n173) );
  NR2OPTPAD1BWP30P140LVT U7 ( .A1(n21), .A2(i_cmd[5]), .ZN(n31) );
  INVD1BWP30P140LVT U8 ( .I(n27), .ZN(n77) );
  INVD4BWP30P140LVT U9 ( .I(n4), .ZN(n163) );
  INVD2BWP30P140LVT U10 ( .I(n170), .ZN(n1) );
  INVD4BWP30P140LVT U11 ( .I(n171), .ZN(n2) );
  INVD8BWP30P140LVT U12 ( .I(n266), .ZN(n3) );
  INVD2BWP30P140LVT U13 ( .I(n173), .ZN(n4) );
  INVD2BWP30P140LVT U14 ( .I(n38), .ZN(n172) );
  INVD2BWP30P140LVT U15 ( .I(n172), .ZN(n258) );
  OR2D4BWP30P140LVT U16 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n21) );
  NR2D1BWP30P140LVT U17 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n18) );
  ND2D1BWP30P140LVT U18 ( .A1(n14), .A2(n13), .ZN(n15) );
  INR2D1BWP30P140LVT U19 ( .A1(n37), .B1(n36), .ZN(n38) );
  INVD1BWP30P140LVT U20 ( .I(n9), .ZN(n178) );
  INVD2BWP30P140LVT U21 ( .I(n1), .ZN(n257) );
  INVD2BWP30P140LVT U22 ( .I(n94), .ZN(n274) );
  OR2D1BWP30P140LVT U23 ( .A1(n42), .A2(n41), .Z(n169) );
  INVD1BWP30P140LVT U24 ( .I(i_cmd[0]), .ZN(n10) );
  INR3D0BWP30P140LVT U25 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n10), .ZN(n8)
         );
  INVD1BWP30P140LVT U26 ( .I(rst), .ZN(n5) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n5), .A2(i_en), .Z(n12) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n31), .A2(n12), .Z(n7) );
  OR2D1BWP30P140LVT U29 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n44) );
  NR2D1BWP30P140LVT U30 ( .A1(n44), .A2(i_cmd[1]), .ZN(n6) );
  ND2OPTIBD2BWP30P140LVT U31 ( .A1(n7), .A2(n6), .ZN(n36) );
  INR2D1BWP30P140LVT U32 ( .A1(n8), .B1(n36), .ZN(n9) );
  INVD1BWP30P140LVT U33 ( .I(n178), .ZN(n89) );
  OR2D4BWP30P140LVT U34 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n33) );
  INVD1BWP30P140LVT U35 ( .I(n33), .ZN(n11) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(n11), .A2(n10), .ZN(n16) );
  INVD1BWP30P140LVT U37 ( .I(i_cmd[3]), .ZN(n14) );
  INVD1BWP30P140LVT U38 ( .I(n12), .ZN(n28) );
  NR2D1BWP30P140LVT U39 ( .A1(i_cmd[4]), .A2(n28), .ZN(n13) );
  NR2D3BWP30P140LVT U40 ( .A1(n16), .A2(n15), .ZN(n24) );
  CKAN2D1BWP30P140LVT U41 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n17) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n18), .A2(n17), .ZN(n19) );
  ND2D1BWP30P140LVT U43 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n20) );
  NR2D1BWP30P140LVT U44 ( .A1(n21), .A2(n20), .ZN(n22) );
  INVD1BWP30P140LVT U45 ( .I(i_cmd[7]), .ZN(n23) );
  INR4D0BWP30P140LVT U46 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n23), .ZN(n26) );
  INVD1BWP30P140LVT U47 ( .I(n24), .ZN(n25) );
  INR2D1BWP30P140LVT U48 ( .A1(n26), .B1(n25), .ZN(n27) );
  INVD2BWP30P140LVT U49 ( .I(n77), .ZN(n281) );
  NR4D0BWP30P140LVT U50 ( .A1(n89), .A2(n266), .A3(n4), .A4(n281), .ZN(n48) );
  NR2D1BWP30P140LVT U51 ( .A1(i_cmd[0]), .A2(n28), .ZN(n30) );
  INVD1BWP30P140LVT U52 ( .I(i_cmd[4]), .ZN(n29) );
  ND3D2BWP30P140LVT U53 ( .A1(n31), .A2(n30), .A3(n29), .ZN(n42) );
  ND2D1BWP30P140LVT U54 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n32) );
  NR2D1BWP30P140LVT U55 ( .A1(n33), .A2(n32), .ZN(n34) );
  IND2D2BWP30P140LVT U56 ( .A1(n45), .B1(n34), .ZN(n171) );
  ND2D1BWP30P140LVT U57 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n35) );
  NR2D1BWP30P140LVT U58 ( .A1(n35), .A2(i_cmd[0]), .ZN(n37) );
  NR2D1BWP30P140LVT U59 ( .A1(n2), .A2(n276), .ZN(n47) );
  INVD1BWP30P140LVT U60 ( .I(i_cmd[2]), .ZN(n40) );
  NR2D1BWP30P140LVT U61 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .ZN(n39) );
  IND3D1BWP30P140LVT U62 ( .A1(n40), .B1(n39), .B2(i_valid[2]), .ZN(n41) );
  INVD2BWP30P140LVT U63 ( .I(n169), .ZN(n275) );
  ND2D1BWP30P140LVT U64 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n43) );
  NR2D1BWP30P140LVT U65 ( .A1(n44), .A2(n43), .ZN(n46) );
  INR2D2BWP30P140LVT U66 ( .A1(n46), .B1(n45), .ZN(n170) );
  ND4D1BWP30P140LVT U67 ( .A1(n48), .A2(n47), .A3(n169), .A4(n1), .ZN(N402) );
  INVD1BWP30P140LVT U68 ( .I(n1), .ZN(n85) );
  AOI22D1BWP30P140LVT U69 ( .A1(n275), .A2(i_data_bus[95]), .B1(n85), .B2(
        i_data_bus[63]), .ZN(n55) );
  AOI22D1BWP30P140LVT U70 ( .A1(n2), .A2(i_data_bus[127]), .B1(n276), .B2(
        i_data_bus[159]), .ZN(n54) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[223]), .ZN(n50) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[191]), .ZN(n49) );
  OAI22D1BWP30P140LVT U73 ( .A1(n3), .A2(n50), .B1(n173), .B2(n49), .ZN(n51)
         );
  AOI21D1BWP30P140LVT U74 ( .A1(n281), .A2(i_data_bus[255]), .B(n51), .ZN(n53)
         );
  ND2D1BWP30P140LVT U75 ( .A1(n89), .A2(i_data_bus[31]), .ZN(n52) );
  ND4D1BWP30P140LVT U76 ( .A1(n55), .A2(n54), .A3(n53), .A4(n52), .ZN(N400) );
  AOI22D1BWP30P140LVT U77 ( .A1(n275), .A2(i_data_bus[94]), .B1(n85), .B2(
        i_data_bus[62]), .ZN(n62) );
  AOI22D1BWP30P140LVT U78 ( .A1(n2), .A2(i_data_bus[126]), .B1(n276), .B2(
        i_data_bus[158]), .ZN(n61) );
  INVD1BWP30P140LVT U79 ( .I(i_data_bus[222]), .ZN(n57) );
  INVD1BWP30P140LVT U80 ( .I(i_data_bus[190]), .ZN(n56) );
  OAI22D1BWP30P140LVT U81 ( .A1(n3), .A2(n57), .B1(n173), .B2(n56), .ZN(n58)
         );
  AOI21D1BWP30P140LVT U82 ( .A1(n269), .A2(i_data_bus[254]), .B(n58), .ZN(n60)
         );
  ND2D1BWP30P140LVT U83 ( .A1(n89), .A2(i_data_bus[30]), .ZN(n59) );
  ND4D1BWP30P140LVT U84 ( .A1(n62), .A2(n61), .A3(n60), .A4(n59), .ZN(N399) );
  AOI22D1BWP30P140LVT U85 ( .A1(n275), .A2(i_data_bus[93]), .B1(n85), .B2(
        i_data_bus[61]), .ZN(n69) );
  AOI22D1BWP30P140LVT U86 ( .A1(n2), .A2(i_data_bus[125]), .B1(n276), .B2(
        i_data_bus[157]), .ZN(n68) );
  INVD1BWP30P140LVT U87 ( .I(i_data_bus[221]), .ZN(n64) );
  INVD1BWP30P140LVT U88 ( .I(i_data_bus[189]), .ZN(n63) );
  OAI22D1BWP30P140LVT U89 ( .A1(n3), .A2(n64), .B1(n163), .B2(n63), .ZN(n65)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n269), .A2(i_data_bus[253]), .B(n65), .ZN(n67)
         );
  ND2D1BWP30P140LVT U91 ( .A1(n89), .A2(i_data_bus[29]), .ZN(n66) );
  ND4D1BWP30P140LVT U92 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(N398) );
  AOI22D1BWP30P140LVT U93 ( .A1(n275), .A2(i_data_bus[92]), .B1(n85), .B2(
        i_data_bus[60]), .ZN(n76) );
  AOI22D1BWP30P140LVT U94 ( .A1(n2), .A2(i_data_bus[124]), .B1(n276), .B2(
        i_data_bus[156]), .ZN(n75) );
  INVD1BWP30P140LVT U95 ( .I(i_data_bus[220]), .ZN(n71) );
  INVD1BWP30P140LVT U96 ( .I(i_data_bus[188]), .ZN(n70) );
  OAI22D1BWP30P140LVT U97 ( .A1(n3), .A2(n71), .B1(n163), .B2(n70), .ZN(n72)
         );
  AOI21D1BWP30P140LVT U98 ( .A1(n281), .A2(i_data_bus[252]), .B(n72), .ZN(n74)
         );
  ND2D1BWP30P140LVT U99 ( .A1(n89), .A2(i_data_bus[28]), .ZN(n73) );
  ND4D1BWP30P140LVT U100 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(N397)
         );
  AOI22D1BWP30P140LVT U101 ( .A1(n275), .A2(i_data_bus[91]), .B1(n85), .B2(
        i_data_bus[59]), .ZN(n84) );
  AOI22D1BWP30P140LVT U102 ( .A1(n2), .A2(i_data_bus[123]), .B1(n276), .B2(
        i_data_bus[155]), .ZN(n83) );
  INVD2BWP30P140LVT U103 ( .I(n77), .ZN(n269) );
  INVD1BWP30P140LVT U104 ( .I(i_data_bus[219]), .ZN(n79) );
  INVD1BWP30P140LVT U105 ( .I(i_data_bus[187]), .ZN(n78) );
  OAI22D1BWP30P140LVT U106 ( .A1(n3), .A2(n79), .B1(n163), .B2(n78), .ZN(n80)
         );
  AOI21D1BWP30P140LVT U107 ( .A1(n269), .A2(i_data_bus[251]), .B(n80), .ZN(n82) );
  ND2D1BWP30P140LVT U108 ( .A1(n89), .A2(i_data_bus[27]), .ZN(n81) );
  ND4D1BWP30P140LVT U109 ( .A1(n84), .A2(n83), .A3(n82), .A4(n81), .ZN(N396)
         );
  AOI22D1BWP30P140LVT U110 ( .A1(n275), .A2(i_data_bus[90]), .B1(n85), .B2(
        i_data_bus[58]), .ZN(n93) );
  AOI22D1BWP30P140LVT U111 ( .A1(n2), .A2(i_data_bus[122]), .B1(n276), .B2(
        i_data_bus[154]), .ZN(n92) );
  INVD1BWP30P140LVT U112 ( .I(i_data_bus[218]), .ZN(n87) );
  INVD1BWP30P140LVT U113 ( .I(i_data_bus[186]), .ZN(n86) );
  OAI22D1BWP30P140LVT U114 ( .A1(n3), .A2(n87), .B1(n163), .B2(n86), .ZN(n88)
         );
  AOI21D1BWP30P140LVT U115 ( .A1(n269), .A2(i_data_bus[250]), .B(n88), .ZN(n91) );
  ND2D1BWP30P140LVT U116 ( .A1(n89), .A2(i_data_bus[26]), .ZN(n90) );
  ND4D1BWP30P140LVT U117 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(N395)
         );
  INVD1BWP30P140LVT U118 ( .I(n170), .ZN(n94) );
  AOI22D1BWP30P140LVT U119 ( .A1(n275), .A2(i_data_bus[89]), .B1(n274), .B2(
        i_data_bus[57]), .ZN(n101) );
  AOI22D1BWP30P140LVT U120 ( .A1(n2), .A2(i_data_bus[121]), .B1(n276), .B2(
        i_data_bus[153]), .ZN(n100) );
  INVD1BWP30P140LVT U121 ( .I(i_data_bus[217]), .ZN(n96) );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[185]), .ZN(n95) );
  OAI22D1BWP30P140LVT U123 ( .A1(n3), .A2(n96), .B1(n163), .B2(n95), .ZN(n97)
         );
  AOI21D1BWP30P140LVT U124 ( .A1(n269), .A2(i_data_bus[249]), .B(n97), .ZN(n99) );
  INVD2BWP30P140LVT U125 ( .I(n178), .ZN(n282) );
  ND2D1BWP30P140LVT U126 ( .A1(n282), .A2(i_data_bus[25]), .ZN(n98) );
  ND4D1BWP30P140LVT U127 ( .A1(n101), .A2(n100), .A3(n99), .A4(n98), .ZN(N394)
         );
  AOI22D1BWP30P140LVT U128 ( .A1(n275), .A2(i_data_bus[88]), .B1(n274), .B2(
        i_data_bus[56]), .ZN(n108) );
  AOI22D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[120]), .B1(n276), .B2(
        i_data_bus[152]), .ZN(n107) );
  INVD1BWP30P140LVT U130 ( .I(i_data_bus[216]), .ZN(n103) );
  INVD1BWP30P140LVT U131 ( .I(i_data_bus[184]), .ZN(n102) );
  OAI22D1BWP30P140LVT U132 ( .A1(n3), .A2(n103), .B1(n163), .B2(n102), .ZN(
        n104) );
  AOI21D1BWP30P140LVT U133 ( .A1(n269), .A2(i_data_bus[248]), .B(n104), .ZN(
        n106) );
  ND2D1BWP30P140LVT U134 ( .A1(n282), .A2(i_data_bus[24]), .ZN(n105) );
  ND4D1BWP30P140LVT U135 ( .A1(n108), .A2(n107), .A3(n106), .A4(n105), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U136 ( .A1(n275), .A2(i_data_bus[87]), .B1(n274), .B2(
        i_data_bus[55]), .ZN(n115) );
  AOI22D1BWP30P140LVT U137 ( .A1(n2), .A2(i_data_bus[119]), .B1(n276), .B2(
        i_data_bus[151]), .ZN(n114) );
  INVD1BWP30P140LVT U138 ( .I(i_data_bus[215]), .ZN(n110) );
  INVD1BWP30P140LVT U139 ( .I(i_data_bus[183]), .ZN(n109) );
  OAI22D1BWP30P140LVT U140 ( .A1(n3), .A2(n110), .B1(n163), .B2(n109), .ZN(
        n111) );
  AOI21D1BWP30P140LVT U141 ( .A1(n269), .A2(i_data_bus[247]), .B(n111), .ZN(
        n113) );
  ND2D1BWP30P140LVT U142 ( .A1(n282), .A2(i_data_bus[23]), .ZN(n112) );
  ND4D1BWP30P140LVT U143 ( .A1(n115), .A2(n114), .A3(n113), .A4(n112), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U144 ( .A1(n275), .A2(i_data_bus[86]), .B1(n274), .B2(
        i_data_bus[54]), .ZN(n122) );
  AOI22D1BWP30P140LVT U145 ( .A1(n2), .A2(i_data_bus[118]), .B1(n276), .B2(
        i_data_bus[150]), .ZN(n121) );
  INVD1BWP30P140LVT U146 ( .I(i_data_bus[214]), .ZN(n117) );
  INVD1BWP30P140LVT U147 ( .I(i_data_bus[182]), .ZN(n116) );
  OAI22D1BWP30P140LVT U148 ( .A1(n3), .A2(n117), .B1(n163), .B2(n116), .ZN(
        n118) );
  AOI21D1BWP30P140LVT U149 ( .A1(n269), .A2(i_data_bus[246]), .B(n118), .ZN(
        n120) );
  ND2D1BWP30P140LVT U150 ( .A1(n282), .A2(i_data_bus[22]), .ZN(n119) );
  ND4D1BWP30P140LVT U151 ( .A1(n122), .A2(n121), .A3(n120), .A4(n119), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U152 ( .A1(n275), .A2(i_data_bus[85]), .B1(n274), .B2(
        i_data_bus[53]), .ZN(n129) );
  AOI22D1BWP30P140LVT U153 ( .A1(n2), .A2(i_data_bus[117]), .B1(n276), .B2(
        i_data_bus[149]), .ZN(n128) );
  INVD1BWP30P140LVT U154 ( .I(i_data_bus[213]), .ZN(n124) );
  INVD1BWP30P140LVT U155 ( .I(i_data_bus[181]), .ZN(n123) );
  OAI22D1BWP30P140LVT U156 ( .A1(n3), .A2(n124), .B1(n163), .B2(n123), .ZN(
        n125) );
  AOI21D1BWP30P140LVT U157 ( .A1(n269), .A2(i_data_bus[245]), .B(n125), .ZN(
        n127) );
  ND2D1BWP30P140LVT U158 ( .A1(n282), .A2(i_data_bus[21]), .ZN(n126) );
  ND4D1BWP30P140LVT U159 ( .A1(n129), .A2(n128), .A3(n127), .A4(n126), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U160 ( .A1(n275), .A2(i_data_bus[84]), .B1(n274), .B2(
        i_data_bus[52]), .ZN(n136) );
  AOI22D1BWP30P140LVT U161 ( .A1(n2), .A2(i_data_bus[116]), .B1(n276), .B2(
        i_data_bus[148]), .ZN(n135) );
  INVD1BWP30P140LVT U162 ( .I(i_data_bus[212]), .ZN(n131) );
  INVD1BWP30P140LVT U163 ( .I(i_data_bus[180]), .ZN(n130) );
  OAI22D1BWP30P140LVT U164 ( .A1(n3), .A2(n131), .B1(n163), .B2(n130), .ZN(
        n132) );
  AOI21D1BWP30P140LVT U165 ( .A1(n269), .A2(i_data_bus[244]), .B(n132), .ZN(
        n134) );
  ND2D1BWP30P140LVT U166 ( .A1(n282), .A2(i_data_bus[20]), .ZN(n133) );
  ND4D1BWP30P140LVT U167 ( .A1(n136), .A2(n135), .A3(n134), .A4(n133), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U168 ( .A1(n275), .A2(i_data_bus[83]), .B1(n274), .B2(
        i_data_bus[51]), .ZN(n143) );
  AOI22D1BWP30P140LVT U169 ( .A1(n2), .A2(i_data_bus[115]), .B1(n276), .B2(
        i_data_bus[147]), .ZN(n142) );
  INVD1BWP30P140LVT U170 ( .I(i_data_bus[211]), .ZN(n138) );
  INVD1BWP30P140LVT U171 ( .I(i_data_bus[179]), .ZN(n137) );
  OAI22D1BWP30P140LVT U172 ( .A1(n3), .A2(n138), .B1(n163), .B2(n137), .ZN(
        n139) );
  AOI21D1BWP30P140LVT U173 ( .A1(n269), .A2(i_data_bus[243]), .B(n139), .ZN(
        n141) );
  ND2D1BWP30P140LVT U174 ( .A1(n282), .A2(i_data_bus[19]), .ZN(n140) );
  ND4D1BWP30P140LVT U175 ( .A1(n143), .A2(n142), .A3(n141), .A4(n140), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U176 ( .A1(n275), .A2(i_data_bus[82]), .B1(n274), .B2(
        i_data_bus[50]), .ZN(n149) );
  AOI22D1BWP30P140LVT U177 ( .A1(n2), .A2(i_data_bus[114]), .B1(n276), .B2(
        i_data_bus[146]), .ZN(n148) );
  INVD1BWP30P140LVT U178 ( .I(i_data_bus[178]), .ZN(n144) );
  MOAI22D1BWP30P140LVT U179 ( .A1(n163), .A2(n144), .B1(n266), .B2(
        i_data_bus[210]), .ZN(n145) );
  AOI21D1BWP30P140LVT U180 ( .A1(n269), .A2(i_data_bus[242]), .B(n145), .ZN(
        n147) );
  ND2D1BWP30P140LVT U181 ( .A1(n282), .A2(i_data_bus[18]), .ZN(n146) );
  ND4D1BWP30P140LVT U182 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U183 ( .A1(n275), .A2(i_data_bus[81]), .B1(n274), .B2(
        i_data_bus[49]), .ZN(n155) );
  AOI22D1BWP30P140LVT U184 ( .A1(n2), .A2(i_data_bus[113]), .B1(n276), .B2(
        i_data_bus[145]), .ZN(n154) );
  INVD1BWP30P140LVT U185 ( .I(i_data_bus[177]), .ZN(n150) );
  MOAI22D1BWP30P140LVT U186 ( .A1(n163), .A2(n150), .B1(n266), .B2(
        i_data_bus[209]), .ZN(n151) );
  AOI21D1BWP30P140LVT U187 ( .A1(n269), .A2(i_data_bus[241]), .B(n151), .ZN(
        n153) );
  ND2D1BWP30P140LVT U188 ( .A1(n282), .A2(i_data_bus[17]), .ZN(n152) );
  ND4D1BWP30P140LVT U189 ( .A1(n155), .A2(n154), .A3(n153), .A4(n152), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U190 ( .A1(n275), .A2(i_data_bus[80]), .B1(n274), .B2(
        i_data_bus[48]), .ZN(n161) );
  AOI22D1BWP30P140LVT U191 ( .A1(n2), .A2(i_data_bus[112]), .B1(n276), .B2(
        i_data_bus[144]), .ZN(n160) );
  INVD1BWP30P140LVT U192 ( .I(i_data_bus[176]), .ZN(n156) );
  MOAI22D1BWP30P140LVT U193 ( .A1(n163), .A2(n156), .B1(n266), .B2(
        i_data_bus[208]), .ZN(n157) );
  AOI21D1BWP30P140LVT U194 ( .A1(n269), .A2(i_data_bus[240]), .B(n157), .ZN(
        n159) );
  ND2D1BWP30P140LVT U195 ( .A1(n282), .A2(i_data_bus[16]), .ZN(n158) );
  ND4D1BWP30P140LVT U196 ( .A1(n161), .A2(n160), .A3(n159), .A4(n158), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U197 ( .A1(n275), .A2(i_data_bus[79]), .B1(n274), .B2(
        i_data_bus[47]), .ZN(n168) );
  AOI22D1BWP30P140LVT U198 ( .A1(n2), .A2(i_data_bus[111]), .B1(n276), .B2(
        i_data_bus[143]), .ZN(n167) );
  INVD1BWP30P140LVT U199 ( .I(i_data_bus[175]), .ZN(n162) );
  MOAI22D1BWP30P140LVT U200 ( .A1(n163), .A2(n162), .B1(n266), .B2(
        i_data_bus[207]), .ZN(n164) );
  AOI21D1BWP30P140LVT U201 ( .A1(n269), .A2(i_data_bus[239]), .B(n164), .ZN(
        n166) );
  ND2D1BWP30P140LVT U202 ( .A1(n282), .A2(i_data_bus[15]), .ZN(n165) );
  ND4D1BWP30P140LVT U203 ( .A1(n168), .A2(n167), .A3(n166), .A4(n165), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U204 ( .A1(n275), .A2(i_data_bus[72]), .B1(n257), .B2(
        i_data_bus[40]), .ZN(n182) );
  AOI22D1BWP30P140LVT U205 ( .A1(n2), .A2(i_data_bus[104]), .B1(n258), .B2(
        i_data_bus[136]), .ZN(n181) );
  INVD2BWP30P140LVT U206 ( .I(n173), .ZN(n174) );
  INVD3BWP30P140LVT U207 ( .I(n174), .ZN(n278) );
  INVD1BWP30P140LVT U208 ( .I(i_data_bus[168]), .ZN(n176) );
  INVD1BWP30P140LVT U209 ( .I(i_data_bus[200]), .ZN(n175) );
  OAI22D1BWP30P140LVT U210 ( .A1(n278), .A2(n176), .B1(n3), .B2(n175), .ZN(
        n177) );
  AOI21OPTREPBD1BWP30P140LVT U211 ( .A1(n269), .A2(i_data_bus[232]), .B(n177), 
        .ZN(n180) );
  INVD2BWP30P140LVT U212 ( .I(n178), .ZN(n261) );
  ND2D1BWP30P140LVT U213 ( .A1(n261), .A2(i_data_bus[8]), .ZN(n179) );
  ND4D1BWP30P140LVT U214 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U215 ( .A1(n275), .A2(i_data_bus[76]), .B1(n257), .B2(
        i_data_bus[44]), .ZN(n189) );
  AOI22D1BWP30P140LVT U216 ( .A1(n2), .A2(i_data_bus[108]), .B1(n258), .B2(
        i_data_bus[140]), .ZN(n188) );
  INVD1BWP30P140LVT U217 ( .I(i_data_bus[204]), .ZN(n184) );
  INVD1BWP30P140LVT U218 ( .I(i_data_bus[172]), .ZN(n183) );
  OAI22D1BWP30P140LVT U219 ( .A1(n3), .A2(n184), .B1(n278), .B2(n183), .ZN(
        n185) );
  AOI21D1BWP30P140LVT U220 ( .A1(n281), .A2(i_data_bus[236]), .B(n185), .ZN(
        n187) );
  ND2D1BWP30P140LVT U221 ( .A1(n261), .A2(i_data_bus[12]), .ZN(n186) );
  ND4D1BWP30P140LVT U222 ( .A1(n189), .A2(n188), .A3(n187), .A4(n186), .ZN(
        N381) );
  AOI22D1BWP30P140LVT U223 ( .A1(n275), .A2(i_data_bus[75]), .B1(n257), .B2(
        i_data_bus[43]), .ZN(n196) );
  AOI22D1BWP30P140LVT U224 ( .A1(n2), .A2(i_data_bus[107]), .B1(n258), .B2(
        i_data_bus[139]), .ZN(n195) );
  INVD1BWP30P140LVT U225 ( .I(i_data_bus[203]), .ZN(n191) );
  INVD1BWP30P140LVT U226 ( .I(i_data_bus[171]), .ZN(n190) );
  OAI22D1BWP30P140LVT U227 ( .A1(n3), .A2(n191), .B1(n278), .B2(n190), .ZN(
        n192) );
  AOI21D1BWP30P140LVT U228 ( .A1(n281), .A2(i_data_bus[235]), .B(n192), .ZN(
        n194) );
  ND2D1BWP30P140LVT U229 ( .A1(n261), .A2(i_data_bus[11]), .ZN(n193) );
  ND4D1BWP30P140LVT U230 ( .A1(n196), .A2(n195), .A3(n194), .A4(n193), .ZN(
        N380) );
  AOI22D1BWP30P140LVT U231 ( .A1(n275), .A2(i_data_bus[74]), .B1(n257), .B2(
        i_data_bus[42]), .ZN(n203) );
  AOI22D1BWP30P140LVT U232 ( .A1(n2), .A2(i_data_bus[106]), .B1(n258), .B2(
        i_data_bus[138]), .ZN(n202) );
  INVD1BWP30P140LVT U233 ( .I(i_data_bus[202]), .ZN(n198) );
  INVD1BWP30P140LVT U234 ( .I(i_data_bus[170]), .ZN(n197) );
  OAI22D1BWP30P140LVT U235 ( .A1(n3), .A2(n198), .B1(n278), .B2(n197), .ZN(
        n199) );
  AOI21D1BWP30P140LVT U236 ( .A1(n281), .A2(i_data_bus[234]), .B(n199), .ZN(
        n201) );
  ND2D1BWP30P140LVT U237 ( .A1(n261), .A2(i_data_bus[10]), .ZN(n200) );
  ND4D1BWP30P140LVT U238 ( .A1(n203), .A2(n202), .A3(n201), .A4(n200), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U239 ( .A1(n275), .A2(i_data_bus[73]), .B1(n257), .B2(
        i_data_bus[41]), .ZN(n210) );
  AOI22D1BWP30P140LVT U240 ( .A1(n2), .A2(i_data_bus[105]), .B1(n258), .B2(
        i_data_bus[137]), .ZN(n209) );
  INVD1BWP30P140LVT U241 ( .I(i_data_bus[201]), .ZN(n205) );
  INVD1BWP30P140LVT U242 ( .I(i_data_bus[169]), .ZN(n204) );
  OAI22D1BWP30P140LVT U243 ( .A1(n3), .A2(n205), .B1(n278), .B2(n204), .ZN(
        n206) );
  AOI21D1BWP30P140LVT U244 ( .A1(n281), .A2(i_data_bus[233]), .B(n206), .ZN(
        n208) );
  ND2D1BWP30P140LVT U245 ( .A1(n261), .A2(i_data_bus[9]), .ZN(n207) );
  ND4D1BWP30P140LVT U246 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U247 ( .A1(n275), .A2(i_data_bus[71]), .B1(n257), .B2(
        i_data_bus[39]), .ZN(n217) );
  AOI22D1BWP30P140LVT U248 ( .A1(n2), .A2(i_data_bus[103]), .B1(n258), .B2(
        i_data_bus[135]), .ZN(n216) );
  INVD1BWP30P140LVT U249 ( .I(i_data_bus[199]), .ZN(n212) );
  INVD1BWP30P140LVT U250 ( .I(i_data_bus[167]), .ZN(n211) );
  OAI22D1BWP30P140LVT U251 ( .A1(n3), .A2(n212), .B1(n278), .B2(n211), .ZN(
        n213) );
  AOI21D1BWP30P140LVT U252 ( .A1(n281), .A2(i_data_bus[231]), .B(n213), .ZN(
        n215) );
  ND2D1BWP30P140LVT U253 ( .A1(n261), .A2(i_data_bus[7]), .ZN(n214) );
  ND4D1BWP30P140LVT U254 ( .A1(n217), .A2(n216), .A3(n215), .A4(n214), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U255 ( .A1(n275), .A2(i_data_bus[70]), .B1(n257), .B2(
        i_data_bus[38]), .ZN(n224) );
  AOI22D1BWP30P140LVT U256 ( .A1(n2), .A2(i_data_bus[102]), .B1(n258), .B2(
        i_data_bus[134]), .ZN(n223) );
  INVD1BWP30P140LVT U257 ( .I(i_data_bus[198]), .ZN(n219) );
  INVD1BWP30P140LVT U258 ( .I(i_data_bus[166]), .ZN(n218) );
  OAI22D1BWP30P140LVT U259 ( .A1(n3), .A2(n219), .B1(n278), .B2(n218), .ZN(
        n220) );
  AOI21D1BWP30P140LVT U260 ( .A1(n281), .A2(i_data_bus[230]), .B(n220), .ZN(
        n222) );
  ND2D1BWP30P140LVT U261 ( .A1(n261), .A2(i_data_bus[6]), .ZN(n221) );
  ND4D1BWP30P140LVT U262 ( .A1(n224), .A2(n223), .A3(n222), .A4(n221), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U263 ( .A1(n275), .A2(i_data_bus[69]), .B1(n257), .B2(
        i_data_bus[37]), .ZN(n231) );
  AOI22D1BWP30P140LVT U264 ( .A1(n2), .A2(i_data_bus[101]), .B1(n258), .B2(
        i_data_bus[133]), .ZN(n230) );
  INVD1BWP30P140LVT U265 ( .I(i_data_bus[197]), .ZN(n226) );
  INVD1BWP30P140LVT U266 ( .I(i_data_bus[165]), .ZN(n225) );
  OAI22D1BWP30P140LVT U267 ( .A1(n3), .A2(n226), .B1(n278), .B2(n225), .ZN(
        n227) );
  AOI21D1BWP30P140LVT U268 ( .A1(n281), .A2(i_data_bus[229]), .B(n227), .ZN(
        n229) );
  ND2D1BWP30P140LVT U269 ( .A1(n261), .A2(i_data_bus[5]), .ZN(n228) );
  ND4D1BWP30P140LVT U270 ( .A1(n231), .A2(n230), .A3(n229), .A4(n228), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U271 ( .A1(n275), .A2(i_data_bus[64]), .B1(n257), .B2(
        i_data_bus[32]), .ZN(n237) );
  AOI22D1BWP30P140LVT U272 ( .A1(n2), .A2(i_data_bus[96]), .B1(n258), .B2(
        i_data_bus[128]), .ZN(n236) );
  INR2D1BWP30P140LVT U273 ( .A1(i_data_bus[192]), .B1(n3), .ZN(n233) );
  INR2D1BWP30P140LVT U274 ( .A1(i_data_bus[160]), .B1(n278), .ZN(n232) );
  AOI211D1BWP30P140LVT U275 ( .A1(i_data_bus[224]), .A2(n281), .B(n233), .C(
        n232), .ZN(n235) );
  ND2D1BWP30P140LVT U276 ( .A1(n261), .A2(i_data_bus[0]), .ZN(n234) );
  ND4D1BWP30P140LVT U277 ( .A1(n237), .A2(n236), .A3(n235), .A4(n234), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U278 ( .A1(n275), .A2(i_data_bus[68]), .B1(n257), .B2(
        i_data_bus[36]), .ZN(n244) );
  AOI22D1BWP30P140LVT U279 ( .A1(n2), .A2(i_data_bus[100]), .B1(n258), .B2(
        i_data_bus[132]), .ZN(n243) );
  INVD1BWP30P140LVT U280 ( .I(i_data_bus[196]), .ZN(n239) );
  INVD1BWP30P140LVT U281 ( .I(i_data_bus[164]), .ZN(n238) );
  OAI22D1BWP30P140LVT U282 ( .A1(n3), .A2(n239), .B1(n278), .B2(n238), .ZN(
        n240) );
  AOI21D1BWP30P140LVT U283 ( .A1(n281), .A2(i_data_bus[228]), .B(n240), .ZN(
        n242) );
  ND2D1BWP30P140LVT U284 ( .A1(n261), .A2(i_data_bus[4]), .ZN(n241) );
  ND4D1BWP30P140LVT U285 ( .A1(n244), .A2(n243), .A3(n242), .A4(n241), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U286 ( .A1(n275), .A2(i_data_bus[67]), .B1(n257), .B2(
        i_data_bus[35]), .ZN(n250) );
  AOI22D1BWP30P140LVT U287 ( .A1(n2), .A2(i_data_bus[99]), .B1(n258), .B2(
        i_data_bus[131]), .ZN(n249) );
  INVD1BWP30P140LVT U288 ( .I(i_data_bus[163]), .ZN(n245) );
  MOAI22D1BWP30P140LVT U289 ( .A1(n278), .A2(n245), .B1(n266), .B2(
        i_data_bus[195]), .ZN(n246) );
  AOI21D1BWP30P140LVT U290 ( .A1(n281), .A2(i_data_bus[227]), .B(n246), .ZN(
        n248) );
  ND2D1BWP30P140LVT U291 ( .A1(n261), .A2(i_data_bus[3]), .ZN(n247) );
  ND4D1BWP30P140LVT U292 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U293 ( .A1(n275), .A2(i_data_bus[66]), .B1(n257), .B2(
        i_data_bus[34]), .ZN(n256) );
  AOI22D1BWP30P140LVT U294 ( .A1(n2), .A2(i_data_bus[98]), .B1(n258), .B2(
        i_data_bus[130]), .ZN(n255) );
  INVD1BWP30P140LVT U295 ( .I(i_data_bus[162]), .ZN(n251) );
  MOAI22D1BWP30P140LVT U296 ( .A1(n278), .A2(n251), .B1(n266), .B2(
        i_data_bus[194]), .ZN(n252) );
  AOI21D1BWP30P140LVT U297 ( .A1(n281), .A2(i_data_bus[226]), .B(n252), .ZN(
        n254) );
  ND2D1BWP30P140LVT U298 ( .A1(n261), .A2(i_data_bus[2]), .ZN(n253) );
  ND4D1BWP30P140LVT U299 ( .A1(n256), .A2(n255), .A3(n254), .A4(n253), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U300 ( .A1(n275), .A2(i_data_bus[65]), .B1(n257), .B2(
        i_data_bus[33]), .ZN(n265) );
  AOI22D1BWP30P140LVT U301 ( .A1(n2), .A2(i_data_bus[97]), .B1(n258), .B2(
        i_data_bus[129]), .ZN(n264) );
  INVD1BWP30P140LVT U302 ( .I(i_data_bus[161]), .ZN(n259) );
  MOAI22D1BWP30P140LVT U303 ( .A1(n278), .A2(n259), .B1(n266), .B2(
        i_data_bus[193]), .ZN(n260) );
  AOI21D1BWP30P140LVT U304 ( .A1(n281), .A2(i_data_bus[225]), .B(n260), .ZN(
        n263) );
  ND2D1BWP30P140LVT U305 ( .A1(n261), .A2(i_data_bus[1]), .ZN(n262) );
  ND4D1BWP30P140LVT U306 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U307 ( .A1(n275), .A2(i_data_bus[78]), .B1(n274), .B2(
        i_data_bus[46]), .ZN(n273) );
  AOI22D1BWP30P140LVT U308 ( .A1(n2), .A2(i_data_bus[110]), .B1(n276), .B2(
        i_data_bus[142]), .ZN(n272) );
  INVD1BWP30P140LVT U309 ( .I(i_data_bus[174]), .ZN(n267) );
  MOAI22D1BWP30P140LVT U310 ( .A1(n278), .A2(n267), .B1(n266), .B2(
        i_data_bus[206]), .ZN(n268) );
  AOI21D1BWP30P140LVT U311 ( .A1(n269), .A2(i_data_bus[238]), .B(n268), .ZN(
        n271) );
  ND2D1BWP30P140LVT U312 ( .A1(n282), .A2(i_data_bus[14]), .ZN(n270) );
  ND4D1BWP30P140LVT U313 ( .A1(n273), .A2(n272), .A3(n271), .A4(n270), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U314 ( .A1(n275), .A2(i_data_bus[77]), .B1(n274), .B2(
        i_data_bus[45]), .ZN(n286) );
  AOI22D1BWP30P140LVT U315 ( .A1(n2), .A2(i_data_bus[109]), .B1(n276), .B2(
        i_data_bus[141]), .ZN(n285) );
  INVD1BWP30P140LVT U316 ( .I(i_data_bus[205]), .ZN(n279) );
  INVD1BWP30P140LVT U317 ( .I(i_data_bus[173]), .ZN(n277) );
  OAI22D1BWP30P140LVT U318 ( .A1(n3), .A2(n279), .B1(n278), .B2(n277), .ZN(
        n280) );
  AOI21D1BWP30P140LVT U319 ( .A1(n281), .A2(i_data_bus[237]), .B(n280), .ZN(
        n284) );
  ND2D1BWP30P140LVT U320 ( .A1(n282), .A2(i_data_bus[13]), .ZN(n283) );
  ND4D1BWP30P140LVT U321 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_15 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  BUFFD4BWP30P140LVT U3 ( .I(n51), .Z(n259) );
  OR2D1BWP30P140LVT U4 ( .A1(n44), .A2(n35), .Z(n126) );
  INR2D1BWP30P140LVT U5 ( .A1(n25), .B1(n24), .ZN(n26) );
  INVD1BWP30P140LVT U6 ( .I(n153), .ZN(n95) );
  INVD3BWP30P140LVT U7 ( .I(n126), .ZN(n1) );
  INVD2BWP30P140LVT U8 ( .I(i_cmd[7]), .ZN(n23) );
  NR2D1BWP30P140LVT U9 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n16) );
  INVD3BWP30P140LVT U10 ( .I(n50), .ZN(n285) );
  ND2OPTIBD2BWP30P140LVT U11 ( .A1(n32), .A2(n31), .ZN(n44) );
  NR2D1BWP30P140LVT U12 ( .A1(n29), .A2(i_cmd[4]), .ZN(n32) );
  NR2D1BWP30P140LVT U13 ( .A1(i_cmd[5]), .A2(n30), .ZN(n31) );
  ND2D1BWP30P140LVT U14 ( .A1(n13), .A2(n12), .ZN(n20) );
  ND2OPTIBD1BWP30P140LVT U15 ( .A1(n4), .A2(n23), .ZN(n30) );
  ND2OPTIBD6BWP30P140LVT U16 ( .A1(n14), .A2(n17), .ZN(n153) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n16), .A2(n15), .Z(n17) );
  INVD1BWP30P140LVT U18 ( .I(n39), .ZN(n50) );
  INVD1BWP30P140LVT U19 ( .I(n10), .ZN(n130) );
  INVD1BWP30P140LVT U20 ( .I(n130), .ZN(n270) );
  INVD1BWP30P140LVT U21 ( .I(n130), .ZN(n292) );
  INR4D0BWP30P140LVT U22 ( .A1(i_valid[2]), .B1(i_cmd[1]), .B2(i_cmd[3]), .B3(
        n40), .ZN(n41) );
  INR2D4BWP30P140LVT U23 ( .A1(n45), .B1(n44), .ZN(n283) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n47), .A2(n46), .Z(n2) );
  INVD1BWP30P140LVT U25 ( .I(i_cmd[0]), .ZN(n3) );
  INR3D0BWP30P140LVT U26 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n3), .ZN(n9) );
  OR2D1BWP30P140LVT U27 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n43) );
  INVD1BWP30P140LVT U28 ( .I(n43), .ZN(n8) );
  INVD1BWP30P140LVT U29 ( .I(i_cmd[6]), .ZN(n4) );
  INVD1BWP30P140LVT U30 ( .I(rst), .ZN(n5) );
  ND2D1BWP30P140LVT U31 ( .A1(n5), .A2(i_en), .ZN(n28) );
  OR2D1BWP30P140LVT U32 ( .A1(i_cmd[1]), .A2(n28), .Z(n6) );
  NR3D0P7BWP30P140LVT U33 ( .A1(n30), .A2(i_cmd[5]), .A3(n6), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U34 ( .A1(n8), .A2(n7), .ZN(n37) );
  INR2D1BWP30P140LVT U35 ( .A1(n9), .B1(n37), .ZN(n10) );
  INVD1BWP30P140LVT U36 ( .I(n130), .ZN(n146) );
  INVD2BWP30P140LVT U37 ( .I(i_cmd[1]), .ZN(n11) );
  INVD2BWP30P140LVT U38 ( .I(i_cmd[2]), .ZN(n40) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(n11), .A2(n40), .ZN(n34) );
  OR2D1BWP30P140LVT U40 ( .A1(n34), .A2(i_cmd[4]), .Z(n18) );
  NR2D1BWP30P140LVT U41 ( .A1(i_cmd[0]), .A2(n28), .ZN(n13) );
  INVD1BWP30P140LVT U42 ( .I(i_cmd[3]), .ZN(n12) );
  NR2OPTPAD1BWP30P140LVT U43 ( .A1(n18), .A2(n20), .ZN(n14) );
  CKAN2D1BWP30P140LVT U44 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n15) );
  NR2D1BWP30P140LVT U45 ( .A1(n30), .A2(n18), .ZN(n22) );
  ND2D1BWP30P140LVT U46 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n19) );
  NR2D1BWP30P140LVT U47 ( .A1(n20), .A2(n19), .ZN(n21) );
  CKND2D2BWP30P140LVT U48 ( .A1(n22), .A2(n21), .ZN(n51) );
  INVD1BWP30P140LVT U49 ( .I(n259), .ZN(n27) );
  INR4D0BWP30P140LVT U50 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n23), .ZN(n25) );
  INVD1BWP30P140LVT U51 ( .I(n14), .ZN(n24) );
  INVD2BWP30P140LVT U52 ( .I(n26), .ZN(n118) );
  INVD2BWP30P140LVT U53 ( .I(n118), .ZN(n291) );
  NR4D0BWP30P140LVT U54 ( .A1(n146), .A2(n95), .A3(n27), .A4(n291), .ZN(n49)
         );
  OR2D1BWP30P140LVT U55 ( .A1(i_cmd[0]), .A2(n28), .Z(n29) );
  ND2OPTIBD1BWP30P140LVT U56 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n33) );
  OR2D1BWP30P140LVT U57 ( .A1(n34), .A2(n33), .Z(n35) );
  ND2OPTIBD1BWP30P140LVT U58 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n36) );
  NR2D1BWP30P140LVT U59 ( .A1(n36), .A2(i_cmd[0]), .ZN(n38) );
  INR2D1BWP30P140LVT U60 ( .A1(n38), .B1(n37), .ZN(n39) );
  NR2D1BWP30P140LVT U61 ( .A1(n1), .A2(n285), .ZN(n48) );
  INR2D2BWP30P140LVT U62 ( .A1(n41), .B1(n44), .ZN(n151) );
  INVD1BWP30P140LVT U63 ( .I(n151), .ZN(n47) );
  ND2D1BWP30P140LVT U64 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n42) );
  NR2D1BWP30P140LVT U65 ( .A1(n43), .A2(n42), .ZN(n45) );
  INVD1BWP30P140LVT U66 ( .I(n283), .ZN(n46) );
  ND3D1BWP30P140LVT U67 ( .A1(n49), .A2(n48), .A3(n2), .ZN(N402) );
  BUFFD4BWP30P140LVT U68 ( .I(n151), .Z(n284) );
  AOI22D1BWP30P140LVT U69 ( .A1(n284), .A2(i_data_bus[68]), .B1(n283), .B2(
        i_data_bus[36]), .ZN(n59) );
  INVD2BWP30P140LVT U70 ( .I(n50), .ZN(n266) );
  AOI22D1BWP30P140LVT U71 ( .A1(n1), .A2(i_data_bus[100]), .B1(n266), .B2(
        i_data_bus[132]), .ZN(n58) );
  INVD1BWP30P140LVT U72 ( .I(i_data_bus[196]), .ZN(n54) );
  INVD2BWP30P140LVT U73 ( .I(n51), .ZN(n52) );
  INVD2BWP30P140LVT U74 ( .I(n52), .ZN(n287) );
  INVD1BWP30P140LVT U75 ( .I(i_data_bus[164]), .ZN(n53) );
  OAI22D1BWP30P140LVT U76 ( .A1(n153), .A2(n54), .B1(n287), .B2(n53), .ZN(n55)
         );
  AOI21D1BWP30P140LVT U77 ( .A1(n291), .A2(i_data_bus[228]), .B(n55), .ZN(n57)
         );
  ND2D1BWP30P140LVT U78 ( .A1(n270), .A2(i_data_bus[4]), .ZN(n56) );
  ND4D1BWP30P140LVT U79 ( .A1(n59), .A2(n58), .A3(n57), .A4(n56), .ZN(N373) );
  AOI22D1BWP30P140LVT U80 ( .A1(n284), .A2(i_data_bus[67]), .B1(n283), .B2(
        i_data_bus[35]), .ZN(n66) );
  AOI22D1BWP30P140LVT U81 ( .A1(n1), .A2(i_data_bus[99]), .B1(n266), .B2(
        i_data_bus[131]), .ZN(n65) );
  INVD1BWP30P140LVT U82 ( .I(i_data_bus[195]), .ZN(n61) );
  INVD1BWP30P140LVT U83 ( .I(i_data_bus[163]), .ZN(n60) );
  OAI22D1BWP30P140LVT U84 ( .A1(n153), .A2(n61), .B1(n287), .B2(n60), .ZN(n62)
         );
  AOI21D1BWP30P140LVT U85 ( .A1(n291), .A2(i_data_bus[227]), .B(n62), .ZN(n64)
         );
  ND2D1BWP30P140LVT U86 ( .A1(n270), .A2(i_data_bus[3]), .ZN(n63) );
  ND4D1BWP30P140LVT U87 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(N372) );
  AOI22D1BWP30P140LVT U88 ( .A1(n284), .A2(i_data_bus[75]), .B1(n283), .B2(
        i_data_bus[43]), .ZN(n73) );
  AOI22D1BWP30P140LVT U89 ( .A1(n1), .A2(i_data_bus[107]), .B1(n266), .B2(
        i_data_bus[139]), .ZN(n72) );
  INVD1BWP30P140LVT U90 ( .I(i_data_bus[203]), .ZN(n68) );
  INVD1BWP30P140LVT U91 ( .I(i_data_bus[171]), .ZN(n67) );
  OAI22D1BWP30P140LVT U92 ( .A1(n153), .A2(n68), .B1(n287), .B2(n67), .ZN(n69)
         );
  AOI21D1BWP30P140LVT U93 ( .A1(n291), .A2(i_data_bus[235]), .B(n69), .ZN(n71)
         );
  ND2D1BWP30P140LVT U94 ( .A1(n270), .A2(i_data_bus[11]), .ZN(n70) );
  ND4D1BWP30P140LVT U95 ( .A1(n73), .A2(n72), .A3(n71), .A4(n70), .ZN(N380) );
  AOI22D1BWP30P140LVT U96 ( .A1(n284), .A2(i_data_bus[69]), .B1(n283), .B2(
        i_data_bus[37]), .ZN(n80) );
  AOI22D1BWP30P140LVT U97 ( .A1(n1), .A2(i_data_bus[101]), .B1(n266), .B2(
        i_data_bus[133]), .ZN(n79) );
  INVD1BWP30P140LVT U98 ( .I(i_data_bus[197]), .ZN(n75) );
  INVD1BWP30P140LVT U99 ( .I(i_data_bus[165]), .ZN(n74) );
  OAI22D1BWP30P140LVT U100 ( .A1(n153), .A2(n75), .B1(n287), .B2(n74), .ZN(n76) );
  AOI21D1BWP30P140LVT U101 ( .A1(n291), .A2(i_data_bus[229]), .B(n76), .ZN(n78) );
  ND2D1BWP30P140LVT U102 ( .A1(n270), .A2(i_data_bus[5]), .ZN(n77) );
  ND4D1BWP30P140LVT U103 ( .A1(n80), .A2(n79), .A3(n78), .A4(n77), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U104 ( .A1(n284), .A2(i_data_bus[66]), .B1(n283), .B2(
        i_data_bus[34]), .ZN(n87) );
  AOI22D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[98]), .B1(n266), .B2(
        i_data_bus[130]), .ZN(n86) );
  INVD1BWP30P140LVT U106 ( .I(i_data_bus[194]), .ZN(n82) );
  INVD1BWP30P140LVT U107 ( .I(i_data_bus[162]), .ZN(n81) );
  OAI22D1BWP30P140LVT U108 ( .A1(n153), .A2(n82), .B1(n287), .B2(n81), .ZN(n83) );
  AOI21D1BWP30P140LVT U109 ( .A1(n291), .A2(i_data_bus[226]), .B(n83), .ZN(n85) );
  ND2D1BWP30P140LVT U110 ( .A1(n270), .A2(i_data_bus[2]), .ZN(n84) );
  ND4D1BWP30P140LVT U111 ( .A1(n87), .A2(n86), .A3(n85), .A4(n84), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U112 ( .A1(n284), .A2(i_data_bus[76]), .B1(n283), .B2(
        i_data_bus[44]), .ZN(n94) );
  AOI22D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[108]), .B1(n266), .B2(
        i_data_bus[140]), .ZN(n93) );
  INVD1BWP30P140LVT U114 ( .I(i_data_bus[172]), .ZN(n89) );
  ND2D1BWP30P140LVT U115 ( .A1(n95), .A2(i_data_bus[204]), .ZN(n88) );
  OAI21D1BWP30P140LVT U116 ( .A1(n287), .A2(n89), .B(n88), .ZN(n90) );
  AOI21D1BWP30P140LVT U117 ( .A1(n291), .A2(i_data_bus[236]), .B(n90), .ZN(n92) );
  ND2D1BWP30P140LVT U118 ( .A1(n270), .A2(i_data_bus[12]), .ZN(n91) );
  ND4D1BWP30P140LVT U119 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .ZN(N381)
         );
  AOI22D1BWP30P140LVT U120 ( .A1(n151), .A2(i_data_bus[93]), .B1(n283), .B2(
        i_data_bus[61]), .ZN(n102) );
  AOI22D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[125]), .B1(n285), .B2(
        i_data_bus[157]), .ZN(n101) );
  INVD1BWP30P140LVT U122 ( .I(n118), .ZN(n113) );
  INVD2BWP30P140LVT U123 ( .I(n95), .ZN(n144) );
  INVD1BWP30P140LVT U124 ( .I(i_data_bus[221]), .ZN(n97) );
  INVD1BWP30P140LVT U125 ( .I(i_data_bus[189]), .ZN(n96) );
  OAI22D1BWP30P140LVT U126 ( .A1(n144), .A2(n97), .B1(n259), .B2(n96), .ZN(n98) );
  AOI21D1BWP30P140LVT U127 ( .A1(n113), .A2(i_data_bus[253]), .B(n98), .ZN(
        n100) );
  ND2D1BWP30P140LVT U128 ( .A1(n146), .A2(i_data_bus[29]), .ZN(n99) );
  ND4D1BWP30P140LVT U129 ( .A1(n102), .A2(n101), .A3(n100), .A4(n99), .ZN(N398) );
  AOI22D1BWP30P140LVT U130 ( .A1(n151), .A2(i_data_bus[94]), .B1(n283), .B2(
        i_data_bus[62]), .ZN(n109) );
  AOI22D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[126]), .B1(n285), .B2(
        i_data_bus[158]), .ZN(n108) );
  INVD1BWP30P140LVT U132 ( .I(i_data_bus[222]), .ZN(n104) );
  INVD1BWP30P140LVT U133 ( .I(i_data_bus[190]), .ZN(n103) );
  OAI22D1BWP30P140LVT U134 ( .A1(n144), .A2(n104), .B1(n259), .B2(n103), .ZN(
        n105) );
  AOI21D1BWP30P140LVT U135 ( .A1(n113), .A2(i_data_bus[254]), .B(n105), .ZN(
        n107) );
  ND2D1BWP30P140LVT U136 ( .A1(n146), .A2(i_data_bus[30]), .ZN(n106) );
  ND4D1BWP30P140LVT U137 ( .A1(n109), .A2(n108), .A3(n107), .A4(n106), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U138 ( .A1(n151), .A2(i_data_bus[92]), .B1(n283), .B2(
        i_data_bus[60]), .ZN(n117) );
  AOI22D1BWP30P140LVT U139 ( .A1(n1), .A2(i_data_bus[124]), .B1(n285), .B2(
        i_data_bus[156]), .ZN(n116) );
  INVD1BWP30P140LVT U140 ( .I(i_data_bus[220]), .ZN(n111) );
  INVD1BWP30P140LVT U141 ( .I(i_data_bus[188]), .ZN(n110) );
  OAI22D1BWP30P140LVT U142 ( .A1(n144), .A2(n111), .B1(n259), .B2(n110), .ZN(
        n112) );
  AOI21D1BWP30P140LVT U143 ( .A1(n113), .A2(i_data_bus[252]), .B(n112), .ZN(
        n115) );
  ND2D1BWP30P140LVT U144 ( .A1(n146), .A2(i_data_bus[28]), .ZN(n114) );
  ND4D1BWP30P140LVT U145 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U146 ( .A1(n151), .A2(i_data_bus[91]), .B1(n283), .B2(
        i_data_bus[59]), .ZN(n125) );
  AOI22D1BWP30P140LVT U147 ( .A1(n1), .A2(i_data_bus[123]), .B1(n285), .B2(
        i_data_bus[155]), .ZN(n124) );
  INVD2BWP30P140LVT U148 ( .I(n118), .ZN(n278) );
  INVD1BWP30P140LVT U149 ( .I(i_data_bus[219]), .ZN(n120) );
  INVD1BWP30P140LVT U150 ( .I(i_data_bus[187]), .ZN(n119) );
  OAI22D1BWP30P140LVT U151 ( .A1(n144), .A2(n120), .B1(n259), .B2(n119), .ZN(
        n121) );
  AOI21D1BWP30P140LVT U152 ( .A1(n278), .A2(i_data_bus[251]), .B(n121), .ZN(
        n123) );
  ND2D1BWP30P140LVT U153 ( .A1(n146), .A2(i_data_bus[27]), .ZN(n122) );
  ND4D1BWP30P140LVT U154 ( .A1(n125), .A2(n124), .A3(n123), .A4(n122), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U155 ( .A1(n284), .A2(i_data_bus[89]), .B1(n283), .B2(
        i_data_bus[57]), .ZN(n134) );
  AOI22D1BWP30P140LVT U156 ( .A1(n1), .A2(i_data_bus[121]), .B1(n285), .B2(
        i_data_bus[153]), .ZN(n133) );
  INVD1BWP30P140LVT U157 ( .I(i_data_bus[217]), .ZN(n128) );
  INVD1BWP30P140LVT U158 ( .I(i_data_bus[185]), .ZN(n127) );
  OAI22D1BWP30P140LVT U159 ( .A1(n144), .A2(n128), .B1(n259), .B2(n127), .ZN(
        n129) );
  AOI21D1BWP30P140LVT U160 ( .A1(n278), .A2(i_data_bus[249]), .B(n129), .ZN(
        n132) );
  ND2D1BWP30P140LVT U161 ( .A1(n292), .A2(i_data_bus[25]), .ZN(n131) );
  ND4D1BWP30P140LVT U162 ( .A1(n134), .A2(n133), .A3(n132), .A4(n131), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U163 ( .A1(n151), .A2(i_data_bus[90]), .B1(n283), .B2(
        i_data_bus[58]), .ZN(n141) );
  AOI22D1BWP30P140LVT U164 ( .A1(n1), .A2(i_data_bus[122]), .B1(n285), .B2(
        i_data_bus[154]), .ZN(n140) );
  INVD1BWP30P140LVT U165 ( .I(i_data_bus[218]), .ZN(n136) );
  INVD1BWP30P140LVT U166 ( .I(i_data_bus[186]), .ZN(n135) );
  OAI22D1BWP30P140LVT U167 ( .A1(n144), .A2(n136), .B1(n259), .B2(n135), .ZN(
        n137) );
  AOI21D1BWP30P140LVT U168 ( .A1(n278), .A2(i_data_bus[250]), .B(n137), .ZN(
        n139) );
  ND2D1BWP30P140LVT U169 ( .A1(n146), .A2(i_data_bus[26]), .ZN(n138) );
  ND4D1BWP30P140LVT U170 ( .A1(n141), .A2(n140), .A3(n139), .A4(n138), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U171 ( .A1(n151), .A2(i_data_bus[95]), .B1(n283), .B2(
        i_data_bus[63]), .ZN(n150) );
  AOI22D1BWP30P140LVT U172 ( .A1(n1), .A2(i_data_bus[127]), .B1(n285), .B2(
        i_data_bus[159]), .ZN(n149) );
  INVD1BWP30P140LVT U173 ( .I(i_data_bus[223]), .ZN(n143) );
  INVD1BWP30P140LVT U174 ( .I(i_data_bus[191]), .ZN(n142) );
  OAI22D1BWP30P140LVT U175 ( .A1(n144), .A2(n143), .B1(n259), .B2(n142), .ZN(
        n145) );
  AOI21D1BWP30P140LVT U176 ( .A1(n291), .A2(i_data_bus[255]), .B(n145), .ZN(
        n148) );
  ND2D1BWP30P140LVT U177 ( .A1(n146), .A2(i_data_bus[31]), .ZN(n147) );
  ND4D1BWP30P140LVT U178 ( .A1(n150), .A2(n149), .A3(n148), .A4(n147), .ZN(
        N400) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n151), .A2(i_data_bus[64]), .Z(n152) );
  AOI21D1BWP30P140LVT U180 ( .A1(n283), .A2(i_data_bus[32]), .B(n152), .ZN(
        n159) );
  AOI22D1BWP30P140LVT U181 ( .A1(n1), .A2(i_data_bus[96]), .B1(n266), .B2(
        i_data_bus[128]), .ZN(n158) );
  BUFFD4BWP30P140LVT U182 ( .I(n153), .Z(n289) );
  INR2D1BWP30P140LVT U183 ( .A1(i_data_bus[192]), .B1(n289), .ZN(n155) );
  INR2D1BWP30P140LVT U184 ( .A1(i_data_bus[160]), .B1(n287), .ZN(n154) );
  AOI211D1BWP30P140LVT U185 ( .A1(i_data_bus[224]), .A2(n291), .B(n155), .C(
        n154), .ZN(n157) );
  ND2D1BWP30P140LVT U186 ( .A1(n270), .A2(i_data_bus[0]), .ZN(n156) );
  ND4D1BWP30P140LVT U187 ( .A1(n159), .A2(n158), .A3(n157), .A4(n156), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U188 ( .A1(n284), .A2(i_data_bus[72]), .B1(n283), .B2(
        i_data_bus[40]), .ZN(n166) );
  AOI22D1BWP30P140LVT U189 ( .A1(n1), .A2(i_data_bus[104]), .B1(n266), .B2(
        i_data_bus[136]), .ZN(n165) );
  INVD1BWP30P140LVT U190 ( .I(i_data_bus[200]), .ZN(n161) );
  INVD1BWP30P140LVT U191 ( .I(i_data_bus[168]), .ZN(n160) );
  OAI22D1BWP30P140LVT U192 ( .A1(n289), .A2(n161), .B1(n287), .B2(n160), .ZN(
        n162) );
  AOI21D1BWP30P140LVT U193 ( .A1(n278), .A2(i_data_bus[232]), .B(n162), .ZN(
        n164) );
  ND2D1BWP30P140LVT U194 ( .A1(n270), .A2(i_data_bus[8]), .ZN(n163) );
  ND4D1BWP30P140LVT U195 ( .A1(n166), .A2(n165), .A3(n164), .A4(n163), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U196 ( .A1(n284), .A2(i_data_bus[70]), .B1(n283), .B2(
        i_data_bus[38]), .ZN(n173) );
  AOI22D1BWP30P140LVT U197 ( .A1(n1), .A2(i_data_bus[102]), .B1(n266), .B2(
        i_data_bus[134]), .ZN(n172) );
  INVD1BWP30P140LVT U198 ( .I(i_data_bus[198]), .ZN(n168) );
  INVD1BWP30P140LVT U199 ( .I(i_data_bus[166]), .ZN(n167) );
  OAI22D1BWP30P140LVT U200 ( .A1(n289), .A2(n168), .B1(n287), .B2(n167), .ZN(
        n169) );
  AOI21D1BWP30P140LVT U201 ( .A1(n291), .A2(i_data_bus[230]), .B(n169), .ZN(
        n171) );
  ND2D1BWP30P140LVT U202 ( .A1(n270), .A2(i_data_bus[6]), .ZN(n170) );
  ND4D1BWP30P140LVT U203 ( .A1(n173), .A2(n172), .A3(n171), .A4(n170), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U204 ( .A1(n284), .A2(i_data_bus[71]), .B1(n283), .B2(
        i_data_bus[39]), .ZN(n180) );
  AOI22D1BWP30P140LVT U205 ( .A1(n1), .A2(i_data_bus[103]), .B1(n266), .B2(
        i_data_bus[135]), .ZN(n179) );
  INVD1BWP30P140LVT U206 ( .I(i_data_bus[199]), .ZN(n175) );
  INVD1BWP30P140LVT U207 ( .I(i_data_bus[167]), .ZN(n174) );
  OAI22D1BWP30P140LVT U208 ( .A1(n289), .A2(n175), .B1(n287), .B2(n174), .ZN(
        n176) );
  AOI21D1BWP30P140LVT U209 ( .A1(n291), .A2(i_data_bus[231]), .B(n176), .ZN(
        n178) );
  ND2D1BWP30P140LVT U210 ( .A1(n270), .A2(i_data_bus[7]), .ZN(n177) );
  ND4D1BWP30P140LVT U211 ( .A1(n180), .A2(n179), .A3(n178), .A4(n177), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U212 ( .A1(n284), .A2(i_data_bus[74]), .B1(n283), .B2(
        i_data_bus[42]), .ZN(n187) );
  AOI22D1BWP30P140LVT U213 ( .A1(n1), .A2(i_data_bus[106]), .B1(n266), .B2(
        i_data_bus[138]), .ZN(n186) );
  INVD1BWP30P140LVT U214 ( .I(i_data_bus[202]), .ZN(n182) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[170]), .ZN(n181) );
  OAI22D1BWP30P140LVT U216 ( .A1(n289), .A2(n182), .B1(n287), .B2(n181), .ZN(
        n183) );
  AOI21D1BWP30P140LVT U217 ( .A1(n291), .A2(i_data_bus[234]), .B(n183), .ZN(
        n185) );
  ND2D1BWP30P140LVT U218 ( .A1(n270), .A2(i_data_bus[10]), .ZN(n184) );
  ND4D1BWP30P140LVT U219 ( .A1(n187), .A2(n186), .A3(n185), .A4(n184), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U220 ( .A1(n284), .A2(i_data_bus[73]), .B1(n283), .B2(
        i_data_bus[41]), .ZN(n194) );
  AOI22D1BWP30P140LVT U221 ( .A1(n1), .A2(i_data_bus[105]), .B1(n266), .B2(
        i_data_bus[137]), .ZN(n193) );
  INVD1BWP30P140LVT U222 ( .I(i_data_bus[201]), .ZN(n189) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[169]), .ZN(n188) );
  OAI22D1BWP30P140LVT U224 ( .A1(n289), .A2(n189), .B1(n287), .B2(n188), .ZN(
        n190) );
  AOI21D1BWP30P140LVT U225 ( .A1(n291), .A2(i_data_bus[233]), .B(n190), .ZN(
        n192) );
  ND2D1BWP30P140LVT U226 ( .A1(n270), .A2(i_data_bus[9]), .ZN(n191) );
  ND4D1BWP30P140LVT U227 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U228 ( .A1(n284), .A2(i_data_bus[84]), .B1(n283), .B2(
        i_data_bus[52]), .ZN(n201) );
  AOI22D1BWP30P140LVT U229 ( .A1(n1), .A2(i_data_bus[116]), .B1(n285), .B2(
        i_data_bus[148]), .ZN(n200) );
  INVD1BWP30P140LVT U230 ( .I(i_data_bus[212]), .ZN(n196) );
  INVD1BWP30P140LVT U231 ( .I(i_data_bus[180]), .ZN(n195) );
  OAI22D1BWP30P140LVT U232 ( .A1(n289), .A2(n196), .B1(n259), .B2(n195), .ZN(
        n197) );
  AOI21D1BWP30P140LVT U233 ( .A1(n278), .A2(i_data_bus[244]), .B(n197), .ZN(
        n199) );
  ND2D1BWP30P140LVT U234 ( .A1(n292), .A2(i_data_bus[20]), .ZN(n198) );
  ND4D1BWP30P140LVT U235 ( .A1(n201), .A2(n200), .A3(n199), .A4(n198), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U236 ( .A1(n284), .A2(i_data_bus[82]), .B1(n283), .B2(
        i_data_bus[50]), .ZN(n208) );
  AOI22D1BWP30P140LVT U237 ( .A1(n1), .A2(i_data_bus[114]), .B1(n285), .B2(
        i_data_bus[146]), .ZN(n207) );
  INVD1BWP30P140LVT U238 ( .I(i_data_bus[210]), .ZN(n203) );
  INVD1BWP30P140LVT U239 ( .I(i_data_bus[178]), .ZN(n202) );
  OAI22D1BWP30P140LVT U240 ( .A1(n289), .A2(n203), .B1(n259), .B2(n202), .ZN(
        n204) );
  AOI21D1BWP30P140LVT U241 ( .A1(n278), .A2(i_data_bus[242]), .B(n204), .ZN(
        n206) );
  ND2D1BWP30P140LVT U242 ( .A1(n292), .A2(i_data_bus[18]), .ZN(n205) );
  ND4D1BWP30P140LVT U243 ( .A1(n208), .A2(n207), .A3(n206), .A4(n205), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U244 ( .A1(n284), .A2(i_data_bus[83]), .B1(n283), .B2(
        i_data_bus[51]), .ZN(n215) );
  AOI22D1BWP30P140LVT U245 ( .A1(n1), .A2(i_data_bus[115]), .B1(n285), .B2(
        i_data_bus[147]), .ZN(n214) );
  INVD1BWP30P140LVT U246 ( .I(i_data_bus[211]), .ZN(n210) );
  INVD1BWP30P140LVT U247 ( .I(i_data_bus[179]), .ZN(n209) );
  OAI22D1BWP30P140LVT U248 ( .A1(n289), .A2(n210), .B1(n259), .B2(n209), .ZN(
        n211) );
  AOI21D1BWP30P140LVT U249 ( .A1(n278), .A2(i_data_bus[243]), .B(n211), .ZN(
        n213) );
  ND2D1BWP30P140LVT U250 ( .A1(n292), .A2(i_data_bus[19]), .ZN(n212) );
  ND4D1BWP30P140LVT U251 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U252 ( .A1(n284), .A2(i_data_bus[87]), .B1(n283), .B2(
        i_data_bus[55]), .ZN(n222) );
  AOI22D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[119]), .B1(n285), .B2(
        i_data_bus[151]), .ZN(n221) );
  INVD1BWP30P140LVT U254 ( .I(i_data_bus[215]), .ZN(n217) );
  INVD1BWP30P140LVT U255 ( .I(i_data_bus[183]), .ZN(n216) );
  OAI22D1BWP30P140LVT U256 ( .A1(n289), .A2(n217), .B1(n259), .B2(n216), .ZN(
        n218) );
  AOI21D1BWP30P140LVT U257 ( .A1(n278), .A2(i_data_bus[247]), .B(n218), .ZN(
        n220) );
  ND2D1BWP30P140LVT U258 ( .A1(n292), .A2(i_data_bus[23]), .ZN(n219) );
  ND4D1BWP30P140LVT U259 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U260 ( .A1(n284), .A2(i_data_bus[85]), .B1(n283), .B2(
        i_data_bus[53]), .ZN(n229) );
  AOI22D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[117]), .B1(n285), .B2(
        i_data_bus[149]), .ZN(n228) );
  INVD1BWP30P140LVT U262 ( .I(i_data_bus[213]), .ZN(n224) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[181]), .ZN(n223) );
  OAI22D1BWP30P140LVT U264 ( .A1(n289), .A2(n224), .B1(n259), .B2(n223), .ZN(
        n225) );
  AOI21D1BWP30P140LVT U265 ( .A1(n278), .A2(i_data_bus[245]), .B(n225), .ZN(
        n227) );
  ND2D1BWP30P140LVT U266 ( .A1(n292), .A2(i_data_bus[21]), .ZN(n226) );
  ND4D1BWP30P140LVT U267 ( .A1(n229), .A2(n228), .A3(n227), .A4(n226), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U268 ( .A1(n284), .A2(i_data_bus[86]), .B1(n283), .B2(
        i_data_bus[54]), .ZN(n236) );
  AOI22D1BWP30P140LVT U269 ( .A1(n1), .A2(i_data_bus[118]), .B1(n285), .B2(
        i_data_bus[150]), .ZN(n235) );
  INVD1BWP30P140LVT U270 ( .I(i_data_bus[214]), .ZN(n231) );
  INVD1BWP30P140LVT U271 ( .I(i_data_bus[182]), .ZN(n230) );
  OAI22D1BWP30P140LVT U272 ( .A1(n289), .A2(n231), .B1(n259), .B2(n230), .ZN(
        n232) );
  AOI21D1BWP30P140LVT U273 ( .A1(n278), .A2(i_data_bus[246]), .B(n232), .ZN(
        n234) );
  ND2D1BWP30P140LVT U274 ( .A1(n292), .A2(i_data_bus[22]), .ZN(n233) );
  ND4D1BWP30P140LVT U275 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U276 ( .A1(n284), .A2(i_data_bus[80]), .B1(n283), .B2(
        i_data_bus[48]), .ZN(n243) );
  AOI22D1BWP30P140LVT U277 ( .A1(n1), .A2(i_data_bus[112]), .B1(n285), .B2(
        i_data_bus[144]), .ZN(n242) );
  INVD1BWP30P140LVT U278 ( .I(i_data_bus[208]), .ZN(n238) );
  INVD1BWP30P140LVT U279 ( .I(i_data_bus[176]), .ZN(n237) );
  OAI22D1BWP30P140LVT U280 ( .A1(n289), .A2(n238), .B1(n259), .B2(n237), .ZN(
        n239) );
  AOI21D1BWP30P140LVT U281 ( .A1(n278), .A2(i_data_bus[240]), .B(n239), .ZN(
        n241) );
  ND2D1BWP30P140LVT U282 ( .A1(n292), .A2(i_data_bus[16]), .ZN(n240) );
  ND4D1BWP30P140LVT U283 ( .A1(n243), .A2(n242), .A3(n241), .A4(n240), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U284 ( .A1(n284), .A2(i_data_bus[81]), .B1(n283), .B2(
        i_data_bus[49]), .ZN(n250) );
  AOI22D1BWP30P140LVT U285 ( .A1(n1), .A2(i_data_bus[113]), .B1(n285), .B2(
        i_data_bus[145]), .ZN(n249) );
  INVD1BWP30P140LVT U286 ( .I(i_data_bus[209]), .ZN(n245) );
  INVD1BWP30P140LVT U287 ( .I(i_data_bus[177]), .ZN(n244) );
  OAI22D1BWP30P140LVT U288 ( .A1(n289), .A2(n245), .B1(n259), .B2(n244), .ZN(
        n246) );
  AOI21D1BWP30P140LVT U289 ( .A1(n278), .A2(i_data_bus[241]), .B(n246), .ZN(
        n248) );
  ND2D1BWP30P140LVT U290 ( .A1(n292), .A2(i_data_bus[17]), .ZN(n247) );
  ND4D1BWP30P140LVT U291 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U292 ( .A1(n284), .A2(i_data_bus[88]), .B1(n283), .B2(
        i_data_bus[56]), .ZN(n257) );
  AOI22D1BWP30P140LVT U293 ( .A1(n1), .A2(i_data_bus[120]), .B1(n285), .B2(
        i_data_bus[152]), .ZN(n256) );
  INVD1BWP30P140LVT U294 ( .I(i_data_bus[216]), .ZN(n252) );
  INVD1BWP30P140LVT U295 ( .I(i_data_bus[184]), .ZN(n251) );
  OAI22D1BWP30P140LVT U296 ( .A1(n289), .A2(n252), .B1(n259), .B2(n251), .ZN(
        n253) );
  AOI21D1BWP30P140LVT U297 ( .A1(n278), .A2(i_data_bus[248]), .B(n253), .ZN(
        n255) );
  ND2D1BWP30P140LVT U298 ( .A1(n292), .A2(i_data_bus[24]), .ZN(n254) );
  ND4D1BWP30P140LVT U299 ( .A1(n257), .A2(n256), .A3(n255), .A4(n254), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U300 ( .A1(n284), .A2(i_data_bus[79]), .B1(n283), .B2(
        i_data_bus[47]), .ZN(n265) );
  AOI22D1BWP30P140LVT U301 ( .A1(n1), .A2(i_data_bus[111]), .B1(n285), .B2(
        i_data_bus[143]), .ZN(n264) );
  INVD1BWP30P140LVT U302 ( .I(i_data_bus[207]), .ZN(n260) );
  INVD1BWP30P140LVT U303 ( .I(i_data_bus[175]), .ZN(n258) );
  OAI22D1BWP30P140LVT U304 ( .A1(n289), .A2(n260), .B1(n259), .B2(n258), .ZN(
        n261) );
  AOI21D1BWP30P140LVT U305 ( .A1(n278), .A2(i_data_bus[239]), .B(n261), .ZN(
        n263) );
  ND2D1BWP30P140LVT U306 ( .A1(n292), .A2(i_data_bus[15]), .ZN(n262) );
  ND4D1BWP30P140LVT U307 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U308 ( .A1(n284), .A2(i_data_bus[65]), .B1(n283), .B2(
        i_data_bus[33]), .ZN(n274) );
  AOI22D1BWP30P140LVT U309 ( .A1(n1), .A2(i_data_bus[97]), .B1(n266), .B2(
        i_data_bus[129]), .ZN(n273) );
  INVD1BWP30P140LVT U310 ( .I(i_data_bus[193]), .ZN(n268) );
  INVD1BWP30P140LVT U311 ( .I(i_data_bus[161]), .ZN(n267) );
  OAI22D1BWP30P140LVT U312 ( .A1(n289), .A2(n268), .B1(n287), .B2(n267), .ZN(
        n269) );
  AOI21D1BWP30P140LVT U313 ( .A1(n291), .A2(i_data_bus[225]), .B(n269), .ZN(
        n272) );
  ND2D1BWP30P140LVT U314 ( .A1(n270), .A2(i_data_bus[1]), .ZN(n271) );
  ND4D1BWP30P140LVT U315 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U316 ( .A1(n284), .A2(i_data_bus[78]), .B1(n283), .B2(
        i_data_bus[46]), .ZN(n282) );
  AOI22D1BWP30P140LVT U317 ( .A1(n1), .A2(i_data_bus[110]), .B1(n285), .B2(
        i_data_bus[142]), .ZN(n281) );
  INVD1BWP30P140LVT U318 ( .I(i_data_bus[206]), .ZN(n276) );
  INVD1BWP30P140LVT U319 ( .I(i_data_bus[174]), .ZN(n275) );
  OAI22D1BWP30P140LVT U320 ( .A1(n289), .A2(n276), .B1(n287), .B2(n275), .ZN(
        n277) );
  AOI21D1BWP30P140LVT U321 ( .A1(n278), .A2(i_data_bus[238]), .B(n277), .ZN(
        n280) );
  ND2D1BWP30P140LVT U322 ( .A1(n292), .A2(i_data_bus[14]), .ZN(n279) );
  ND4D1BWP30P140LVT U323 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U324 ( .A1(n284), .A2(i_data_bus[77]), .B1(n283), .B2(
        i_data_bus[45]), .ZN(n296) );
  AOI22D1BWP30P140LVT U325 ( .A1(n1), .A2(i_data_bus[109]), .B1(n285), .B2(
        i_data_bus[141]), .ZN(n295) );
  INVD1BWP30P140LVT U326 ( .I(i_data_bus[205]), .ZN(n288) );
  INVD1BWP30P140LVT U327 ( .I(i_data_bus[173]), .ZN(n286) );
  OAI22D1BWP30P140LVT U328 ( .A1(n289), .A2(n288), .B1(n287), .B2(n286), .ZN(
        n290) );
  AOI21D1BWP30P140LVT U329 ( .A1(n291), .A2(i_data_bus[237]), .B(n290), .ZN(
        n294) );
  ND2D1BWP30P140LVT U330 ( .A1(n292), .A2(i_data_bus[13]), .ZN(n293) );
  ND4D1BWP30P140LVT U331 ( .A1(n296), .A2(n295), .A3(n294), .A4(n293), .ZN(
        N382) );
endmodule


module crossbar_8_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA8_0 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [63:0] i_cmd;
  input clk, rst, i_en;

  wire   [63:0] o_inner_cmd_wire;
  wire   [255:0] bottom_half_0__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_0__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_1__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_1__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_2__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_2__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_3__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_3__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_4__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_4__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_5__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_5__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_6__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_6__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_7__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_7__inner_valid_i_mux_tree_wire;

  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 top_half_0__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[0]), .i_data_bus(
        i_data_bus[31:0]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[0], 
        bottom_half_6__inner_valid_i_mux_tree_wire[0], 
        bottom_half_5__inner_valid_i_mux_tree_wire[0], 
        bottom_half_4__inner_valid_i_mux_tree_wire[0], 
        bottom_half_3__inner_valid_i_mux_tree_wire[0], 
        bottom_half_2__inner_valid_i_mux_tree_wire[0], 
        bottom_half_1__inner_valid_i_mux_tree_wire[0], 
        bottom_half_0__inner_valid_i_mux_tree_wire[0]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_6__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_5__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_4__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_3__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_2__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_1__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_0__inner_data_i_mux_tree_wire[31:0]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_15 top_half_1__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[1]), .i_data_bus(
        i_data_bus[63:32]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[1], 
        bottom_half_6__inner_valid_i_mux_tree_wire[1], 
        bottom_half_5__inner_valid_i_mux_tree_wire[1], 
        bottom_half_4__inner_valid_i_mux_tree_wire[1], 
        bottom_half_3__inner_valid_i_mux_tree_wire[1], 
        bottom_half_2__inner_valid_i_mux_tree_wire[1], 
        bottom_half_1__inner_valid_i_mux_tree_wire[1], 
        bottom_half_0__inner_valid_i_mux_tree_wire[1]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_6__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_5__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_4__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_3__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_2__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_1__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_0__inner_data_i_mux_tree_wire[63:32]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_14 top_half_2__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[2]), .i_data_bus(
        i_data_bus[95:64]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[2], 
        bottom_half_6__inner_valid_i_mux_tree_wire[2], 
        bottom_half_5__inner_valid_i_mux_tree_wire[2], 
        bottom_half_4__inner_valid_i_mux_tree_wire[2], 
        bottom_half_3__inner_valid_i_mux_tree_wire[2], 
        bottom_half_2__inner_valid_i_mux_tree_wire[2], 
        bottom_half_1__inner_valid_i_mux_tree_wire[2], 
        bottom_half_0__inner_valid_i_mux_tree_wire[2]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_6__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_5__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_4__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_3__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_2__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_1__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_0__inner_data_i_mux_tree_wire[95:64]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_13 top_half_3__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[3]), .i_data_bus(
        i_data_bus[127:96]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[3], 
        bottom_half_6__inner_valid_i_mux_tree_wire[3], 
        bottom_half_5__inner_valid_i_mux_tree_wire[3], 
        bottom_half_4__inner_valid_i_mux_tree_wire[3], 
        bottom_half_3__inner_valid_i_mux_tree_wire[3], 
        bottom_half_2__inner_valid_i_mux_tree_wire[3], 
        bottom_half_1__inner_valid_i_mux_tree_wire[3], 
        bottom_half_0__inner_valid_i_mux_tree_wire[3]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_6__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_5__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_4__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_3__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_2__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_1__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_0__inner_data_i_mux_tree_wire[127:96]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_12 top_half_4__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[4]), .i_data_bus(
        i_data_bus[159:128]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[4], 
        bottom_half_6__inner_valid_i_mux_tree_wire[4], 
        bottom_half_5__inner_valid_i_mux_tree_wire[4], 
        bottom_half_4__inner_valid_i_mux_tree_wire[4], 
        bottom_half_3__inner_valid_i_mux_tree_wire[4], 
        bottom_half_2__inner_valid_i_mux_tree_wire[4], 
        bottom_half_1__inner_valid_i_mux_tree_wire[4], 
        bottom_half_0__inner_valid_i_mux_tree_wire[4]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_6__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_5__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_4__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_3__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_2__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_1__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_0__inner_data_i_mux_tree_wire[159:128]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_11 top_half_5__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[5]), .i_data_bus(
        i_data_bus[191:160]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[5], 
        bottom_half_6__inner_valid_i_mux_tree_wire[5], 
        bottom_half_5__inner_valid_i_mux_tree_wire[5], 
        bottom_half_4__inner_valid_i_mux_tree_wire[5], 
        bottom_half_3__inner_valid_i_mux_tree_wire[5], 
        bottom_half_2__inner_valid_i_mux_tree_wire[5], 
        bottom_half_1__inner_valid_i_mux_tree_wire[5], 
        bottom_half_0__inner_valid_i_mux_tree_wire[5]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_6__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_5__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_4__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_3__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_2__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_1__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_0__inner_data_i_mux_tree_wire[191:160]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_10 top_half_6__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[6]), .i_data_bus(
        i_data_bus[223:192]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[6], 
        bottom_half_6__inner_valid_i_mux_tree_wire[6], 
        bottom_half_5__inner_valid_i_mux_tree_wire[6], 
        bottom_half_4__inner_valid_i_mux_tree_wire[6], 
        bottom_half_3__inner_valid_i_mux_tree_wire[6], 
        bottom_half_2__inner_valid_i_mux_tree_wire[6], 
        bottom_half_1__inner_valid_i_mux_tree_wire[6], 
        bottom_half_0__inner_valid_i_mux_tree_wire[6]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_6__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_5__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_4__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_3__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_2__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_1__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_0__inner_data_i_mux_tree_wire[223:192]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_9 top_half_7__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[7]), .i_data_bus(
        i_data_bus[255:224]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[7], 
        bottom_half_6__inner_valid_i_mux_tree_wire[7], 
        bottom_half_5__inner_valid_i_mux_tree_wire[7], 
        bottom_half_4__inner_valid_i_mux_tree_wire[7], 
        bottom_half_3__inner_valid_i_mux_tree_wire[7], 
        bottom_half_2__inner_valid_i_mux_tree_wire[7], 
        bottom_half_1__inner_valid_i_mux_tree_wire[7], 
        bottom_half_0__inner_valid_i_mux_tree_wire[7]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_6__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_5__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_4__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_3__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_2__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_1__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_0__inner_data_i_mux_tree_wire[255:224]}), .i_en(i_en) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 i_cmd_id_0__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[0]), .o_cmd_1(
        o_inner_cmd_wire[8]), .o_cmd_2(o_inner_cmd_wire[16]), .o_cmd_3(
        o_inner_cmd_wire[24]), .o_cmd_4(o_inner_cmd_wire[32]), .o_cmd_5(
        o_inner_cmd_wire[40]), .o_cmd_6(o_inner_cmd_wire[48]), .o_cmd_7(
        o_inner_cmd_wire[56]), .i_en(i_en), .i_cmd(i_cmd[7:0]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_15 i_cmd_id_1__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[1]), .o_cmd_1(
        o_inner_cmd_wire[9]), .o_cmd_2(o_inner_cmd_wire[17]), .o_cmd_3(
        o_inner_cmd_wire[25]), .o_cmd_4(o_inner_cmd_wire[33]), .o_cmd_5(
        o_inner_cmd_wire[41]), .o_cmd_6(o_inner_cmd_wire[49]), .o_cmd_7(
        o_inner_cmd_wire[57]), .i_en(i_en), .i_cmd(i_cmd[15:8]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_14 i_cmd_id_2__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[2]), .o_cmd_1(
        o_inner_cmd_wire[10]), .o_cmd_2(o_inner_cmd_wire[18]), .o_cmd_3(
        o_inner_cmd_wire[26]), .o_cmd_4(o_inner_cmd_wire[34]), .o_cmd_5(
        o_inner_cmd_wire[42]), .o_cmd_6(o_inner_cmd_wire[50]), .o_cmd_7(
        o_inner_cmd_wire[58]), .i_en(i_en), .i_cmd(i_cmd[23:16]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_13 i_cmd_id_3__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[3]), .o_cmd_1(
        o_inner_cmd_wire[11]), .o_cmd_2(o_inner_cmd_wire[19]), .o_cmd_3(
        o_inner_cmd_wire[27]), .o_cmd_4(o_inner_cmd_wire[35]), .o_cmd_5(
        o_inner_cmd_wire[43]), .o_cmd_6(o_inner_cmd_wire[51]), .o_cmd_7(
        o_inner_cmd_wire[59]), .i_en(i_en), .i_cmd(i_cmd[31:24]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_12 i_cmd_id_4__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[4]), .o_cmd_1(
        o_inner_cmd_wire[12]), .o_cmd_2(o_inner_cmd_wire[20]), .o_cmd_3(
        o_inner_cmd_wire[28]), .o_cmd_4(o_inner_cmd_wire[36]), .o_cmd_5(
        o_inner_cmd_wire[44]), .o_cmd_6(o_inner_cmd_wire[52]), .o_cmd_7(
        o_inner_cmd_wire[60]), .i_en(i_en), .i_cmd(i_cmd[39:32]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_11 i_cmd_id_5__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[5]), .o_cmd_1(
        o_inner_cmd_wire[13]), .o_cmd_2(o_inner_cmd_wire[21]), .o_cmd_3(
        o_inner_cmd_wire[29]), .o_cmd_4(o_inner_cmd_wire[37]), .o_cmd_5(
        o_inner_cmd_wire[45]), .o_cmd_6(o_inner_cmd_wire[53]), .o_cmd_7(
        o_inner_cmd_wire[61]), .i_en(i_en), .i_cmd(i_cmd[47:40]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_10 i_cmd_id_6__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[6]), .o_cmd_1(
        o_inner_cmd_wire[14]), .o_cmd_2(o_inner_cmd_wire[22]), .o_cmd_3(
        o_inner_cmd_wire[30]), .o_cmd_4(o_inner_cmd_wire[38]), .o_cmd_5(
        o_inner_cmd_wire[46]), .o_cmd_6(o_inner_cmd_wire[54]), .o_cmd_7(
        o_inner_cmd_wire[62]), .i_en(i_en), .i_cmd(i_cmd[55:48]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_9 i_cmd_id_7__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[7]), .o_cmd_1(
        o_inner_cmd_wire[15]), .o_cmd_2(o_inner_cmd_wire[23]), .o_cmd_3(
        o_inner_cmd_wire[31]), .o_cmd_4(o_inner_cmd_wire[39]), .o_cmd_5(
        o_inner_cmd_wire[47]), .o_cmd_6(o_inner_cmd_wire[55]), .o_cmd_7(
        o_inner_cmd_wire[63]), .i_en(i_en), .i_cmd(i_cmd[63:56]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_0 bottom_half_0__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_0__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_0__inner_data_i_mux_tree_wire), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[7:0]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_15 bottom_half_1__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_1__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_1__inner_data_i_mux_tree_wire), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[15:8]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_14 bottom_half_2__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_2__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_2__inner_data_i_mux_tree_wire), .o_valid(o_valid[2]), 
        .o_data_bus(o_data_bus[95:64]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[23:16]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_13 bottom_half_3__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_3__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_3__inner_data_i_mux_tree_wire), .o_valid(o_valid[3]), 
        .o_data_bus(o_data_bus[127:96]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[31:24]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_12 bottom_half_4__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_4__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_4__inner_data_i_mux_tree_wire), .o_valid(o_valid[4]), 
        .o_data_bus(o_data_bus[159:128]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[39:32]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_11 bottom_half_5__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_5__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_5__inner_data_i_mux_tree_wire), .o_valid(o_valid[5]), 
        .o_data_bus(o_data_bus[191:160]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[47:40]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_10 bottom_half_6__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_6__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_6__inner_data_i_mux_tree_wire), .o_valid(o_valid[6]), 
        .o_data_bus(o_data_bus[223:192]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[55:48]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_9 bottom_half_7__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_7__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_7__inner_data_i_mux_tree_wire), .o_valid(o_valid[7]), 
        .o_data_bus(o_data_bus[255:224]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[63:56]) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_8 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), 
        .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), 
        .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), 
        .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), 
        .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), 
        .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), 
        .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), 
        .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), 
        .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), 
        .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), 
        .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_8 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_1 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INR2D6BWP30P140LVT U3 ( .A1(n43), .B1(n42), .ZN(n280) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n36), .A2(n35), .Z(n1) );
  ND2D2BWP30P140LVT U5 ( .A1(n3), .A2(n1), .ZN(n72) );
  NR2OPTPAD1BWP30P140LVT U6 ( .A1(n19), .A2(n34), .ZN(n23) );
  INVD3BWP30P140LVT U7 ( .I(n271), .ZN(n177) );
  INVD2BWP30P140LVT U8 ( .I(n71), .ZN(n279) );
  ND2OPTIBD2BWP30P140LVT U9 ( .A1(n48), .A2(n1), .ZN(n71) );
  NR2D2BWP30P140LVT U10 ( .A1(n19), .A2(n21), .ZN(n25) );
  OR2D1BWP30P140LVT U11 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n50) );
  ND2D1BWP30P140LVT U12 ( .A1(n23), .A2(n22), .ZN(n74) );
  ND2D1BWP30P140LVT U13 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n20) );
  INVD1BWP30P140LVT U14 ( .I(n50), .ZN(n43) );
  ND2D1BWP30P140LVT U15 ( .A1(n8), .A2(n7), .ZN(n38) );
  AN2D2BWP30P140LVT U16 ( .A1(n37), .A2(n1), .Z(n2) );
  INVD1BWP30P140LVT U17 ( .I(n72), .ZN(n174) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n52), .A2(n51), .Z(n3) );
  INVD1BWP30P140LVT U19 ( .I(n28), .ZN(n73) );
  INVD1BWP30P140LVT U20 ( .I(i_cmd[0]), .ZN(n4) );
  INR3D0BWP30P140LVT U21 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n4), .ZN(n10)
         );
  OR2D2BWP30P140LVT U22 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n34) );
  NR2OPTPAD1BWP30P140LVT U23 ( .A1(n34), .A2(i_cmd[5]), .ZN(n8) );
  INVD1BWP30P140LVT U24 ( .I(rst), .ZN(n5) );
  ND2D1BWP30P140LVT U25 ( .A1(n5), .A2(i_en), .ZN(n33) );
  INVD1BWP30P140LVT U26 ( .I(n33), .ZN(n6) );
  INR2D1BWP30P140LVT U27 ( .A1(n6), .B1(i_cmd[1]), .ZN(n7) );
  IND2D1BWP30P140LVT U28 ( .A1(n38), .B1(n43), .ZN(n9) );
  INR2D1BWP30P140LVT U29 ( .A1(n10), .B1(n9), .ZN(n11) );
  INVD2BWP30P140LVT U30 ( .I(n11), .ZN(n179) );
  INVD1BWP30P140LVT U31 ( .I(n179), .ZN(n169) );
  ND2D1BWP30P140LVT U32 ( .A1(i_cmd[6]), .A2(i_valid[6]), .ZN(n17) );
  NR2D1BWP30P140LVT U33 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n16) );
  OR2D4BWP30P140LVT U34 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .Z(n31) );
  INVD1BWP30P140LVT U35 ( .I(n31), .ZN(n13) );
  NR2OPTPAD1BWP30P140LVT U36 ( .A1(i_cmd[0]), .A2(n33), .ZN(n12) );
  ND2OPTIBD2BWP30P140LVT U37 ( .A1(n13), .A2(n12), .ZN(n19) );
  INVD1BWP30P140LVT U38 ( .I(i_cmd[3]), .ZN(n15) );
  INVD1BWP30P140LVT U39 ( .I(i_cmd[4]), .ZN(n14) );
  ND2OPTIBD1BWP30P140LVT U40 ( .A1(n15), .A2(n14), .ZN(n21) );
  IND3D4BWP30P140LVT U41 ( .A1(n17), .B1(n16), .B2(n25), .ZN(n18) );
  INVD4BWP30P140LVT U42 ( .I(n18), .ZN(n271) );
  NR2D1BWP30P140LVT U43 ( .A1(n21), .A2(n20), .ZN(n22) );
  BUFFD4BWP30P140LVT U44 ( .I(n74), .Z(n244) );
  INVD1BWP30P140LVT U45 ( .I(n244), .ZN(n29) );
  INVD1BWP30P140LVT U46 ( .I(i_cmd[7]), .ZN(n24) );
  INR4D0BWP30P140LVT U47 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n24), .ZN(n27) );
  INVD1BWP30P140LVT U48 ( .I(n25), .ZN(n26) );
  INR2D1BWP30P140LVT U49 ( .A1(n27), .B1(n26), .ZN(n28) );
  INVD2BWP30P140LVT U50 ( .I(n73), .ZN(n286) );
  NR4D0BWP30P140LVT U51 ( .A1(n169), .A2(n271), .A3(n29), .A4(n286), .ZN(n54)
         );
  NR2D1BWP30P140LVT U52 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n51) );
  ND2D1BWP30P140LVT U53 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n30) );
  OR2D1BWP30P140LVT U54 ( .A1(n31), .A2(n30), .Z(n32) );
  INR2D1BWP30P140LVT U55 ( .A1(n51), .B1(n32), .ZN(n37) );
  NR2D1BWP30P140LVT U56 ( .A1(i_cmd[5]), .A2(n33), .ZN(n36) );
  INVD1BWP30P140LVT U57 ( .I(n34), .ZN(n35) );
  INVD1BWP30P140LVT U58 ( .I(n38), .ZN(n41) );
  ND2D1BWP30P140LVT U59 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n39) );
  NR2D1BWP30P140LVT U60 ( .A1(n39), .A2(i_cmd[0]), .ZN(n40) );
  ND2D2BWP30P140LVT U61 ( .A1(n41), .A2(n40), .ZN(n42) );
  NR2D1BWP30P140LVT U62 ( .A1(n2), .A2(n280), .ZN(n53) );
  NR2D1BWP30P140LVT U63 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .ZN(n44) );
  ND2D1BWP30P140LVT U64 ( .A1(n51), .A2(n44), .ZN(n47) );
  INVD1BWP30P140LVT U65 ( .I(i_cmd[2]), .ZN(n46) );
  INVD1BWP30P140LVT U66 ( .I(i_valid[2]), .ZN(n45) );
  NR3D0P7BWP30P140LVT U67 ( .A1(n47), .A2(n46), .A3(n45), .ZN(n48) );
  ND2D1BWP30P140LVT U68 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n49) );
  NR2D1BWP30P140LVT U69 ( .A1(n50), .A2(n49), .ZN(n52) );
  ND4D1BWP30P140LVT U70 ( .A1(n54), .A2(n53), .A3(n71), .A4(n72), .ZN(N402) );
  INR2D1BWP30P140LVT U71 ( .A1(i_data_bus[63]), .B1(n72), .ZN(n56) );
  INR2D1BWP30P140LVT U72 ( .A1(i_data_bus[95]), .B1(n71), .ZN(n55) );
  NR2D1BWP30P140LVT U73 ( .A1(n56), .A2(n55), .ZN(n63) );
  AOI22D1BWP30P140LVT U74 ( .A1(n2), .A2(i_data_bus[127]), .B1(n280), .B2(
        i_data_bus[159]), .ZN(n62) );
  INVD1BWP30P140LVT U75 ( .I(i_data_bus[223]), .ZN(n58) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[191]), .ZN(n57) );
  OAI22D1BWP30P140LVT U77 ( .A1(n177), .A2(n58), .B1(n244), .B2(n57), .ZN(n59)
         );
  AOI21D1BWP30P140LVT U78 ( .A1(n286), .A2(i_data_bus[255]), .B(n59), .ZN(n61)
         );
  ND2D1BWP30P140LVT U79 ( .A1(n169), .A2(i_data_bus[31]), .ZN(n60) );
  ND4D1BWP30P140LVT U80 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(N400) );
  AOI22D1BWP30P140LVT U81 ( .A1(n279), .A2(i_data_bus[94]), .B1(n174), .B2(
        i_data_bus[62]), .ZN(n70) );
  AOI22D1BWP30P140LVT U82 ( .A1(n2), .A2(i_data_bus[126]), .B1(n280), .B2(
        i_data_bus[158]), .ZN(n69) );
  INVD1BWP30P140LVT U83 ( .I(i_data_bus[222]), .ZN(n65) );
  INVD1BWP30P140LVT U84 ( .I(i_data_bus[190]), .ZN(n64) );
  OAI22D1BWP30P140LVT U85 ( .A1(n177), .A2(n65), .B1(n244), .B2(n64), .ZN(n66)
         );
  AOI21D1BWP30P140LVT U86 ( .A1(n274), .A2(i_data_bus[254]), .B(n66), .ZN(n68)
         );
  ND2D1BWP30P140LVT U87 ( .A1(n169), .A2(i_data_bus[30]), .ZN(n67) );
  ND4D1BWP30P140LVT U88 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(N399) );
  INVD2BWP30P140LVT U89 ( .I(n71), .ZN(n263) );
  INVD2BWP30P140LVT U90 ( .I(n72), .ZN(n262) );
  AOI22D1BWP30P140LVT U91 ( .A1(n263), .A2(i_data_bus[72]), .B1(n262), .B2(
        i_data_bus[40]), .ZN(n82) );
  AOI22D1BWP30P140LVT U92 ( .A1(n2), .A2(i_data_bus[104]), .B1(n280), .B2(
        i_data_bus[136]), .ZN(n81) );
  INVD2BWP30P140LVT U93 ( .I(n73), .ZN(n274) );
  INVD2BWP30P140LVT U94 ( .I(n74), .ZN(n75) );
  INVD3BWP30P140LVT U95 ( .I(n75), .ZN(n282) );
  INVD1BWP30P140LVT U96 ( .I(i_data_bus[168]), .ZN(n77) );
  INVD1BWP30P140LVT U97 ( .I(i_data_bus[200]), .ZN(n76) );
  OAI22D1BWP30P140LVT U98 ( .A1(n282), .A2(n77), .B1(n177), .B2(n76), .ZN(n78)
         );
  AOI21OPTREPBD1BWP30P140LVT U99 ( .A1(n274), .A2(i_data_bus[232]), .B(n78), 
        .ZN(n80) );
  INVD2BWP30P140LVT U100 ( .I(n179), .ZN(n266) );
  ND2D1BWP30P140LVT U101 ( .A1(n266), .A2(i_data_bus[8]), .ZN(n79) );
  ND4D1BWP30P140LVT U102 ( .A1(n82), .A2(n81), .A3(n80), .A4(n79), .ZN(N377)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n263), .A2(i_data_bus[76]), .B1(n262), .B2(
        i_data_bus[44]), .ZN(n89) );
  AOI22D1BWP30P140LVT U104 ( .A1(n2), .A2(i_data_bus[108]), .B1(n280), .B2(
        i_data_bus[140]), .ZN(n88) );
  INVD6BWP30P140LVT U105 ( .I(n271), .ZN(n284) );
  INVD1BWP30P140LVT U106 ( .I(i_data_bus[204]), .ZN(n84) );
  INVD1BWP30P140LVT U107 ( .I(i_data_bus[172]), .ZN(n83) );
  OAI22D1BWP30P140LVT U108 ( .A1(n284), .A2(n84), .B1(n282), .B2(n83), .ZN(n85) );
  AOI21D1BWP30P140LVT U109 ( .A1(n286), .A2(i_data_bus[236]), .B(n85), .ZN(n87) );
  ND2D1BWP30P140LVT U110 ( .A1(n266), .A2(i_data_bus[12]), .ZN(n86) );
  ND4D1BWP30P140LVT U111 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(N381)
         );
  AOI22D1BWP30P140LVT U112 ( .A1(n263), .A2(i_data_bus[75]), .B1(n262), .B2(
        i_data_bus[43]), .ZN(n96) );
  AOI22D1BWP30P140LVT U113 ( .A1(n2), .A2(i_data_bus[107]), .B1(n280), .B2(
        i_data_bus[139]), .ZN(n95) );
  INVD1BWP30P140LVT U114 ( .I(i_data_bus[203]), .ZN(n91) );
  INVD1BWP30P140LVT U115 ( .I(i_data_bus[171]), .ZN(n90) );
  OAI22D1BWP30P140LVT U116 ( .A1(n284), .A2(n91), .B1(n282), .B2(n90), .ZN(n92) );
  AOI21D1BWP30P140LVT U117 ( .A1(n286), .A2(i_data_bus[235]), .B(n92), .ZN(n94) );
  ND2D1BWP30P140LVT U118 ( .A1(n266), .A2(i_data_bus[11]), .ZN(n93) );
  ND4D1BWP30P140LVT U119 ( .A1(n96), .A2(n95), .A3(n94), .A4(n93), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U120 ( .A1(n263), .A2(i_data_bus[74]), .B1(n262), .B2(
        i_data_bus[42]), .ZN(n103) );
  AOI22D1BWP30P140LVT U121 ( .A1(n2), .A2(i_data_bus[106]), .B1(n280), .B2(
        i_data_bus[138]), .ZN(n102) );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[202]), .ZN(n98) );
  INVD1BWP30P140LVT U123 ( .I(i_data_bus[170]), .ZN(n97) );
  OAI22D1BWP30P140LVT U124 ( .A1(n284), .A2(n98), .B1(n282), .B2(n97), .ZN(n99) );
  AOI21D1BWP30P140LVT U125 ( .A1(n286), .A2(i_data_bus[234]), .B(n99), .ZN(
        n101) );
  ND2D1BWP30P140LVT U126 ( .A1(n266), .A2(i_data_bus[10]), .ZN(n100) );
  ND4D1BWP30P140LVT U127 ( .A1(n103), .A2(n102), .A3(n101), .A4(n100), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U128 ( .A1(n263), .A2(i_data_bus[73]), .B1(n262), .B2(
        i_data_bus[41]), .ZN(n110) );
  AOI22D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[105]), .B1(n280), .B2(
        i_data_bus[137]), .ZN(n109) );
  INVD1BWP30P140LVT U130 ( .I(i_data_bus[201]), .ZN(n105) );
  INVD1BWP30P140LVT U131 ( .I(i_data_bus[169]), .ZN(n104) );
  OAI22D1BWP30P140LVT U132 ( .A1(n284), .A2(n105), .B1(n282), .B2(n104), .ZN(
        n106) );
  AOI21D1BWP30P140LVT U133 ( .A1(n286), .A2(i_data_bus[233]), .B(n106), .ZN(
        n108) );
  ND2D1BWP30P140LVT U134 ( .A1(n266), .A2(i_data_bus[9]), .ZN(n107) );
  ND4D1BWP30P140LVT U135 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U136 ( .A1(n263), .A2(i_data_bus[71]), .B1(n262), .B2(
        i_data_bus[39]), .ZN(n117) );
  AOI22D1BWP30P140LVT U137 ( .A1(n2), .A2(i_data_bus[103]), .B1(n280), .B2(
        i_data_bus[135]), .ZN(n116) );
  INVD1BWP30P140LVT U138 ( .I(i_data_bus[199]), .ZN(n112) );
  INVD1BWP30P140LVT U139 ( .I(i_data_bus[167]), .ZN(n111) );
  OAI22D1BWP30P140LVT U140 ( .A1(n284), .A2(n112), .B1(n282), .B2(n111), .ZN(
        n113) );
  AOI21D1BWP30P140LVT U141 ( .A1(n286), .A2(i_data_bus[231]), .B(n113), .ZN(
        n115) );
  ND2D1BWP30P140LVT U142 ( .A1(n266), .A2(i_data_bus[7]), .ZN(n114) );
  ND4D1BWP30P140LVT U143 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U144 ( .A1(n263), .A2(i_data_bus[70]), .B1(n262), .B2(
        i_data_bus[38]), .ZN(n124) );
  AOI22D1BWP30P140LVT U145 ( .A1(n2), .A2(i_data_bus[102]), .B1(n280), .B2(
        i_data_bus[134]), .ZN(n123) );
  INVD1BWP30P140LVT U146 ( .I(i_data_bus[198]), .ZN(n119) );
  INVD1BWP30P140LVT U147 ( .I(i_data_bus[166]), .ZN(n118) );
  OAI22D1BWP30P140LVT U148 ( .A1(n284), .A2(n119), .B1(n282), .B2(n118), .ZN(
        n120) );
  AOI21D1BWP30P140LVT U149 ( .A1(n286), .A2(i_data_bus[230]), .B(n120), .ZN(
        n122) );
  ND2D1BWP30P140LVT U150 ( .A1(n266), .A2(i_data_bus[6]), .ZN(n121) );
  ND4D1BWP30P140LVT U151 ( .A1(n124), .A2(n123), .A3(n122), .A4(n121), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U152 ( .A1(n263), .A2(i_data_bus[69]), .B1(n262), .B2(
        i_data_bus[37]), .ZN(n131) );
  AOI22D1BWP30P140LVT U153 ( .A1(n2), .A2(i_data_bus[101]), .B1(n280), .B2(
        i_data_bus[133]), .ZN(n130) );
  INVD1BWP30P140LVT U154 ( .I(i_data_bus[197]), .ZN(n126) );
  INVD1BWP30P140LVT U155 ( .I(i_data_bus[165]), .ZN(n125) );
  OAI22D1BWP30P140LVT U156 ( .A1(n284), .A2(n126), .B1(n282), .B2(n125), .ZN(
        n127) );
  AOI21D1BWP30P140LVT U157 ( .A1(n286), .A2(i_data_bus[229]), .B(n127), .ZN(
        n129) );
  ND2D1BWP30P140LVT U158 ( .A1(n266), .A2(i_data_bus[5]), .ZN(n128) );
  ND4D1BWP30P140LVT U159 ( .A1(n131), .A2(n130), .A3(n129), .A4(n128), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U160 ( .A1(n263), .A2(i_data_bus[68]), .B1(n262), .B2(
        i_data_bus[36]), .ZN(n138) );
  AOI22D1BWP30P140LVT U161 ( .A1(n2), .A2(i_data_bus[100]), .B1(n280), .B2(
        i_data_bus[132]), .ZN(n137) );
  INVD1BWP30P140LVT U162 ( .I(i_data_bus[196]), .ZN(n133) );
  INVD1BWP30P140LVT U163 ( .I(i_data_bus[164]), .ZN(n132) );
  OAI22D1BWP30P140LVT U164 ( .A1(n284), .A2(n133), .B1(n282), .B2(n132), .ZN(
        n134) );
  AOI21D1BWP30P140LVT U165 ( .A1(n286), .A2(i_data_bus[228]), .B(n134), .ZN(
        n136) );
  ND2D1BWP30P140LVT U166 ( .A1(n266), .A2(i_data_bus[4]), .ZN(n135) );
  ND4D1BWP30P140LVT U167 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U168 ( .A1(n263), .A2(i_data_bus[67]), .B1(n262), .B2(
        i_data_bus[35]), .ZN(n144) );
  AOI22D1BWP30P140LVT U169 ( .A1(n2), .A2(i_data_bus[99]), .B1(n280), .B2(
        i_data_bus[131]), .ZN(n143) );
  INVD1BWP30P140LVT U170 ( .I(i_data_bus[163]), .ZN(n139) );
  MOAI22D1BWP30P140LVT U171 ( .A1(n282), .A2(n139), .B1(n271), .B2(
        i_data_bus[195]), .ZN(n140) );
  AOI21D1BWP30P140LVT U172 ( .A1(n286), .A2(i_data_bus[227]), .B(n140), .ZN(
        n142) );
  ND2D1BWP30P140LVT U173 ( .A1(n266), .A2(i_data_bus[3]), .ZN(n141) );
  ND4D1BWP30P140LVT U174 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U175 ( .A1(n279), .A2(i_data_bus[93]), .B1(n174), .B2(
        i_data_bus[61]), .ZN(n151) );
  AOI22D1BWP30P140LVT U176 ( .A1(n2), .A2(i_data_bus[125]), .B1(n280), .B2(
        i_data_bus[157]), .ZN(n150) );
  INVD1BWP30P140LVT U177 ( .I(i_data_bus[221]), .ZN(n146) );
  INVD1BWP30P140LVT U178 ( .I(i_data_bus[189]), .ZN(n145) );
  OAI22D1BWP30P140LVT U179 ( .A1(n177), .A2(n146), .B1(n244), .B2(n145), .ZN(
        n147) );
  AOI21D1BWP30P140LVT U180 ( .A1(n274), .A2(i_data_bus[253]), .B(n147), .ZN(
        n149) );
  ND2D1BWP30P140LVT U181 ( .A1(n169), .A2(i_data_bus[29]), .ZN(n148) );
  ND4D1BWP30P140LVT U182 ( .A1(n151), .A2(n150), .A3(n149), .A4(n148), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U183 ( .A1(n279), .A2(i_data_bus[92]), .B1(n174), .B2(
        i_data_bus[60]), .ZN(n158) );
  AOI22D1BWP30P140LVT U184 ( .A1(n2), .A2(i_data_bus[124]), .B1(n280), .B2(
        i_data_bus[156]), .ZN(n157) );
  INVD1BWP30P140LVT U185 ( .I(i_data_bus[220]), .ZN(n153) );
  INVD1BWP30P140LVT U186 ( .I(i_data_bus[188]), .ZN(n152) );
  OAI22D1BWP30P140LVT U187 ( .A1(n177), .A2(n153), .B1(n244), .B2(n152), .ZN(
        n154) );
  AOI21D1BWP30P140LVT U188 ( .A1(n286), .A2(i_data_bus[252]), .B(n154), .ZN(
        n156) );
  ND2D1BWP30P140LVT U189 ( .A1(n169), .A2(i_data_bus[28]), .ZN(n155) );
  ND4D1BWP30P140LVT U190 ( .A1(n158), .A2(n157), .A3(n156), .A4(n155), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U191 ( .A1(n279), .A2(i_data_bus[91]), .B1(n174), .B2(
        i_data_bus[59]), .ZN(n165) );
  AOI22D1BWP30P140LVT U192 ( .A1(n2), .A2(i_data_bus[123]), .B1(n280), .B2(
        i_data_bus[155]), .ZN(n164) );
  INVD1BWP30P140LVT U193 ( .I(i_data_bus[219]), .ZN(n160) );
  INVD1BWP30P140LVT U194 ( .I(i_data_bus[187]), .ZN(n159) );
  OAI22D1BWP30P140LVT U195 ( .A1(n177), .A2(n160), .B1(n244), .B2(n159), .ZN(
        n161) );
  AOI21D1BWP30P140LVT U196 ( .A1(n274), .A2(i_data_bus[251]), .B(n161), .ZN(
        n163) );
  ND2D1BWP30P140LVT U197 ( .A1(n169), .A2(i_data_bus[27]), .ZN(n162) );
  ND4D1BWP30P140LVT U198 ( .A1(n165), .A2(n164), .A3(n163), .A4(n162), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U199 ( .A1(n279), .A2(i_data_bus[90]), .B1(n174), .B2(
        i_data_bus[58]), .ZN(n173) );
  AOI22D1BWP30P140LVT U200 ( .A1(n2), .A2(i_data_bus[122]), .B1(n280), .B2(
        i_data_bus[154]), .ZN(n172) );
  INVD1BWP30P140LVT U201 ( .I(i_data_bus[218]), .ZN(n167) );
  INVD1BWP30P140LVT U202 ( .I(i_data_bus[186]), .ZN(n166) );
  OAI22D1BWP30P140LVT U203 ( .A1(n177), .A2(n167), .B1(n244), .B2(n166), .ZN(
        n168) );
  AOI21D1BWP30P140LVT U204 ( .A1(n274), .A2(i_data_bus[250]), .B(n168), .ZN(
        n171) );
  ND2D1BWP30P140LVT U205 ( .A1(n169), .A2(i_data_bus[26]), .ZN(n170) );
  ND4D1BWP30P140LVT U206 ( .A1(n173), .A2(n172), .A3(n171), .A4(n170), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U207 ( .A1(n279), .A2(i_data_bus[89]), .B1(n174), .B2(
        i_data_bus[57]), .ZN(n183) );
  AOI22D1BWP30P140LVT U208 ( .A1(n2), .A2(i_data_bus[121]), .B1(n280), .B2(
        i_data_bus[153]), .ZN(n182) );
  INVD1BWP30P140LVT U209 ( .I(i_data_bus[217]), .ZN(n176) );
  INVD1BWP30P140LVT U210 ( .I(i_data_bus[185]), .ZN(n175) );
  OAI22D1BWP30P140LVT U211 ( .A1(n177), .A2(n176), .B1(n244), .B2(n175), .ZN(
        n178) );
  AOI21D1BWP30P140LVT U212 ( .A1(n274), .A2(i_data_bus[249]), .B(n178), .ZN(
        n181) );
  INVD2BWP30P140LVT U213 ( .I(n179), .ZN(n287) );
  ND2D1BWP30P140LVT U214 ( .A1(n287), .A2(i_data_bus[25]), .ZN(n180) );
  ND4D1BWP30P140LVT U215 ( .A1(n183), .A2(n182), .A3(n181), .A4(n180), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U216 ( .A1(n279), .A2(i_data_bus[88]), .B1(n262), .B2(
        i_data_bus[56]), .ZN(n190) );
  AOI22D1BWP30P140LVT U217 ( .A1(n2), .A2(i_data_bus[120]), .B1(n280), .B2(
        i_data_bus[152]), .ZN(n189) );
  INVD1BWP30P140LVT U218 ( .I(i_data_bus[216]), .ZN(n185) );
  INVD1BWP30P140LVT U219 ( .I(i_data_bus[184]), .ZN(n184) );
  OAI22D1BWP30P140LVT U220 ( .A1(n284), .A2(n185), .B1(n244), .B2(n184), .ZN(
        n186) );
  AOI21D1BWP30P140LVT U221 ( .A1(n274), .A2(i_data_bus[248]), .B(n186), .ZN(
        n188) );
  ND2D1BWP30P140LVT U222 ( .A1(n287), .A2(i_data_bus[24]), .ZN(n187) );
  ND4D1BWP30P140LVT U223 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U224 ( .A1(n279), .A2(i_data_bus[87]), .B1(n262), .B2(
        i_data_bus[55]), .ZN(n197) );
  AOI22D1BWP30P140LVT U225 ( .A1(n2), .A2(i_data_bus[119]), .B1(n280), .B2(
        i_data_bus[151]), .ZN(n196) );
  INVD1BWP30P140LVT U226 ( .I(i_data_bus[215]), .ZN(n192) );
  INVD1BWP30P140LVT U227 ( .I(i_data_bus[183]), .ZN(n191) );
  OAI22D1BWP30P140LVT U228 ( .A1(n284), .A2(n192), .B1(n244), .B2(n191), .ZN(
        n193) );
  AOI21D1BWP30P140LVT U229 ( .A1(n274), .A2(i_data_bus[247]), .B(n193), .ZN(
        n195) );
  ND2D1BWP30P140LVT U230 ( .A1(n287), .A2(i_data_bus[23]), .ZN(n194) );
  ND4D1BWP30P140LVT U231 ( .A1(n197), .A2(n196), .A3(n195), .A4(n194), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U232 ( .A1(n279), .A2(i_data_bus[86]), .B1(n174), .B2(
        i_data_bus[54]), .ZN(n204) );
  AOI22D1BWP30P140LVT U233 ( .A1(n2), .A2(i_data_bus[118]), .B1(n280), .B2(
        i_data_bus[150]), .ZN(n203) );
  INVD1BWP30P140LVT U234 ( .I(i_data_bus[214]), .ZN(n199) );
  INVD1BWP30P140LVT U235 ( .I(i_data_bus[182]), .ZN(n198) );
  OAI22D1BWP30P140LVT U236 ( .A1(n284), .A2(n199), .B1(n244), .B2(n198), .ZN(
        n200) );
  AOI21D1BWP30P140LVT U237 ( .A1(n274), .A2(i_data_bus[246]), .B(n200), .ZN(
        n202) );
  ND2D1BWP30P140LVT U238 ( .A1(n287), .A2(i_data_bus[22]), .ZN(n201) );
  ND4D1BWP30P140LVT U239 ( .A1(n204), .A2(n203), .A3(n202), .A4(n201), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U240 ( .A1(n279), .A2(i_data_bus[85]), .B1(n262), .B2(
        i_data_bus[53]), .ZN(n211) );
  AOI22D1BWP30P140LVT U241 ( .A1(n2), .A2(i_data_bus[117]), .B1(n280), .B2(
        i_data_bus[149]), .ZN(n210) );
  INVD1BWP30P140LVT U242 ( .I(i_data_bus[213]), .ZN(n206) );
  INVD1BWP30P140LVT U243 ( .I(i_data_bus[181]), .ZN(n205) );
  OAI22D1BWP30P140LVT U244 ( .A1(n284), .A2(n206), .B1(n244), .B2(n205), .ZN(
        n207) );
  AOI21D1BWP30P140LVT U245 ( .A1(n274), .A2(i_data_bus[245]), .B(n207), .ZN(
        n209) );
  ND2D1BWP30P140LVT U246 ( .A1(n287), .A2(i_data_bus[21]), .ZN(n208) );
  ND4D1BWP30P140LVT U247 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U248 ( .A1(n279), .A2(i_data_bus[84]), .B1(n262), .B2(
        i_data_bus[52]), .ZN(n218) );
  AOI22D1BWP30P140LVT U249 ( .A1(n2), .A2(i_data_bus[116]), .B1(n280), .B2(
        i_data_bus[148]), .ZN(n217) );
  INVD1BWP30P140LVT U250 ( .I(i_data_bus[212]), .ZN(n213) );
  INVD1BWP30P140LVT U251 ( .I(i_data_bus[180]), .ZN(n212) );
  OAI22D1BWP30P140LVT U252 ( .A1(n284), .A2(n213), .B1(n244), .B2(n212), .ZN(
        n214) );
  AOI21D1BWP30P140LVT U253 ( .A1(n274), .A2(i_data_bus[244]), .B(n214), .ZN(
        n216) );
  ND2D1BWP30P140LVT U254 ( .A1(n287), .A2(i_data_bus[20]), .ZN(n215) );
  ND4D1BWP30P140LVT U255 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U256 ( .A1(n279), .A2(i_data_bus[83]), .B1(n174), .B2(
        i_data_bus[51]), .ZN(n224) );
  AOI22D1BWP30P140LVT U257 ( .A1(n2), .A2(i_data_bus[115]), .B1(n280), .B2(
        i_data_bus[147]), .ZN(n223) );
  INVD1BWP30P140LVT U258 ( .I(i_data_bus[179]), .ZN(n219) );
  MOAI22D1BWP30P140LVT U259 ( .A1(n244), .A2(n219), .B1(n271), .B2(
        i_data_bus[211]), .ZN(n220) );
  AOI21D1BWP30P140LVT U260 ( .A1(n274), .A2(i_data_bus[243]), .B(n220), .ZN(
        n222) );
  ND2D1BWP30P140LVT U261 ( .A1(n287), .A2(i_data_bus[19]), .ZN(n221) );
  ND4D1BWP30P140LVT U262 ( .A1(n224), .A2(n223), .A3(n222), .A4(n221), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U263 ( .A1(n279), .A2(i_data_bus[82]), .B1(n262), .B2(
        i_data_bus[50]), .ZN(n230) );
  AOI22D1BWP30P140LVT U264 ( .A1(n2), .A2(i_data_bus[114]), .B1(n280), .B2(
        i_data_bus[146]), .ZN(n229) );
  INVD1BWP30P140LVT U265 ( .I(i_data_bus[178]), .ZN(n225) );
  MOAI22D1BWP30P140LVT U266 ( .A1(n244), .A2(n225), .B1(n271), .B2(
        i_data_bus[210]), .ZN(n226) );
  AOI21D1BWP30P140LVT U267 ( .A1(n274), .A2(i_data_bus[242]), .B(n226), .ZN(
        n228) );
  ND2D1BWP30P140LVT U268 ( .A1(n287), .A2(i_data_bus[18]), .ZN(n227) );
  ND4D1BWP30P140LVT U269 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U270 ( .A1(n279), .A2(i_data_bus[81]), .B1(n262), .B2(
        i_data_bus[49]), .ZN(n236) );
  AOI22D1BWP30P140LVT U271 ( .A1(n2), .A2(i_data_bus[113]), .B1(n280), .B2(
        i_data_bus[145]), .ZN(n235) );
  INVD1BWP30P140LVT U272 ( .I(i_data_bus[177]), .ZN(n231) );
  MOAI22D1BWP30P140LVT U273 ( .A1(n244), .A2(n231), .B1(n271), .B2(
        i_data_bus[209]), .ZN(n232) );
  AOI21D1BWP30P140LVT U274 ( .A1(n274), .A2(i_data_bus[241]), .B(n232), .ZN(
        n234) );
  ND2D1BWP30P140LVT U275 ( .A1(n287), .A2(i_data_bus[17]), .ZN(n233) );
  ND4D1BWP30P140LVT U276 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U277 ( .A1(n279), .A2(i_data_bus[80]), .B1(n174), .B2(
        i_data_bus[48]), .ZN(n242) );
  AOI22D1BWP30P140LVT U278 ( .A1(n2), .A2(i_data_bus[112]), .B1(n280), .B2(
        i_data_bus[144]), .ZN(n241) );
  INVD1BWP30P140LVT U279 ( .I(i_data_bus[176]), .ZN(n237) );
  MOAI22D1BWP30P140LVT U280 ( .A1(n244), .A2(n237), .B1(n271), .B2(
        i_data_bus[208]), .ZN(n238) );
  AOI21D1BWP30P140LVT U281 ( .A1(n274), .A2(i_data_bus[240]), .B(n238), .ZN(
        n240) );
  ND2D1BWP30P140LVT U282 ( .A1(n287), .A2(i_data_bus[16]), .ZN(n239) );
  ND4D1BWP30P140LVT U283 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U284 ( .A1(n279), .A2(i_data_bus[79]), .B1(n262), .B2(
        i_data_bus[47]), .ZN(n249) );
  AOI22D1BWP30P140LVT U285 ( .A1(n2), .A2(i_data_bus[111]), .B1(n280), .B2(
        i_data_bus[143]), .ZN(n248) );
  INVD1BWP30P140LVT U286 ( .I(i_data_bus[175]), .ZN(n243) );
  MOAI22D1BWP30P140LVT U287 ( .A1(n244), .A2(n243), .B1(n271), .B2(
        i_data_bus[207]), .ZN(n245) );
  AOI21D1BWP30P140LVT U288 ( .A1(n274), .A2(i_data_bus[239]), .B(n245), .ZN(
        n247) );
  ND2D1BWP30P140LVT U289 ( .A1(n287), .A2(i_data_bus[15]), .ZN(n246) );
  ND4D1BWP30P140LVT U290 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U291 ( .A1(n263), .A2(i_data_bus[64]), .B1(n262), .B2(
        i_data_bus[32]), .ZN(n255) );
  AOI22D1BWP30P140LVT U292 ( .A1(n2), .A2(i_data_bus[96]), .B1(n280), .B2(
        i_data_bus[128]), .ZN(n254) );
  INR2D1BWP30P140LVT U293 ( .A1(i_data_bus[192]), .B1(n284), .ZN(n251) );
  INR2D1BWP30P140LVT U294 ( .A1(i_data_bus[160]), .B1(n282), .ZN(n250) );
  AOI211D1BWP30P140LVT U295 ( .A1(i_data_bus[224]), .A2(n286), .B(n251), .C(
        n250), .ZN(n253) );
  ND2D1BWP30P140LVT U296 ( .A1(n266), .A2(i_data_bus[0]), .ZN(n252) );
  ND4D1BWP30P140LVT U297 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U298 ( .A1(n263), .A2(i_data_bus[66]), .B1(n262), .B2(
        i_data_bus[34]), .ZN(n261) );
  AOI22D1BWP30P140LVT U299 ( .A1(n2), .A2(i_data_bus[98]), .B1(n280), .B2(
        i_data_bus[130]), .ZN(n260) );
  INVD1BWP30P140LVT U300 ( .I(i_data_bus[162]), .ZN(n256) );
  MOAI22D1BWP30P140LVT U301 ( .A1(n282), .A2(n256), .B1(n271), .B2(
        i_data_bus[194]), .ZN(n257) );
  AOI21D1BWP30P140LVT U302 ( .A1(n286), .A2(i_data_bus[226]), .B(n257), .ZN(
        n259) );
  ND2D1BWP30P140LVT U303 ( .A1(n266), .A2(i_data_bus[2]), .ZN(n258) );
  ND4D1BWP30P140LVT U304 ( .A1(n261), .A2(n260), .A3(n259), .A4(n258), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U305 ( .A1(n263), .A2(i_data_bus[65]), .B1(n262), .B2(
        i_data_bus[33]), .ZN(n270) );
  AOI22D1BWP30P140LVT U306 ( .A1(n2), .A2(i_data_bus[97]), .B1(n280), .B2(
        i_data_bus[129]), .ZN(n269) );
  INVD1BWP30P140LVT U307 ( .I(i_data_bus[161]), .ZN(n264) );
  MOAI22D1BWP30P140LVT U308 ( .A1(n282), .A2(n264), .B1(n271), .B2(
        i_data_bus[193]), .ZN(n265) );
  AOI21D1BWP30P140LVT U309 ( .A1(n286), .A2(i_data_bus[225]), .B(n265), .ZN(
        n268) );
  ND2D1BWP30P140LVT U310 ( .A1(n266), .A2(i_data_bus[1]), .ZN(n267) );
  ND4D1BWP30P140LVT U311 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U312 ( .A1(n279), .A2(i_data_bus[78]), .B1(n262), .B2(
        i_data_bus[46]), .ZN(n278) );
  AOI22D1BWP30P140LVT U313 ( .A1(n2), .A2(i_data_bus[110]), .B1(n280), .B2(
        i_data_bus[142]), .ZN(n277) );
  INVD1BWP30P140LVT U314 ( .I(i_data_bus[174]), .ZN(n272) );
  MOAI22D1BWP30P140LVT U315 ( .A1(n282), .A2(n272), .B1(n271), .B2(
        i_data_bus[206]), .ZN(n273) );
  AOI21D1BWP30P140LVT U316 ( .A1(n274), .A2(i_data_bus[238]), .B(n273), .ZN(
        n276) );
  ND2D1BWP30P140LVT U317 ( .A1(n287), .A2(i_data_bus[14]), .ZN(n275) );
  ND4D1BWP30P140LVT U318 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U319 ( .A1(n279), .A2(i_data_bus[77]), .B1(n174), .B2(
        i_data_bus[45]), .ZN(n291) );
  AOI22D1BWP30P140LVT U320 ( .A1(n2), .A2(i_data_bus[109]), .B1(n280), .B2(
        i_data_bus[141]), .ZN(n290) );
  INVD1BWP30P140LVT U321 ( .I(i_data_bus[205]), .ZN(n283) );
  INVD1BWP30P140LVT U322 ( .I(i_data_bus[173]), .ZN(n281) );
  OAI22D1BWP30P140LVT U323 ( .A1(n284), .A2(n283), .B1(n282), .B2(n281), .ZN(
        n285) );
  AOI21D1BWP30P140LVT U324 ( .A1(n286), .A2(i_data_bus[237]), .B(n285), .ZN(
        n289) );
  ND2D1BWP30P140LVT U325 ( .A1(n287), .A2(i_data_bus[13]), .ZN(n288) );
  ND4D1BWP30P140LVT U326 ( .A1(n291), .A2(n290), .A3(n289), .A4(n288), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_2 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n165), .ZN(n270) );
  INVD1BWP30P140LVT U4 ( .I(n166), .ZN(n47) );
  CKND2D3BWP30P140LVT U5 ( .A1(n21), .A2(n23), .ZN(n169) );
  NR2OPTPAD2BWP30P140LVT U6 ( .A1(n15), .A2(n14), .ZN(n23) );
  INVD1BWP30P140LVT U7 ( .I(n169), .ZN(n1) );
  INVD4BWP30P140LVT U8 ( .I(n47), .ZN(n2) );
  INVD3BWP30P140LVT U9 ( .I(n167), .ZN(n3) );
  ND2OPTPAD2BWP30P140LVT U10 ( .A1(n10), .A2(n9), .ZN(n15) );
  NR2OPTPAD2BWP30P140LVT U11 ( .A1(n20), .A2(i_cmd[5]), .ZN(n30) );
  INVD2BWP30P140LVT U12 ( .I(n262), .ZN(n275) );
  INVD3BWP30P140LVT U13 ( .I(n168), .ZN(n254) );
  NR2D1BWP30P140LVT U14 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n17) );
  INVD4BWP30P140LVT U15 ( .I(n168), .ZN(n271) );
  ND2OPTIBD1BWP30P140LVT U16 ( .A1(n13), .A2(n12), .ZN(n14) );
  INVD2BWP30P140LVT U17 ( .I(n1), .ZN(n159) );
  INVD1BWP30P140LVT U18 ( .I(n37), .ZN(n168) );
  ND2D1BWP30P140LVT U19 ( .A1(n17), .A2(n16), .ZN(n18) );
  IND2D2BWP30P140LVT U20 ( .A1(n41), .B1(n33), .ZN(n167) );
  INVD1BWP30P140LVT U21 ( .I(n8), .ZN(n175) );
  INR2D1BWP30P140LVT U22 ( .A1(n44), .B1(n41), .ZN(n166) );
  OR2D1BWP30P140LVT U23 ( .A1(n41), .A2(n40), .Z(n165) );
  INVD1BWP30P140LVT U24 ( .I(n26), .ZN(n76) );
  ND3D1BWP30P140LVT U25 ( .A1(n30), .A2(n29), .A3(n28), .ZN(n41) );
  INVD1BWP30P140LVT U26 ( .I(i_cmd[0]), .ZN(n9) );
  INR3D0BWP30P140LVT U27 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n9), .ZN(n7) );
  OR2D4BWP30P140LVT U28 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n20) );
  INVD1BWP30P140LVT U29 ( .I(rst), .ZN(n4) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n4), .A2(i_en), .Z(n11) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n30), .A2(n11), .Z(n6) );
  OR2D1BWP30P140LVT U32 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n43) );
  NR2D1BWP30P140LVT U33 ( .A1(n43), .A2(i_cmd[1]), .ZN(n5) );
  ND2OPTIBD1BWP30P140LVT U34 ( .A1(n6), .A2(n5), .ZN(n35) );
  INR2D1BWP30P140LVT U35 ( .A1(n7), .B1(n35), .ZN(n8) );
  OR2D4BWP30P140LVT U36 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n32) );
  INVD2BWP30P140LVT U37 ( .I(n32), .ZN(n10) );
  INVD1BWP30P140LVT U38 ( .I(i_cmd[3]), .ZN(n13) );
  INVD1BWP30P140LVT U39 ( .I(n11), .ZN(n27) );
  NR2D1BWP30P140LVT U40 ( .A1(i_cmd[4]), .A2(n27), .ZN(n12) );
  CKAN2D1BWP30P140LVT U41 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n16) );
  INR2D4BWP30P140LVT U42 ( .A1(n23), .B1(n18), .ZN(n262) );
  ND2D1BWP30P140LVT U43 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n19) );
  NR2D1BWP30P140LVT U44 ( .A1(n20), .A2(n19), .ZN(n21) );
  INVD1BWP30P140LVT U45 ( .I(i_cmd[7]), .ZN(n22) );
  INR4D0BWP30P140LVT U46 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n22), .ZN(n25) );
  INVD1BWP30P140LVT U47 ( .I(n23), .ZN(n24) );
  INR2D1BWP30P140LVT U48 ( .A1(n25), .B1(n24), .ZN(n26) );
  INVD2BWP30P140LVT U49 ( .I(n76), .ZN(n277) );
  NR4D0BWP30P140LVT U50 ( .A1(n278), .A2(n262), .A3(n1), .A4(n277), .ZN(n46)
         );
  NR2D1BWP30P140LVT U51 ( .A1(i_cmd[0]), .A2(n27), .ZN(n29) );
  INVD1BWP30P140LVT U52 ( .I(i_cmd[4]), .ZN(n28) );
  ND2D1BWP30P140LVT U53 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n31) );
  NR2D1BWP30P140LVT U54 ( .A1(n32), .A2(n31), .ZN(n33) );
  ND2D1BWP30P140LVT U55 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n34) );
  NR2D1BWP30P140LVT U56 ( .A1(n34), .A2(i_cmd[0]), .ZN(n36) );
  INR2D1BWP30P140LVT U57 ( .A1(n36), .B1(n35), .ZN(n37) );
  NR2D1BWP30P140LVT U58 ( .A1(n3), .A2(n271), .ZN(n45) );
  INVD1BWP30P140LVT U59 ( .I(i_cmd[2]), .ZN(n39) );
  NR2D1BWP30P140LVT U60 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .ZN(n38) );
  IND3D1BWP30P140LVT U61 ( .A1(n39), .B1(n38), .B2(i_valid[2]), .ZN(n40) );
  ND2D1BWP30P140LVT U62 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n42) );
  NR2D1BWP30P140LVT U63 ( .A1(n43), .A2(n42), .ZN(n44) );
  ND4D1BWP30P140LVT U64 ( .A1(n46), .A2(n45), .A3(n165), .A4(n47), .ZN(N402)
         );
  AOI22D1BWP30P140LVT U65 ( .A1(n270), .A2(i_data_bus[95]), .B1(n2), .B2(
        i_data_bus[63]), .ZN(n54) );
  AOI22D1BWP30P140LVT U66 ( .A1(n3), .A2(i_data_bus[127]), .B1(n271), .B2(
        i_data_bus[159]), .ZN(n53) );
  INVD2BWP30P140LVT U67 ( .I(n262), .ZN(n172) );
  INVD1BWP30P140LVT U68 ( .I(i_data_bus[223]), .ZN(n49) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[191]), .ZN(n48) );
  OAI22D1BWP30P140LVT U70 ( .A1(n172), .A2(n49), .B1(n169), .B2(n48), .ZN(n50)
         );
  AOI21D1BWP30P140LVT U71 ( .A1(n277), .A2(i_data_bus[255]), .B(n50), .ZN(n52)
         );
  ND2D1BWP30P140LVT U72 ( .A1(n257), .A2(i_data_bus[31]), .ZN(n51) );
  ND4D1BWP30P140LVT U73 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(N400) );
  AOI22D1BWP30P140LVT U74 ( .A1(n270), .A2(i_data_bus[94]), .B1(n2), .B2(
        i_data_bus[62]), .ZN(n61) );
  AOI22D1BWP30P140LVT U75 ( .A1(n3), .A2(i_data_bus[126]), .B1(n271), .B2(
        i_data_bus[158]), .ZN(n60) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[222]), .ZN(n56) );
  INVD1BWP30P140LVT U77 ( .I(i_data_bus[190]), .ZN(n55) );
  OAI22D1BWP30P140LVT U78 ( .A1(n172), .A2(n56), .B1(n169), .B2(n55), .ZN(n57)
         );
  AOI21D1BWP30P140LVT U79 ( .A1(n265), .A2(i_data_bus[254]), .B(n57), .ZN(n59)
         );
  ND2D1BWP30P140LVT U80 ( .A1(n278), .A2(i_data_bus[30]), .ZN(n58) );
  ND4D1BWP30P140LVT U81 ( .A1(n61), .A2(n60), .A3(n59), .A4(n58), .ZN(N399) );
  AOI22D1BWP30P140LVT U82 ( .A1(n270), .A2(i_data_bus[93]), .B1(n2), .B2(
        i_data_bus[61]), .ZN(n68) );
  AOI22D1BWP30P140LVT U83 ( .A1(n3), .A2(i_data_bus[125]), .B1(n271), .B2(
        i_data_bus[157]), .ZN(n67) );
  INVD1BWP30P140LVT U84 ( .I(i_data_bus[221]), .ZN(n63) );
  INVD1BWP30P140LVT U85 ( .I(i_data_bus[189]), .ZN(n62) );
  OAI22D1BWP30P140LVT U86 ( .A1(n172), .A2(n63), .B1(n159), .B2(n62), .ZN(n64)
         );
  AOI21D1BWP30P140LVT U87 ( .A1(n265), .A2(i_data_bus[253]), .B(n64), .ZN(n66)
         );
  ND2D1BWP30P140LVT U88 ( .A1(n257), .A2(i_data_bus[29]), .ZN(n65) );
  ND4D1BWP30P140LVT U89 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(N398) );
  AOI22D1BWP30P140LVT U90 ( .A1(n270), .A2(i_data_bus[92]), .B1(n2), .B2(
        i_data_bus[60]), .ZN(n75) );
  AOI22D1BWP30P140LVT U91 ( .A1(n3), .A2(i_data_bus[124]), .B1(n271), .B2(
        i_data_bus[156]), .ZN(n74) );
  INVD1BWP30P140LVT U92 ( .I(i_data_bus[220]), .ZN(n70) );
  INVD1BWP30P140LVT U93 ( .I(i_data_bus[188]), .ZN(n69) );
  OAI22D1BWP30P140LVT U94 ( .A1(n172), .A2(n70), .B1(n159), .B2(n69), .ZN(n71)
         );
  AOI21D1BWP30P140LVT U95 ( .A1(n265), .A2(i_data_bus[252]), .B(n71), .ZN(n73)
         );
  ND2D1BWP30P140LVT U96 ( .A1(n278), .A2(i_data_bus[28]), .ZN(n72) );
  ND4D1BWP30P140LVT U97 ( .A1(n75), .A2(n74), .A3(n73), .A4(n72), .ZN(N397) );
  AOI22D1BWP30P140LVT U98 ( .A1(n270), .A2(i_data_bus[91]), .B1(n2), .B2(
        i_data_bus[59]), .ZN(n83) );
  AOI22D1BWP30P140LVT U99 ( .A1(n3), .A2(i_data_bus[123]), .B1(n271), .B2(
        i_data_bus[155]), .ZN(n82) );
  INVD2BWP30P140LVT U100 ( .I(n76), .ZN(n265) );
  INVD1BWP30P140LVT U101 ( .I(i_data_bus[219]), .ZN(n78) );
  INVD1BWP30P140LVT U102 ( .I(i_data_bus[187]), .ZN(n77) );
  OAI22D1BWP30P140LVT U103 ( .A1(n172), .A2(n78), .B1(n159), .B2(n77), .ZN(n79) );
  AOI21D1BWP30P140LVT U104 ( .A1(n265), .A2(i_data_bus[251]), .B(n79), .ZN(n81) );
  ND2D1BWP30P140LVT U105 ( .A1(n257), .A2(i_data_bus[27]), .ZN(n80) );
  ND4D1BWP30P140LVT U106 ( .A1(n83), .A2(n82), .A3(n81), .A4(n80), .ZN(N396)
         );
  AOI22D1BWP30P140LVT U107 ( .A1(n270), .A2(i_data_bus[90]), .B1(n2), .B2(
        i_data_bus[58]), .ZN(n90) );
  AOI22D1BWP30P140LVT U108 ( .A1(n3), .A2(i_data_bus[122]), .B1(n271), .B2(
        i_data_bus[154]), .ZN(n89) );
  INVD1BWP30P140LVT U109 ( .I(i_data_bus[218]), .ZN(n85) );
  INVD1BWP30P140LVT U110 ( .I(i_data_bus[186]), .ZN(n84) );
  OAI22D1BWP30P140LVT U111 ( .A1(n172), .A2(n85), .B1(n159), .B2(n84), .ZN(n86) );
  AOI21D1BWP30P140LVT U112 ( .A1(n265), .A2(i_data_bus[250]), .B(n86), .ZN(n88) );
  ND2D1BWP30P140LVT U113 ( .A1(n8), .A2(i_data_bus[26]), .ZN(n87) );
  ND4D1BWP30P140LVT U114 ( .A1(n90), .A2(n89), .A3(n88), .A4(n87), .ZN(N395)
         );
  AOI22D1BWP30P140LVT U115 ( .A1(n270), .A2(i_data_bus[89]), .B1(n2), .B2(
        i_data_bus[57]), .ZN(n97) );
  AOI22D1BWP30P140LVT U116 ( .A1(n3), .A2(i_data_bus[121]), .B1(n271), .B2(
        i_data_bus[153]), .ZN(n96) );
  INVD1BWP30P140LVT U117 ( .I(i_data_bus[217]), .ZN(n92) );
  INVD1BWP30P140LVT U118 ( .I(i_data_bus[185]), .ZN(n91) );
  OAI22D1BWP30P140LVT U119 ( .A1(n172), .A2(n92), .B1(n159), .B2(n91), .ZN(n93) );
  AOI21D1BWP30P140LVT U120 ( .A1(n265), .A2(i_data_bus[249]), .B(n93), .ZN(n95) );
  INVD2BWP30P140LVT U121 ( .I(n175), .ZN(n278) );
  ND2D1BWP30P140LVT U122 ( .A1(n278), .A2(i_data_bus[25]), .ZN(n94) );
  ND4D1BWP30P140LVT U123 ( .A1(n97), .A2(n96), .A3(n95), .A4(n94), .ZN(N394)
         );
  AOI22D1BWP30P140LVT U124 ( .A1(n270), .A2(i_data_bus[88]), .B1(n2), .B2(
        i_data_bus[56]), .ZN(n104) );
  AOI22D1BWP30P140LVT U125 ( .A1(n3), .A2(i_data_bus[120]), .B1(n271), .B2(
        i_data_bus[152]), .ZN(n103) );
  INVD1BWP30P140LVT U126 ( .I(i_data_bus[216]), .ZN(n99) );
  INVD1BWP30P140LVT U127 ( .I(i_data_bus[184]), .ZN(n98) );
  OAI22D1BWP30P140LVT U128 ( .A1(n275), .A2(n99), .B1(n159), .B2(n98), .ZN(
        n100) );
  AOI21D1BWP30P140LVT U129 ( .A1(n265), .A2(i_data_bus[248]), .B(n100), .ZN(
        n102) );
  ND2D1BWP30P140LVT U130 ( .A1(n278), .A2(i_data_bus[24]), .ZN(n101) );
  ND4D1BWP30P140LVT U131 ( .A1(n104), .A2(n103), .A3(n102), .A4(n101), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U132 ( .A1(n270), .A2(i_data_bus[87]), .B1(n2), .B2(
        i_data_bus[55]), .ZN(n111) );
  AOI22D1BWP30P140LVT U133 ( .A1(n3), .A2(i_data_bus[119]), .B1(n271), .B2(
        i_data_bus[151]), .ZN(n110) );
  INVD1BWP30P140LVT U134 ( .I(i_data_bus[215]), .ZN(n106) );
  INVD1BWP30P140LVT U135 ( .I(i_data_bus[183]), .ZN(n105) );
  OAI22D1BWP30P140LVT U136 ( .A1(n275), .A2(n106), .B1(n159), .B2(n105), .ZN(
        n107) );
  AOI21D1BWP30P140LVT U137 ( .A1(n265), .A2(i_data_bus[247]), .B(n107), .ZN(
        n109) );
  ND2D1BWP30P140LVT U138 ( .A1(n278), .A2(i_data_bus[23]), .ZN(n108) );
  ND4D1BWP30P140LVT U139 ( .A1(n111), .A2(n110), .A3(n109), .A4(n108), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U140 ( .A1(n270), .A2(i_data_bus[86]), .B1(n2), .B2(
        i_data_bus[54]), .ZN(n118) );
  AOI22D1BWP30P140LVT U141 ( .A1(n3), .A2(i_data_bus[118]), .B1(n271), .B2(
        i_data_bus[150]), .ZN(n117) );
  INVD1BWP30P140LVT U142 ( .I(i_data_bus[214]), .ZN(n113) );
  INVD1BWP30P140LVT U143 ( .I(i_data_bus[182]), .ZN(n112) );
  OAI22D1BWP30P140LVT U144 ( .A1(n275), .A2(n113), .B1(n159), .B2(n112), .ZN(
        n114) );
  AOI21D1BWP30P140LVT U145 ( .A1(n265), .A2(i_data_bus[246]), .B(n114), .ZN(
        n116) );
  ND2D1BWP30P140LVT U146 ( .A1(n278), .A2(i_data_bus[22]), .ZN(n115) );
  ND4D1BWP30P140LVT U147 ( .A1(n118), .A2(n117), .A3(n116), .A4(n115), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U148 ( .A1(n270), .A2(i_data_bus[85]), .B1(n2), .B2(
        i_data_bus[53]), .ZN(n125) );
  AOI22D1BWP30P140LVT U149 ( .A1(n3), .A2(i_data_bus[117]), .B1(n271), .B2(
        i_data_bus[149]), .ZN(n124) );
  INVD1BWP30P140LVT U150 ( .I(i_data_bus[213]), .ZN(n120) );
  INVD1BWP30P140LVT U151 ( .I(i_data_bus[181]), .ZN(n119) );
  OAI22D1BWP30P140LVT U152 ( .A1(n275), .A2(n120), .B1(n159), .B2(n119), .ZN(
        n121) );
  AOI21D1BWP30P140LVT U153 ( .A1(n265), .A2(i_data_bus[245]), .B(n121), .ZN(
        n123) );
  ND2D1BWP30P140LVT U154 ( .A1(n278), .A2(i_data_bus[21]), .ZN(n122) );
  ND4D1BWP30P140LVT U155 ( .A1(n125), .A2(n124), .A3(n123), .A4(n122), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U156 ( .A1(n270), .A2(i_data_bus[84]), .B1(n2), .B2(
        i_data_bus[52]), .ZN(n132) );
  AOI22D1BWP30P140LVT U157 ( .A1(n3), .A2(i_data_bus[116]), .B1(n271), .B2(
        i_data_bus[148]), .ZN(n131) );
  INVD1BWP30P140LVT U158 ( .I(i_data_bus[212]), .ZN(n127) );
  INVD1BWP30P140LVT U159 ( .I(i_data_bus[180]), .ZN(n126) );
  OAI22D1BWP30P140LVT U160 ( .A1(n275), .A2(n127), .B1(n159), .B2(n126), .ZN(
        n128) );
  AOI21D1BWP30P140LVT U161 ( .A1(n265), .A2(i_data_bus[244]), .B(n128), .ZN(
        n130) );
  ND2D1BWP30P140LVT U162 ( .A1(n278), .A2(i_data_bus[20]), .ZN(n129) );
  ND4D1BWP30P140LVT U163 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U164 ( .A1(n270), .A2(i_data_bus[83]), .B1(n2), .B2(
        i_data_bus[51]), .ZN(n139) );
  AOI22D1BWP30P140LVT U165 ( .A1(n3), .A2(i_data_bus[115]), .B1(n271), .B2(
        i_data_bus[147]), .ZN(n138) );
  INVD1BWP30P140LVT U166 ( .I(i_data_bus[211]), .ZN(n134) );
  INVD1BWP30P140LVT U167 ( .I(i_data_bus[179]), .ZN(n133) );
  OAI22D1BWP30P140LVT U168 ( .A1(n275), .A2(n134), .B1(n159), .B2(n133), .ZN(
        n135) );
  AOI21D1BWP30P140LVT U169 ( .A1(n265), .A2(i_data_bus[243]), .B(n135), .ZN(
        n137) );
  ND2D1BWP30P140LVT U170 ( .A1(n278), .A2(i_data_bus[19]), .ZN(n136) );
  ND4D1BWP30P140LVT U171 ( .A1(n139), .A2(n138), .A3(n137), .A4(n136), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U172 ( .A1(n270), .A2(i_data_bus[82]), .B1(n2), .B2(
        i_data_bus[50]), .ZN(n145) );
  AOI22D1BWP30P140LVT U173 ( .A1(n3), .A2(i_data_bus[114]), .B1(n271), .B2(
        i_data_bus[146]), .ZN(n144) );
  INVD1BWP30P140LVT U174 ( .I(i_data_bus[178]), .ZN(n140) );
  MOAI22D1BWP30P140LVT U175 ( .A1(n159), .A2(n140), .B1(n262), .B2(
        i_data_bus[210]), .ZN(n141) );
  AOI21D1BWP30P140LVT U176 ( .A1(n265), .A2(i_data_bus[242]), .B(n141), .ZN(
        n143) );
  ND2D1BWP30P140LVT U177 ( .A1(n278), .A2(i_data_bus[18]), .ZN(n142) );
  ND4D1BWP30P140LVT U178 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U179 ( .A1(n270), .A2(i_data_bus[81]), .B1(n2), .B2(
        i_data_bus[49]), .ZN(n151) );
  AOI22D1BWP30P140LVT U180 ( .A1(n3), .A2(i_data_bus[113]), .B1(n271), .B2(
        i_data_bus[145]), .ZN(n150) );
  INVD1BWP30P140LVT U181 ( .I(i_data_bus[177]), .ZN(n146) );
  MOAI22D1BWP30P140LVT U182 ( .A1(n159), .A2(n146), .B1(n262), .B2(
        i_data_bus[209]), .ZN(n147) );
  AOI21D1BWP30P140LVT U183 ( .A1(n265), .A2(i_data_bus[241]), .B(n147), .ZN(
        n149) );
  ND2D1BWP30P140LVT U184 ( .A1(n278), .A2(i_data_bus[17]), .ZN(n148) );
  ND4D1BWP30P140LVT U185 ( .A1(n151), .A2(n150), .A3(n149), .A4(n148), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U186 ( .A1(n270), .A2(i_data_bus[80]), .B1(n2), .B2(
        i_data_bus[48]), .ZN(n157) );
  AOI22D1BWP30P140LVT U187 ( .A1(n3), .A2(i_data_bus[112]), .B1(n271), .B2(
        i_data_bus[144]), .ZN(n156) );
  INVD1BWP30P140LVT U188 ( .I(i_data_bus[176]), .ZN(n152) );
  MOAI22D1BWP30P140LVT U189 ( .A1(n159), .A2(n152), .B1(n262), .B2(
        i_data_bus[208]), .ZN(n153) );
  AOI21D1BWP30P140LVT U190 ( .A1(n265), .A2(i_data_bus[240]), .B(n153), .ZN(
        n155) );
  ND2D1BWP30P140LVT U191 ( .A1(n278), .A2(i_data_bus[16]), .ZN(n154) );
  ND4D1BWP30P140LVT U192 ( .A1(n157), .A2(n156), .A3(n155), .A4(n154), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U193 ( .A1(n270), .A2(i_data_bus[79]), .B1(n2), .B2(
        i_data_bus[47]), .ZN(n164) );
  AOI22D1BWP30P140LVT U194 ( .A1(n3), .A2(i_data_bus[111]), .B1(n271), .B2(
        i_data_bus[143]), .ZN(n163) );
  INVD1BWP30P140LVT U195 ( .I(i_data_bus[175]), .ZN(n158) );
  MOAI22D1BWP30P140LVT U196 ( .A1(n159), .A2(n158), .B1(n262), .B2(
        i_data_bus[207]), .ZN(n160) );
  AOI21D1BWP30P140LVT U197 ( .A1(n265), .A2(i_data_bus[239]), .B(n160), .ZN(
        n162) );
  ND2D1BWP30P140LVT U198 ( .A1(n278), .A2(i_data_bus[15]), .ZN(n161) );
  ND4D1BWP30P140LVT U199 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U200 ( .A1(n270), .A2(i_data_bus[72]), .B1(n2), .B2(
        i_data_bus[40]), .ZN(n179) );
  AOI22D1BWP30P140LVT U201 ( .A1(n3), .A2(i_data_bus[104]), .B1(n254), .B2(
        i_data_bus[136]), .ZN(n178) );
  INVD1BWP30P140LVT U202 ( .I(n169), .ZN(n170) );
  INVD2BWP30P140LVT U203 ( .I(n170), .ZN(n273) );
  INVD1BWP30P140LVT U204 ( .I(i_data_bus[168]), .ZN(n173) );
  INVD1BWP30P140LVT U205 ( .I(i_data_bus[200]), .ZN(n171) );
  OAI22D1BWP30P140LVT U206 ( .A1(n273), .A2(n173), .B1(n172), .B2(n171), .ZN(
        n174) );
  AOI21D1BWP30P140LVT U207 ( .A1(n265), .A2(i_data_bus[232]), .B(n174), .ZN(
        n177) );
  INVD2BWP30P140LVT U208 ( .I(n175), .ZN(n257) );
  ND2D1BWP30P140LVT U209 ( .A1(n257), .A2(i_data_bus[8]), .ZN(n176) );
  ND4D1BWP30P140LVT U210 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U211 ( .A1(n270), .A2(i_data_bus[76]), .B1(n2), .B2(
        i_data_bus[44]), .ZN(n186) );
  AOI22D1BWP30P140LVT U212 ( .A1(n3), .A2(i_data_bus[108]), .B1(n254), .B2(
        i_data_bus[140]), .ZN(n185) );
  INVD1BWP30P140LVT U213 ( .I(i_data_bus[204]), .ZN(n181) );
  INVD1BWP30P140LVT U214 ( .I(i_data_bus[172]), .ZN(n180) );
  OAI22D1BWP30P140LVT U215 ( .A1(n275), .A2(n181), .B1(n273), .B2(n180), .ZN(
        n182) );
  AOI21D1BWP30P140LVT U216 ( .A1(n277), .A2(i_data_bus[236]), .B(n182), .ZN(
        n184) );
  ND2D1BWP30P140LVT U217 ( .A1(n257), .A2(i_data_bus[12]), .ZN(n183) );
  ND4D1BWP30P140LVT U218 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(
        N381) );
  AOI22D1BWP30P140LVT U219 ( .A1(n270), .A2(i_data_bus[75]), .B1(n2), .B2(
        i_data_bus[43]), .ZN(n193) );
  AOI22D1BWP30P140LVT U220 ( .A1(n3), .A2(i_data_bus[107]), .B1(n254), .B2(
        i_data_bus[139]), .ZN(n192) );
  INVD1BWP30P140LVT U221 ( .I(i_data_bus[203]), .ZN(n188) );
  INVD1BWP30P140LVT U222 ( .I(i_data_bus[171]), .ZN(n187) );
  OAI22D1BWP30P140LVT U223 ( .A1(n275), .A2(n188), .B1(n273), .B2(n187), .ZN(
        n189) );
  AOI21D1BWP30P140LVT U224 ( .A1(n277), .A2(i_data_bus[235]), .B(n189), .ZN(
        n191) );
  ND2D1BWP30P140LVT U225 ( .A1(n257), .A2(i_data_bus[11]), .ZN(n190) );
  ND4D1BWP30P140LVT U226 ( .A1(n193), .A2(n192), .A3(n191), .A4(n190), .ZN(
        N380) );
  AOI22D1BWP30P140LVT U227 ( .A1(n270), .A2(i_data_bus[74]), .B1(n2), .B2(
        i_data_bus[42]), .ZN(n200) );
  AOI22D1BWP30P140LVT U228 ( .A1(n3), .A2(i_data_bus[106]), .B1(n254), .B2(
        i_data_bus[138]), .ZN(n199) );
  INVD1BWP30P140LVT U229 ( .I(i_data_bus[202]), .ZN(n195) );
  INVD1BWP30P140LVT U230 ( .I(i_data_bus[170]), .ZN(n194) );
  OAI22D1BWP30P140LVT U231 ( .A1(n275), .A2(n195), .B1(n273), .B2(n194), .ZN(
        n196) );
  AOI21D1BWP30P140LVT U232 ( .A1(n277), .A2(i_data_bus[234]), .B(n196), .ZN(
        n198) );
  ND2D1BWP30P140LVT U233 ( .A1(n257), .A2(i_data_bus[10]), .ZN(n197) );
  ND4D1BWP30P140LVT U234 ( .A1(n200), .A2(n199), .A3(n198), .A4(n197), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U235 ( .A1(n270), .A2(i_data_bus[73]), .B1(n2), .B2(
        i_data_bus[41]), .ZN(n207) );
  AOI22D1BWP30P140LVT U236 ( .A1(n3), .A2(i_data_bus[105]), .B1(n254), .B2(
        i_data_bus[137]), .ZN(n206) );
  INVD1BWP30P140LVT U237 ( .I(i_data_bus[201]), .ZN(n202) );
  INVD1BWP30P140LVT U238 ( .I(i_data_bus[169]), .ZN(n201) );
  OAI22D1BWP30P140LVT U239 ( .A1(n275), .A2(n202), .B1(n273), .B2(n201), .ZN(
        n203) );
  AOI21D1BWP30P140LVT U240 ( .A1(n277), .A2(i_data_bus[233]), .B(n203), .ZN(
        n205) );
  ND2D1BWP30P140LVT U241 ( .A1(n257), .A2(i_data_bus[9]), .ZN(n204) );
  ND4D1BWP30P140LVT U242 ( .A1(n207), .A2(n206), .A3(n205), .A4(n204), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U243 ( .A1(n270), .A2(i_data_bus[71]), .B1(n2), .B2(
        i_data_bus[39]), .ZN(n214) );
  AOI22D1BWP30P140LVT U244 ( .A1(n3), .A2(i_data_bus[103]), .B1(n254), .B2(
        i_data_bus[135]), .ZN(n213) );
  INVD1BWP30P140LVT U245 ( .I(i_data_bus[199]), .ZN(n209) );
  INVD1BWP30P140LVT U246 ( .I(i_data_bus[167]), .ZN(n208) );
  OAI22D1BWP30P140LVT U247 ( .A1(n275), .A2(n209), .B1(n273), .B2(n208), .ZN(
        n210) );
  AOI21D1BWP30P140LVT U248 ( .A1(n277), .A2(i_data_bus[231]), .B(n210), .ZN(
        n212) );
  ND2D1BWP30P140LVT U249 ( .A1(n257), .A2(i_data_bus[7]), .ZN(n211) );
  ND4D1BWP30P140LVT U250 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U251 ( .A1(n270), .A2(i_data_bus[70]), .B1(n2), .B2(
        i_data_bus[38]), .ZN(n221) );
  AOI22D1BWP30P140LVT U252 ( .A1(n3), .A2(i_data_bus[102]), .B1(n254), .B2(
        i_data_bus[134]), .ZN(n220) );
  INVD1BWP30P140LVT U253 ( .I(i_data_bus[198]), .ZN(n216) );
  INVD1BWP30P140LVT U254 ( .I(i_data_bus[166]), .ZN(n215) );
  OAI22D1BWP30P140LVT U255 ( .A1(n275), .A2(n216), .B1(n273), .B2(n215), .ZN(
        n217) );
  AOI21D1BWP30P140LVT U256 ( .A1(n277), .A2(i_data_bus[230]), .B(n217), .ZN(
        n219) );
  ND2D1BWP30P140LVT U257 ( .A1(n257), .A2(i_data_bus[6]), .ZN(n218) );
  ND4D1BWP30P140LVT U258 ( .A1(n221), .A2(n220), .A3(n219), .A4(n218), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U259 ( .A1(n270), .A2(i_data_bus[69]), .B1(n2), .B2(
        i_data_bus[37]), .ZN(n228) );
  AOI22D1BWP30P140LVT U260 ( .A1(n3), .A2(i_data_bus[101]), .B1(n254), .B2(
        i_data_bus[133]), .ZN(n227) );
  INVD1BWP30P140LVT U261 ( .I(i_data_bus[197]), .ZN(n223) );
  INVD1BWP30P140LVT U262 ( .I(i_data_bus[165]), .ZN(n222) );
  OAI22D1BWP30P140LVT U263 ( .A1(n275), .A2(n223), .B1(n273), .B2(n222), .ZN(
        n224) );
  AOI21D1BWP30P140LVT U264 ( .A1(n277), .A2(i_data_bus[229]), .B(n224), .ZN(
        n226) );
  ND2D1BWP30P140LVT U265 ( .A1(n257), .A2(i_data_bus[5]), .ZN(n225) );
  ND4D1BWP30P140LVT U266 ( .A1(n228), .A2(n227), .A3(n226), .A4(n225), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U267 ( .A1(n270), .A2(i_data_bus[64]), .B1(n2), .B2(
        i_data_bus[32]), .ZN(n234) );
  AOI22D1BWP30P140LVT U268 ( .A1(n3), .A2(i_data_bus[96]), .B1(n254), .B2(
        i_data_bus[128]), .ZN(n233) );
  INR2D1BWP30P140LVT U269 ( .A1(i_data_bus[192]), .B1(n275), .ZN(n230) );
  INR2D1BWP30P140LVT U270 ( .A1(i_data_bus[160]), .B1(n273), .ZN(n229) );
  AOI211D1BWP30P140LVT U271 ( .A1(i_data_bus[224]), .A2(n277), .B(n230), .C(
        n229), .ZN(n232) );
  ND2D1BWP30P140LVT U272 ( .A1(n257), .A2(i_data_bus[0]), .ZN(n231) );
  ND4D1BWP30P140LVT U273 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U274 ( .A1(n270), .A2(i_data_bus[68]), .B1(n2), .B2(
        i_data_bus[36]), .ZN(n241) );
  AOI22D1BWP30P140LVT U275 ( .A1(n3), .A2(i_data_bus[100]), .B1(n254), .B2(
        i_data_bus[132]), .ZN(n240) );
  INVD1BWP30P140LVT U276 ( .I(i_data_bus[196]), .ZN(n236) );
  INVD1BWP30P140LVT U277 ( .I(i_data_bus[164]), .ZN(n235) );
  OAI22D1BWP30P140LVT U278 ( .A1(n275), .A2(n236), .B1(n273), .B2(n235), .ZN(
        n237) );
  AOI21D1BWP30P140LVT U279 ( .A1(n277), .A2(i_data_bus[228]), .B(n237), .ZN(
        n239) );
  ND2D1BWP30P140LVT U280 ( .A1(n257), .A2(i_data_bus[4]), .ZN(n238) );
  ND4D1BWP30P140LVT U281 ( .A1(n241), .A2(n240), .A3(n239), .A4(n238), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U282 ( .A1(n270), .A2(i_data_bus[67]), .B1(n2), .B2(
        i_data_bus[35]), .ZN(n247) );
  AOI22D1BWP30P140LVT U283 ( .A1(n3), .A2(i_data_bus[99]), .B1(n254), .B2(
        i_data_bus[131]), .ZN(n246) );
  INVD1BWP30P140LVT U284 ( .I(i_data_bus[163]), .ZN(n242) );
  MOAI22D1BWP30P140LVT U285 ( .A1(n273), .A2(n242), .B1(n262), .B2(
        i_data_bus[195]), .ZN(n243) );
  AOI21D1BWP30P140LVT U286 ( .A1(n277), .A2(i_data_bus[227]), .B(n243), .ZN(
        n245) );
  ND2D1BWP30P140LVT U287 ( .A1(n257), .A2(i_data_bus[3]), .ZN(n244) );
  ND4D1BWP30P140LVT U288 ( .A1(n247), .A2(n246), .A3(n245), .A4(n244), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U289 ( .A1(n270), .A2(i_data_bus[66]), .B1(n2), .B2(
        i_data_bus[34]), .ZN(n253) );
  AOI22D1BWP30P140LVT U290 ( .A1(n3), .A2(i_data_bus[98]), .B1(n254), .B2(
        i_data_bus[130]), .ZN(n252) );
  INVD1BWP30P140LVT U291 ( .I(i_data_bus[162]), .ZN(n248) );
  MOAI22D1BWP30P140LVT U292 ( .A1(n273), .A2(n248), .B1(n262), .B2(
        i_data_bus[194]), .ZN(n249) );
  AOI21D1BWP30P140LVT U293 ( .A1(n277), .A2(i_data_bus[226]), .B(n249), .ZN(
        n251) );
  ND2D1BWP30P140LVT U294 ( .A1(n257), .A2(i_data_bus[2]), .ZN(n250) );
  ND4D1BWP30P140LVT U295 ( .A1(n253), .A2(n252), .A3(n251), .A4(n250), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U296 ( .A1(n270), .A2(i_data_bus[65]), .B1(n2), .B2(
        i_data_bus[33]), .ZN(n261) );
  AOI22D1BWP30P140LVT U297 ( .A1(n3), .A2(i_data_bus[97]), .B1(n254), .B2(
        i_data_bus[129]), .ZN(n260) );
  INVD1BWP30P140LVT U298 ( .I(i_data_bus[161]), .ZN(n255) );
  MOAI22D1BWP30P140LVT U299 ( .A1(n273), .A2(n255), .B1(n262), .B2(
        i_data_bus[193]), .ZN(n256) );
  AOI21D1BWP30P140LVT U300 ( .A1(n277), .A2(i_data_bus[225]), .B(n256), .ZN(
        n259) );
  ND2D1BWP30P140LVT U301 ( .A1(n257), .A2(i_data_bus[1]), .ZN(n258) );
  ND4D1BWP30P140LVT U302 ( .A1(n261), .A2(n260), .A3(n259), .A4(n258), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U303 ( .A1(n270), .A2(i_data_bus[78]), .B1(n2), .B2(
        i_data_bus[46]), .ZN(n269) );
  AOI22D1BWP30P140LVT U304 ( .A1(n3), .A2(i_data_bus[110]), .B1(n271), .B2(
        i_data_bus[142]), .ZN(n268) );
  INVD1BWP30P140LVT U305 ( .I(i_data_bus[174]), .ZN(n263) );
  MOAI22D1BWP30P140LVT U306 ( .A1(n273), .A2(n263), .B1(n262), .B2(
        i_data_bus[206]), .ZN(n264) );
  AOI21D1BWP30P140LVT U307 ( .A1(n265), .A2(i_data_bus[238]), .B(n264), .ZN(
        n267) );
  ND2D1BWP30P140LVT U308 ( .A1(n278), .A2(i_data_bus[14]), .ZN(n266) );
  ND4D1BWP30P140LVT U309 ( .A1(n269), .A2(n268), .A3(n267), .A4(n266), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U310 ( .A1(n270), .A2(i_data_bus[77]), .B1(n2), .B2(
        i_data_bus[45]), .ZN(n282) );
  AOI22D1BWP30P140LVT U311 ( .A1(n3), .A2(i_data_bus[109]), .B1(n271), .B2(
        i_data_bus[141]), .ZN(n281) );
  INVD1BWP30P140LVT U312 ( .I(i_data_bus[205]), .ZN(n274) );
  INVD1BWP30P140LVT U313 ( .I(i_data_bus[173]), .ZN(n272) );
  OAI22D1BWP30P140LVT U314 ( .A1(n275), .A2(n274), .B1(n273), .B2(n272), .ZN(
        n276) );
  AOI21D1BWP30P140LVT U315 ( .A1(n277), .A2(i_data_bus[237]), .B(n276), .ZN(
        n280) );
  ND2D1BWP30P140LVT U316 ( .A1(n278), .A2(i_data_bus[13]), .ZN(n279) );
  ND4D1BWP30P140LVT U317 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_3 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n53), .ZN(n1) );
  INVD6BWP30P140LVT U4 ( .I(n22), .ZN(n284) );
  INVD1BWP30P140LVT U5 ( .I(n31), .ZN(n65) );
  CKND2D2BWP30P140LVT U6 ( .A1(n28), .A2(n27), .ZN(n36) );
  INVD2BWP30P140LVT U7 ( .I(n157), .ZN(n2) );
  INR2D2BWP30P140LVT U8 ( .A1(n39), .B1(n36), .ZN(n32) );
  INVD1BWP30P140LVT U9 ( .I(n2), .ZN(n201) );
  INVD2BWP30P140LVT U10 ( .I(n65), .ZN(n269) );
  INVD2BWP30P140LVT U11 ( .I(n65), .ZN(n291) );
  INR2D1BWP30P140LVT U12 ( .A1(n11), .B1(n13), .ZN(n157) );
  INVD1BWP30P140LVT U13 ( .I(n15), .ZN(n158) );
  INVD1BWP30P140LVT U14 ( .I(n157), .ZN(n64) );
  AOI21D1BWP30P140LVT U15 ( .A1(n151), .A2(i_data_bus[254]), .B(n44), .ZN(n50)
         );
  BUFFD3BWP30P140LVT U16 ( .I(n67), .Z(n139) );
  ND2OPTIBD1BWP30P140LVT U17 ( .A1(n41), .A2(n40), .ZN(n67) );
  INVD1BWP30P140LVT U18 ( .I(n139), .ZN(n140) );
  INR2D1BWP30P140LVT U19 ( .A1(n9), .B1(n13), .ZN(n156) );
  INVD1BWP30P140LVT U20 ( .I(i_cmd[2]), .ZN(n3) );
  INR4D0BWP30P140LVT U21 ( .A1(i_valid[2]), .B1(i_cmd[1]), .B2(i_cmd[3]), .B3(
        n3), .ZN(n9) );
  INVD1BWP30P140LVT U22 ( .I(i_cmd[4]), .ZN(n4) );
  INVD1BWP30P140LVT U23 ( .I(i_cmd[0]), .ZN(n45) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n4), .A2(n45), .Z(n8) );
  INVD1BWP30P140LVT U25 ( .I(rst), .ZN(n5) );
  ND2D1BWP30P140LVT U26 ( .A1(n5), .A2(i_en), .ZN(n26) );
  NR2OPTPAD1BWP30P140LVT U27 ( .A1(i_cmd[5]), .A2(n26), .ZN(n18) );
  INVD1BWP30P140LVT U28 ( .I(n18), .ZN(n6) );
  OR2D2BWP30P140LVT U29 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n37) );
  NR2OPTPAD1BWP30P140LVT U30 ( .A1(n6), .A2(n37), .ZN(n7) );
  ND2OPTIBD2BWP30P140LVT U31 ( .A1(n8), .A2(n7), .ZN(n13) );
  INVD1BWP30P140LVT U32 ( .I(n156), .ZN(n53) );
  OR2D1BWP30P140LVT U33 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n16) );
  ND2D1BWP30P140LVT U34 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n10) );
  NR2D1BWP30P140LVT U35 ( .A1(n16), .A2(n10), .ZN(n11) );
  AOI22D1BWP30P140LVT U36 ( .A1(n1), .A2(i_data_bus[94]), .B1(n201), .B2(
        i_data_bus[62]), .ZN(n52) );
  OR2D4BWP30P140LVT U37 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .Z(n25) );
  ND2D1BWP30P140LVT U38 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n12) );
  NR2D1BWP30P140LVT U39 ( .A1(n25), .A2(n12), .ZN(n14) );
  INR2D1BWP30P140LVT U40 ( .A1(n14), .B1(n13), .ZN(n15) );
  INVD1BWP30P140LVT U41 ( .I(n16), .ZN(n19) );
  NR2D1BWP30P140LVT U42 ( .A1(n37), .A2(i_cmd[1]), .ZN(n17) );
  ND3D2BWP30P140LVT U43 ( .A1(n19), .A2(n18), .A3(n17), .ZN(n46) );
  ND2D1BWP30P140LVT U44 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n20) );
  OR2D1BWP30P140LVT U45 ( .A1(n20), .A2(i_cmd[0]), .Z(n21) );
  OR2D4BWP30P140LVT U46 ( .A1(n46), .A2(n21), .Z(n22) );
  AOI22D1BWP30P140LVT U47 ( .A1(n275), .A2(i_data_bus[126]), .B1(n284), .B2(
        i_data_bus[158]), .ZN(n51) );
  INVD1BWP30P140LVT U48 ( .I(i_cmd[7]), .ZN(n24) );
  INVD1BWP30P140LVT U49 ( .I(i_valid[7]), .ZN(n23) );
  NR4D0BWP30P140LVT U50 ( .A1(n24), .A2(n23), .A3(i_cmd[6]), .A4(i_cmd[5]), 
        .ZN(n30) );
  NR2D1BWP30P140LVT U51 ( .A1(i_cmd[3]), .A2(i_cmd[0]), .ZN(n39) );
  INVD2BWP30P140LVT U52 ( .I(n25), .ZN(n28) );
  NR2D1BWP30P140LVT U53 ( .A1(i_cmd[4]), .A2(n26), .ZN(n27) );
  INVD1BWP30P140LVT U54 ( .I(n32), .ZN(n29) );
  INR2D1BWP30P140LVT U55 ( .A1(n30), .B1(n29), .ZN(n31) );
  INVD1BWP30P140LVT U56 ( .I(n65), .ZN(n151) );
  ND2OPTIBD1BWP30P140LVT U57 ( .A1(i_cmd[6]), .A2(i_valid[6]), .ZN(n34) );
  NR2D1BWP30P140LVT U58 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n33) );
  IND3D2BWP30P140LVT U59 ( .A1(n34), .B1(n33), .B2(n32), .ZN(n35) );
  INVD2BWP30P140LVT U60 ( .I(n35), .ZN(n66) );
  INVD1BWP30P140LVT U61 ( .I(n66), .ZN(n239) );
  INVD1BWP30P140LVT U62 ( .I(i_data_bus[222]), .ZN(n43) );
  NR2D1BWP30P140LVT U63 ( .A1(n37), .A2(n36), .ZN(n41) );
  ND2OPTIBD1BWP30P140LVT U64 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n38) );
  INR2D1BWP30P140LVT U65 ( .A1(n39), .B1(n38), .ZN(n40) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[190]), .ZN(n42) );
  OAI22D1BWP30P140LVT U67 ( .A1(n239), .A2(n43), .B1(n139), .B2(n42), .ZN(n44)
         );
  INR3D0BWP30P140LVT U68 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n45), .ZN(n47)
         );
  INR2D1BWP30P140LVT U69 ( .A1(n47), .B1(n46), .ZN(n48) );
  INVD2BWP30P140LVT U70 ( .I(n48), .ZN(n59) );
  INVD2BWP30P140LVT U71 ( .I(n59), .ZN(n278) );
  ND2D1BWP30P140LVT U72 ( .A1(n278), .A2(i_data_bus[30]), .ZN(n49) );
  ND4D1BWP30P140LVT U73 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(N399) );
  NR4D0BWP30P140LVT U74 ( .A1(n278), .A2(n66), .A3(n140), .A4(n291), .ZN(n55)
         );
  NR2D1BWP30P140LVT U75 ( .A1(n15), .A2(n284), .ZN(n54) );
  ND4D1BWP30P140LVT U76 ( .A1(n55), .A2(n54), .A3(n53), .A4(n2), .ZN(N402) );
  AOI22D1BWP30P140LVT U77 ( .A1(n1), .A2(i_data_bus[95]), .B1(n201), .B2(
        i_data_bus[63]), .ZN(n63) );
  AOI22D1BWP30P140LVT U78 ( .A1(n285), .A2(i_data_bus[127]), .B1(n284), .B2(
        i_data_bus[159]), .ZN(n62) );
  INVD1BWP30P140LVT U79 ( .I(i_data_bus[223]), .ZN(n57) );
  INVD1BWP30P140LVT U80 ( .I(i_data_bus[191]), .ZN(n56) );
  OAI22D1BWP30P140LVT U81 ( .A1(n239), .A2(n57), .B1(n139), .B2(n56), .ZN(n58)
         );
  AOI21D1BWP30P140LVT U82 ( .A1(n291), .A2(i_data_bus[255]), .B(n58), .ZN(n61)
         );
  INVD2BWP30P140LVT U83 ( .I(n59), .ZN(n292) );
  ND2OPTIBD1BWP30P140LVT U84 ( .A1(n292), .A2(i_data_bus[31]), .ZN(n60) );
  ND4D1BWP30P140LVT U85 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(N400) );
  INVD2BWP30P140LVT U86 ( .I(n64), .ZN(n274) );
  AOI22D1BWP30P140LVT U87 ( .A1(n1), .A2(i_data_bus[72]), .B1(n274), .B2(
        i_data_bus[40]), .ZN(n75) );
  INVD2BWP30P140LVT U88 ( .I(n158), .ZN(n275) );
  AOI22D1BWP30P140LVT U89 ( .A1(n275), .A2(i_data_bus[104]), .B1(n284), .B2(
        i_data_bus[136]), .ZN(n74) );
  INVD3BWP30P140LVT U90 ( .I(n66), .ZN(n289) );
  INVD1BWP30P140LVT U91 ( .I(i_data_bus[200]), .ZN(n70) );
  INVD1BWP30P140LVT U92 ( .I(n67), .ZN(n68) );
  INVD2BWP30P140LVT U93 ( .I(n68), .ZN(n287) );
  INVD1BWP30P140LVT U94 ( .I(i_data_bus[168]), .ZN(n69) );
  OAI22D1BWP30P140LVT U95 ( .A1(n289), .A2(n70), .B1(n287), .B2(n69), .ZN(n71)
         );
  AOI21D1BWP30P140LVT U96 ( .A1(n269), .A2(i_data_bus[232]), .B(n71), .ZN(n73)
         );
  ND2D1BWP30P140LVT U97 ( .A1(n278), .A2(i_data_bus[8]), .ZN(n72) );
  ND4D1BWP30P140LVT U98 ( .A1(n75), .A2(n74), .A3(n73), .A4(n72), .ZN(N377) );
  AOI22D1BWP30P140LVT U99 ( .A1(n1), .A2(i_data_bus[73]), .B1(n274), .B2(
        i_data_bus[41]), .ZN(n82) );
  AOI22D1BWP30P140LVT U100 ( .A1(n275), .A2(i_data_bus[105]), .B1(n284), .B2(
        i_data_bus[137]), .ZN(n81) );
  INVD1BWP30P140LVT U101 ( .I(i_data_bus[201]), .ZN(n77) );
  INVD1BWP30P140LVT U102 ( .I(i_data_bus[169]), .ZN(n76) );
  OAI22D1BWP30P140LVT U103 ( .A1(n289), .A2(n77), .B1(n287), .B2(n76), .ZN(n78) );
  AOI21D1BWP30P140LVT U104 ( .A1(n291), .A2(i_data_bus[233]), .B(n78), .ZN(n80) );
  ND2D1BWP30P140LVT U105 ( .A1(n278), .A2(i_data_bus[9]), .ZN(n79) );
  ND4D1BWP30P140LVT U106 ( .A1(n82), .A2(n81), .A3(n80), .A4(n79), .ZN(N378)
         );
  AOI22D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[74]), .B1(n274), .B2(
        i_data_bus[42]), .ZN(n89) );
  AOI22D1BWP30P140LVT U108 ( .A1(n275), .A2(i_data_bus[106]), .B1(n284), .B2(
        i_data_bus[138]), .ZN(n88) );
  INVD1BWP30P140LVT U109 ( .I(i_data_bus[202]), .ZN(n84) );
  INVD1BWP30P140LVT U110 ( .I(i_data_bus[170]), .ZN(n83) );
  OAI22D1BWP30P140LVT U111 ( .A1(n289), .A2(n84), .B1(n287), .B2(n83), .ZN(n85) );
  AOI21D1BWP30P140LVT U112 ( .A1(n291), .A2(i_data_bus[234]), .B(n85), .ZN(n87) );
  ND2D1BWP30P140LVT U113 ( .A1(n278), .A2(i_data_bus[10]), .ZN(n86) );
  ND4D1BWP30P140LVT U114 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(N379)
         );
  AOI22D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[68]), .B1(n274), .B2(
        i_data_bus[36]), .ZN(n96) );
  AOI22D1BWP30P140LVT U116 ( .A1(n275), .A2(i_data_bus[100]), .B1(n284), .B2(
        i_data_bus[132]), .ZN(n95) );
  INVD1BWP30P140LVT U117 ( .I(i_data_bus[196]), .ZN(n91) );
  INVD1BWP30P140LVT U118 ( .I(i_data_bus[164]), .ZN(n90) );
  OAI22D1BWP30P140LVT U119 ( .A1(n289), .A2(n91), .B1(n287), .B2(n90), .ZN(n92) );
  AOI21D1BWP30P140LVT U120 ( .A1(n291), .A2(i_data_bus[228]), .B(n92), .ZN(n94) );
  ND2D1BWP30P140LVT U121 ( .A1(n278), .A2(i_data_bus[4]), .ZN(n93) );
  ND4D1BWP30P140LVT U122 ( .A1(n96), .A2(n95), .A3(n94), .A4(n93), .ZN(N373)
         );
  AOI22D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[76]), .B1(n274), .B2(
        i_data_bus[44]), .ZN(n103) );
  AOI22D1BWP30P140LVT U124 ( .A1(n275), .A2(i_data_bus[108]), .B1(n284), .B2(
        i_data_bus[140]), .ZN(n102) );
  INVD1BWP30P140LVT U125 ( .I(i_data_bus[204]), .ZN(n98) );
  INVD1BWP30P140LVT U126 ( .I(i_data_bus[172]), .ZN(n97) );
  OAI22D1BWP30P140LVT U127 ( .A1(n289), .A2(n98), .B1(n287), .B2(n97), .ZN(n99) );
  AOI21D1BWP30P140LVT U128 ( .A1(n291), .A2(i_data_bus[236]), .B(n99), .ZN(
        n101) );
  ND2D1BWP30P140LVT U129 ( .A1(n278), .A2(i_data_bus[12]), .ZN(n100) );
  ND4D1BWP30P140LVT U130 ( .A1(n103), .A2(n102), .A3(n101), .A4(n100), .ZN(
        N381) );
  AOI22D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[75]), .B1(n274), .B2(
        i_data_bus[43]), .ZN(n110) );
  AOI22D1BWP30P140LVT U132 ( .A1(n275), .A2(i_data_bus[107]), .B1(n284), .B2(
        i_data_bus[139]), .ZN(n109) );
  INVD1BWP30P140LVT U133 ( .I(i_data_bus[203]), .ZN(n105) );
  INVD1BWP30P140LVT U134 ( .I(i_data_bus[171]), .ZN(n104) );
  OAI22D1BWP30P140LVT U135 ( .A1(n289), .A2(n105), .B1(n287), .B2(n104), .ZN(
        n106) );
  AOI21D1BWP30P140LVT U136 ( .A1(n291), .A2(i_data_bus[235]), .B(n106), .ZN(
        n108) );
  ND2D1BWP30P140LVT U137 ( .A1(n278), .A2(i_data_bus[11]), .ZN(n107) );
  ND4D1BWP30P140LVT U138 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .ZN(
        N380) );
  AOI22D1BWP30P140LVT U139 ( .A1(n1), .A2(i_data_bus[70]), .B1(n274), .B2(
        i_data_bus[38]), .ZN(n117) );
  AOI22D1BWP30P140LVT U140 ( .A1(n275), .A2(i_data_bus[102]), .B1(n284), .B2(
        i_data_bus[134]), .ZN(n116) );
  INVD1BWP30P140LVT U141 ( .I(i_data_bus[198]), .ZN(n112) );
  INVD1BWP30P140LVT U142 ( .I(i_data_bus[166]), .ZN(n111) );
  OAI22D1BWP30P140LVT U143 ( .A1(n289), .A2(n112), .B1(n287), .B2(n111), .ZN(
        n113) );
  AOI21D1BWP30P140LVT U144 ( .A1(n291), .A2(i_data_bus[230]), .B(n113), .ZN(
        n115) );
  ND2D1BWP30P140LVT U145 ( .A1(n278), .A2(i_data_bus[6]), .ZN(n114) );
  ND4D1BWP30P140LVT U146 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U147 ( .A1(n1), .A2(i_data_bus[71]), .B1(n274), .B2(
        i_data_bus[39]), .ZN(n124) );
  AOI22D1BWP30P140LVT U148 ( .A1(n275), .A2(i_data_bus[103]), .B1(n284), .B2(
        i_data_bus[135]), .ZN(n123) );
  INVD1BWP30P140LVT U149 ( .I(i_data_bus[199]), .ZN(n119) );
  INVD1BWP30P140LVT U150 ( .I(i_data_bus[167]), .ZN(n118) );
  OAI22D1BWP30P140LVT U151 ( .A1(n289), .A2(n119), .B1(n287), .B2(n118), .ZN(
        n120) );
  AOI21D1BWP30P140LVT U152 ( .A1(n291), .A2(i_data_bus[231]), .B(n120), .ZN(
        n122) );
  ND2D1BWP30P140LVT U153 ( .A1(n278), .A2(i_data_bus[7]), .ZN(n121) );
  ND4D1BWP30P140LVT U154 ( .A1(n124), .A2(n123), .A3(n122), .A4(n121), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U155 ( .A1(n1), .A2(i_data_bus[69]), .B1(n274), .B2(
        i_data_bus[37]), .ZN(n131) );
  AOI22D1BWP30P140LVT U156 ( .A1(n275), .A2(i_data_bus[101]), .B1(n284), .B2(
        i_data_bus[133]), .ZN(n130) );
  INVD1BWP30P140LVT U157 ( .I(i_data_bus[197]), .ZN(n126) );
  INVD1BWP30P140LVT U158 ( .I(i_data_bus[165]), .ZN(n125) );
  OAI22D1BWP30P140LVT U159 ( .A1(n289), .A2(n126), .B1(n287), .B2(n125), .ZN(
        n127) );
  AOI21D1BWP30P140LVT U160 ( .A1(n291), .A2(i_data_bus[229]), .B(n127), .ZN(
        n129) );
  ND2D1BWP30P140LVT U161 ( .A1(n278), .A2(i_data_bus[5]), .ZN(n128) );
  ND4D1BWP30P140LVT U162 ( .A1(n131), .A2(n130), .A3(n129), .A4(n128), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U163 ( .A1(n1), .A2(i_data_bus[67]), .B1(n274), .B2(
        i_data_bus[35]), .ZN(n138) );
  AOI22D1BWP30P140LVT U164 ( .A1(n275), .A2(i_data_bus[99]), .B1(n284), .B2(
        i_data_bus[131]), .ZN(n137) );
  INVD1BWP30P140LVT U165 ( .I(i_data_bus[195]), .ZN(n133) );
  INVD1BWP30P140LVT U166 ( .I(i_data_bus[163]), .ZN(n132) );
  OAI22D1BWP30P140LVT U167 ( .A1(n289), .A2(n133), .B1(n287), .B2(n132), .ZN(
        n134) );
  AOI21D1BWP30P140LVT U168 ( .A1(n291), .A2(i_data_bus[227]), .B(n134), .ZN(
        n136) );
  ND2D1BWP30P140LVT U169 ( .A1(n278), .A2(i_data_bus[3]), .ZN(n135) );
  ND4D1BWP30P140LVT U170 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U171 ( .A1(n1), .A2(i_data_bus[93]), .B1(n201), .B2(
        i_data_bus[61]), .ZN(n147) );
  AOI22D1BWP30P140LVT U172 ( .A1(n285), .A2(i_data_bus[125]), .B1(n284), .B2(
        i_data_bus[157]), .ZN(n146) );
  INVD1BWP30P140LVT U173 ( .I(i_data_bus[221]), .ZN(n142) );
  INVD1BWP30P140LVT U174 ( .I(i_data_bus[189]), .ZN(n141) );
  OAI22D1BWP30P140LVT U175 ( .A1(n239), .A2(n142), .B1(n139), .B2(n141), .ZN(
        n143) );
  AOI21D1BWP30P140LVT U176 ( .A1(n151), .A2(i_data_bus[253]), .B(n143), .ZN(
        n145) );
  ND2OPTIBD1BWP30P140LVT U177 ( .A1(n292), .A2(i_data_bus[29]), .ZN(n144) );
  ND4D1BWP30P140LVT U178 ( .A1(n147), .A2(n146), .A3(n145), .A4(n144), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U179 ( .A1(n1), .A2(i_data_bus[92]), .B1(n201), .B2(
        i_data_bus[60]), .ZN(n155) );
  AOI22D1BWP30P140LVT U180 ( .A1(n275), .A2(i_data_bus[124]), .B1(n284), .B2(
        i_data_bus[156]), .ZN(n154) );
  INVD1BWP30P140LVT U181 ( .I(i_data_bus[220]), .ZN(n149) );
  INVD1BWP30P140LVT U182 ( .I(i_data_bus[188]), .ZN(n148) );
  OAI22D1BWP30P140LVT U183 ( .A1(n239), .A2(n149), .B1(n139), .B2(n148), .ZN(
        n150) );
  AOI21D1BWP30P140LVT U184 ( .A1(n151), .A2(i_data_bus[252]), .B(n150), .ZN(
        n153) );
  ND2OPTIBD1BWP30P140LVT U185 ( .A1(n292), .A2(i_data_bus[28]), .ZN(n152) );
  ND4D1BWP30P140LVT U186 ( .A1(n155), .A2(n154), .A3(n153), .A4(n152), .ZN(
        N397) );
  INVD2BWP30P140LVT U187 ( .I(n2), .ZN(n283) );
  AOI22D1BWP30P140LVT U188 ( .A1(n1), .A2(i_data_bus[88]), .B1(n283), .B2(
        i_data_bus[56]), .ZN(n165) );
  INVD2BWP30P140LVT U189 ( .I(n158), .ZN(n285) );
  AOI22D1BWP30P140LVT U190 ( .A1(n285), .A2(i_data_bus[120]), .B1(n284), .B2(
        i_data_bus[152]), .ZN(n164) );
  INVD1BWP30P140LVT U191 ( .I(i_data_bus[216]), .ZN(n160) );
  INVD1BWP30P140LVT U192 ( .I(i_data_bus[184]), .ZN(n159) );
  OAI22D1BWP30P140LVT U193 ( .A1(n289), .A2(n160), .B1(n139), .B2(n159), .ZN(
        n161) );
  AOI21D1BWP30P140LVT U194 ( .A1(n269), .A2(i_data_bus[248]), .B(n161), .ZN(
        n163) );
  ND2OPTIBD1BWP30P140LVT U195 ( .A1(n292), .A2(i_data_bus[24]), .ZN(n162) );
  ND4D1BWP30P140LVT U196 ( .A1(n165), .A2(n164), .A3(n163), .A4(n162), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U197 ( .A1(n1), .A2(i_data_bus[80]), .B1(n283), .B2(
        i_data_bus[48]), .ZN(n172) );
  AOI22D1BWP30P140LVT U198 ( .A1(n285), .A2(i_data_bus[112]), .B1(n284), .B2(
        i_data_bus[144]), .ZN(n171) );
  INVD1BWP30P140LVT U199 ( .I(i_data_bus[208]), .ZN(n167) );
  INVD1BWP30P140LVT U200 ( .I(i_data_bus[176]), .ZN(n166) );
  OAI22D1BWP30P140LVT U201 ( .A1(n289), .A2(n167), .B1(n139), .B2(n166), .ZN(
        n168) );
  AOI21D1BWP30P140LVT U202 ( .A1(n269), .A2(i_data_bus[240]), .B(n168), .ZN(
        n170) );
  ND2OPTIBD1BWP30P140LVT U203 ( .A1(n292), .A2(i_data_bus[16]), .ZN(n169) );
  ND4D1BWP30P140LVT U204 ( .A1(n172), .A2(n171), .A3(n170), .A4(n169), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U205 ( .A1(n1), .A2(i_data_bus[87]), .B1(n283), .B2(
        i_data_bus[55]), .ZN(n179) );
  AOI22D1BWP30P140LVT U206 ( .A1(n285), .A2(i_data_bus[119]), .B1(n284), .B2(
        i_data_bus[151]), .ZN(n178) );
  INVD1BWP30P140LVT U207 ( .I(i_data_bus[215]), .ZN(n174) );
  INVD1BWP30P140LVT U208 ( .I(i_data_bus[183]), .ZN(n173) );
  OAI22D1BWP30P140LVT U209 ( .A1(n289), .A2(n174), .B1(n139), .B2(n173), .ZN(
        n175) );
  AOI21D1BWP30P140LVT U210 ( .A1(n269), .A2(i_data_bus[247]), .B(n175), .ZN(
        n177) );
  ND2OPTIBD1BWP30P140LVT U211 ( .A1(n292), .A2(i_data_bus[23]), .ZN(n176) );
  ND4D1BWP30P140LVT U212 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U213 ( .A1(n1), .A2(i_data_bus[90]), .B1(n201), .B2(
        i_data_bus[58]), .ZN(n186) );
  AOI22D1BWP30P140LVT U214 ( .A1(n285), .A2(i_data_bus[122]), .B1(n284), .B2(
        i_data_bus[154]), .ZN(n185) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[218]), .ZN(n181) );
  INVD1BWP30P140LVT U216 ( .I(i_data_bus[186]), .ZN(n180) );
  OAI22D1BWP30P140LVT U217 ( .A1(n239), .A2(n181), .B1(n139), .B2(n180), .ZN(
        n182) );
  AOI21D1BWP30P140LVT U218 ( .A1(n269), .A2(i_data_bus[250]), .B(n182), .ZN(
        n184) );
  ND2OPTIBD1BWP30P140LVT U219 ( .A1(n292), .A2(i_data_bus[26]), .ZN(n183) );
  ND4D1BWP30P140LVT U220 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U221 ( .A1(n1), .A2(i_data_bus[85]), .B1(n283), .B2(
        i_data_bus[53]), .ZN(n193) );
  AOI22D1BWP30P140LVT U222 ( .A1(n285), .A2(i_data_bus[117]), .B1(n284), .B2(
        i_data_bus[149]), .ZN(n192) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[213]), .ZN(n188) );
  INVD1BWP30P140LVT U224 ( .I(i_data_bus[181]), .ZN(n187) );
  OAI22D1BWP30P140LVT U225 ( .A1(n289), .A2(n188), .B1(n139), .B2(n187), .ZN(
        n189) );
  AOI21D1BWP30P140LVT U226 ( .A1(n269), .A2(i_data_bus[245]), .B(n189), .ZN(
        n191) );
  ND2OPTIBD1BWP30P140LVT U227 ( .A1(n292), .A2(i_data_bus[21]), .ZN(n190) );
  ND4D1BWP30P140LVT U228 ( .A1(n193), .A2(n192), .A3(n191), .A4(n190), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U229 ( .A1(n1), .A2(i_data_bus[86]), .B1(n283), .B2(
        i_data_bus[54]), .ZN(n200) );
  AOI22D1BWP30P140LVT U230 ( .A1(n285), .A2(i_data_bus[118]), .B1(n284), .B2(
        i_data_bus[150]), .ZN(n199) );
  INVD1BWP30P140LVT U231 ( .I(i_data_bus[214]), .ZN(n195) );
  INVD1BWP30P140LVT U232 ( .I(i_data_bus[182]), .ZN(n194) );
  OAI22D1BWP30P140LVT U233 ( .A1(n289), .A2(n195), .B1(n139), .B2(n194), .ZN(
        n196) );
  AOI21D1BWP30P140LVT U234 ( .A1(n269), .A2(i_data_bus[246]), .B(n196), .ZN(
        n198) );
  ND2OPTIBD1BWP30P140LVT U235 ( .A1(n292), .A2(i_data_bus[22]), .ZN(n197) );
  ND4D1BWP30P140LVT U236 ( .A1(n200), .A2(n199), .A3(n198), .A4(n197), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U237 ( .A1(n1), .A2(i_data_bus[91]), .B1(n201), .B2(
        i_data_bus[59]), .ZN(n208) );
  AOI22D1BWP30P140LVT U238 ( .A1(n275), .A2(i_data_bus[123]), .B1(n284), .B2(
        i_data_bus[155]), .ZN(n207) );
  INVD1BWP30P140LVT U239 ( .I(i_data_bus[219]), .ZN(n203) );
  INVD1BWP30P140LVT U240 ( .I(i_data_bus[187]), .ZN(n202) );
  OAI22D1BWP30P140LVT U241 ( .A1(n239), .A2(n203), .B1(n139), .B2(n202), .ZN(
        n204) );
  AOI21D1BWP30P140LVT U242 ( .A1(n269), .A2(i_data_bus[251]), .B(n204), .ZN(
        n206) );
  ND2OPTIBD1BWP30P140LVT U243 ( .A1(n292), .A2(i_data_bus[27]), .ZN(n205) );
  ND4D1BWP30P140LVT U244 ( .A1(n208), .A2(n207), .A3(n206), .A4(n205), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U245 ( .A1(n1), .A2(i_data_bus[83]), .B1(n283), .B2(
        i_data_bus[51]), .ZN(n215) );
  AOI22D1BWP30P140LVT U246 ( .A1(n285), .A2(i_data_bus[115]), .B1(n284), .B2(
        i_data_bus[147]), .ZN(n214) );
  INVD1BWP30P140LVT U247 ( .I(i_data_bus[211]), .ZN(n210) );
  INVD1BWP30P140LVT U248 ( .I(i_data_bus[179]), .ZN(n209) );
  OAI22D1BWP30P140LVT U249 ( .A1(n289), .A2(n210), .B1(n139), .B2(n209), .ZN(
        n211) );
  AOI21D1BWP30P140LVT U250 ( .A1(n269), .A2(i_data_bus[243]), .B(n211), .ZN(
        n213) );
  ND2OPTIBD1BWP30P140LVT U251 ( .A1(n292), .A2(i_data_bus[19]), .ZN(n212) );
  ND4D1BWP30P140LVT U252 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[84]), .B1(n283), .B2(
        i_data_bus[52]), .ZN(n222) );
  AOI22D1BWP30P140LVT U254 ( .A1(n285), .A2(i_data_bus[116]), .B1(n284), .B2(
        i_data_bus[148]), .ZN(n221) );
  INVD1BWP30P140LVT U255 ( .I(i_data_bus[212]), .ZN(n217) );
  INVD1BWP30P140LVT U256 ( .I(i_data_bus[180]), .ZN(n216) );
  OAI22D1BWP30P140LVT U257 ( .A1(n289), .A2(n217), .B1(n139), .B2(n216), .ZN(
        n218) );
  AOI21D1BWP30P140LVT U258 ( .A1(n269), .A2(i_data_bus[244]), .B(n218), .ZN(
        n220) );
  ND2OPTIBD1BWP30P140LVT U259 ( .A1(n292), .A2(i_data_bus[20]), .ZN(n219) );
  ND4D1BWP30P140LVT U260 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[81]), .B1(n283), .B2(
        i_data_bus[49]), .ZN(n229) );
  AOI22D1BWP30P140LVT U262 ( .A1(n285), .A2(i_data_bus[113]), .B1(n284), .B2(
        i_data_bus[145]), .ZN(n228) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[209]), .ZN(n224) );
  INVD1BWP30P140LVT U264 ( .I(i_data_bus[177]), .ZN(n223) );
  OAI22D1BWP30P140LVT U265 ( .A1(n289), .A2(n224), .B1(n139), .B2(n223), .ZN(
        n225) );
  AOI21D1BWP30P140LVT U266 ( .A1(n269), .A2(i_data_bus[241]), .B(n225), .ZN(
        n227) );
  ND2OPTIBD1BWP30P140LVT U267 ( .A1(n292), .A2(i_data_bus[17]), .ZN(n226) );
  ND4D1BWP30P140LVT U268 ( .A1(n229), .A2(n228), .A3(n227), .A4(n226), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U269 ( .A1(n1), .A2(i_data_bus[82]), .B1(n283), .B2(
        i_data_bus[50]), .ZN(n236) );
  AOI22D1BWP30P140LVT U270 ( .A1(n285), .A2(i_data_bus[114]), .B1(n284), .B2(
        i_data_bus[146]), .ZN(n235) );
  INVD1BWP30P140LVT U271 ( .I(i_data_bus[210]), .ZN(n231) );
  INVD1BWP30P140LVT U272 ( .I(i_data_bus[178]), .ZN(n230) );
  OAI22D1BWP30P140LVT U273 ( .A1(n289), .A2(n231), .B1(n139), .B2(n230), .ZN(
        n232) );
  AOI21D1BWP30P140LVT U274 ( .A1(n269), .A2(i_data_bus[242]), .B(n232), .ZN(
        n234) );
  ND2OPTIBD1BWP30P140LVT U275 ( .A1(n292), .A2(i_data_bus[18]), .ZN(n233) );
  ND4D1BWP30P140LVT U276 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U277 ( .A1(n1), .A2(i_data_bus[89]), .B1(n283), .B2(
        i_data_bus[57]), .ZN(n244) );
  AOI22D1BWP30P140LVT U278 ( .A1(n285), .A2(i_data_bus[121]), .B1(n284), .B2(
        i_data_bus[153]), .ZN(n243) );
  INVD1BWP30P140LVT U279 ( .I(i_data_bus[217]), .ZN(n238) );
  INVD1BWP30P140LVT U280 ( .I(i_data_bus[185]), .ZN(n237) );
  OAI22D1BWP30P140LVT U281 ( .A1(n239), .A2(n238), .B1(n139), .B2(n237), .ZN(
        n240) );
  AOI21D1BWP30P140LVT U282 ( .A1(n269), .A2(i_data_bus[249]), .B(n240), .ZN(
        n242) );
  ND2OPTIBD1BWP30P140LVT U283 ( .A1(n292), .A2(i_data_bus[25]), .ZN(n241) );
  ND4D1BWP30P140LVT U284 ( .A1(n244), .A2(n243), .A3(n242), .A4(n241), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U285 ( .A1(n1), .A2(i_data_bus[66]), .B1(n274), .B2(
        i_data_bus[34]), .ZN(n251) );
  AOI22D1BWP30P140LVT U286 ( .A1(n275), .A2(i_data_bus[98]), .B1(n284), .B2(
        i_data_bus[130]), .ZN(n250) );
  INVD1BWP30P140LVT U287 ( .I(i_data_bus[194]), .ZN(n246) );
  INVD1BWP30P140LVT U288 ( .I(i_data_bus[162]), .ZN(n245) );
  OAI22D1BWP30P140LVT U289 ( .A1(n289), .A2(n246), .B1(n287), .B2(n245), .ZN(
        n247) );
  AOI21D1BWP30P140LVT U290 ( .A1(n291), .A2(i_data_bus[226]), .B(n247), .ZN(
        n249) );
  ND2D1BWP30P140LVT U291 ( .A1(n278), .A2(i_data_bus[2]), .ZN(n248) );
  ND4D1BWP30P140LVT U292 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U293 ( .A1(n1), .A2(i_data_bus[65]), .B1(n274), .B2(
        i_data_bus[33]), .ZN(n258) );
  AOI22D1BWP30P140LVT U294 ( .A1(n275), .A2(i_data_bus[97]), .B1(n284), .B2(
        i_data_bus[129]), .ZN(n257) );
  INVD1BWP30P140LVT U295 ( .I(i_data_bus[193]), .ZN(n253) );
  INVD1BWP30P140LVT U296 ( .I(i_data_bus[161]), .ZN(n252) );
  OAI22D1BWP30P140LVT U297 ( .A1(n289), .A2(n253), .B1(n287), .B2(n252), .ZN(
        n254) );
  AOI21D1BWP30P140LVT U298 ( .A1(n291), .A2(i_data_bus[225]), .B(n254), .ZN(
        n256) );
  ND2D1BWP30P140LVT U299 ( .A1(n278), .A2(i_data_bus[1]), .ZN(n255) );
  ND4D1BWP30P140LVT U300 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U301 ( .A1(n1), .A2(i_data_bus[79]), .B1(n283), .B2(
        i_data_bus[47]), .ZN(n265) );
  AOI22D1BWP30P140LVT U302 ( .A1(n285), .A2(i_data_bus[111]), .B1(n284), .B2(
        i_data_bus[143]), .ZN(n264) );
  INVD1BWP30P140LVT U303 ( .I(i_data_bus[207]), .ZN(n260) );
  INVD1BWP30P140LVT U304 ( .I(i_data_bus[175]), .ZN(n259) );
  OAI22D1BWP30P140LVT U305 ( .A1(n289), .A2(n260), .B1(n139), .B2(n259), .ZN(
        n261) );
  AOI21D1BWP30P140LVT U306 ( .A1(n269), .A2(i_data_bus[239]), .B(n261), .ZN(
        n263) );
  ND2OPTIBD1BWP30P140LVT U307 ( .A1(n292), .A2(i_data_bus[15]), .ZN(n262) );
  ND4D1BWP30P140LVT U308 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U309 ( .A1(n1), .A2(i_data_bus[78]), .B1(n283), .B2(
        i_data_bus[46]), .ZN(n273) );
  AOI22D1BWP30P140LVT U310 ( .A1(n285), .A2(i_data_bus[110]), .B1(n284), .B2(
        i_data_bus[142]), .ZN(n272) );
  INVD1BWP30P140LVT U311 ( .I(i_data_bus[206]), .ZN(n267) );
  INVD1BWP30P140LVT U312 ( .I(i_data_bus[174]), .ZN(n266) );
  OAI22D1BWP30P140LVT U313 ( .A1(n289), .A2(n267), .B1(n287), .B2(n266), .ZN(
        n268) );
  AOI21D1BWP30P140LVT U314 ( .A1(n269), .A2(i_data_bus[238]), .B(n268), .ZN(
        n271) );
  ND2OPTIBD1BWP30P140LVT U315 ( .A1(n292), .A2(i_data_bus[14]), .ZN(n270) );
  ND4D1BWP30P140LVT U316 ( .A1(n273), .A2(n272), .A3(n271), .A4(n270), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U317 ( .A1(n1), .A2(i_data_bus[64]), .B1(n274), .B2(
        i_data_bus[32]), .ZN(n282) );
  AOI22D1BWP30P140LVT U318 ( .A1(n275), .A2(i_data_bus[96]), .B1(n284), .B2(
        i_data_bus[128]), .ZN(n281) );
  INR2D1BWP30P140LVT U319 ( .A1(i_data_bus[192]), .B1(n289), .ZN(n277) );
  INR2D1BWP30P140LVT U320 ( .A1(i_data_bus[160]), .B1(n287), .ZN(n276) );
  AOI211D1BWP30P140LVT U321 ( .A1(i_data_bus[224]), .A2(n291), .B(n277), .C(
        n276), .ZN(n280) );
  ND2D1BWP30P140LVT U322 ( .A1(n278), .A2(i_data_bus[0]), .ZN(n279) );
  ND4D1BWP30P140LVT U323 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U324 ( .A1(n1), .A2(i_data_bus[77]), .B1(n283), .B2(
        i_data_bus[45]), .ZN(n296) );
  AOI22D1BWP30P140LVT U325 ( .A1(n285), .A2(i_data_bus[109]), .B1(n284), .B2(
        i_data_bus[141]), .ZN(n295) );
  INVD1BWP30P140LVT U326 ( .I(i_data_bus[205]), .ZN(n288) );
  INVD1BWP30P140LVT U327 ( .I(i_data_bus[173]), .ZN(n286) );
  OAI22D1BWP30P140LVT U328 ( .A1(n289), .A2(n288), .B1(n287), .B2(n286), .ZN(
        n290) );
  AOI21D1BWP30P140LVT U329 ( .A1(n291), .A2(i_data_bus[237]), .B(n290), .ZN(
        n294) );
  ND2OPTIBD1BWP30P140LVT U330 ( .A1(n292), .A2(i_data_bus[13]), .ZN(n293) );
  ND4D1BWP30P140LVT U331 ( .A1(n296), .A2(n295), .A3(n294), .A4(n293), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_4 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n56), .ZN(n284) );
  INVD2BWP30P140LVT U4 ( .I(n275), .ZN(n2) );
  INVD4BWP30P140LVT U5 ( .I(n275), .ZN(n289) );
  INVD3BWP30P140LVT U6 ( .I(n121), .ZN(n1) );
  INVD3BWP30P140LVT U7 ( .I(n161), .ZN(n3) );
  INVD2BWP30P140LVT U8 ( .I(n265), .ZN(n4) );
  INVD2BWP30P140LVT U9 ( .I(n157), .ZN(n147) );
  OAI22D1BWP30P140LVT U10 ( .A1(n2), .A2(n159), .B1(n226), .B2(n158), .ZN(n160) );
  ND2D1BWP30P140LVT U11 ( .A1(n16), .A2(n45), .ZN(n50) );
  INVD1BWP30P140LVT U12 ( .I(n35), .ZN(n51) );
  NR2D1BWP30P140LVT U13 ( .A1(n48), .A2(n46), .ZN(n35) );
  ND2OPTIBD1BWP30P140LVT U14 ( .A1(n5), .A2(n9), .ZN(n23) );
  INVD2BWP30P140LVT U15 ( .I(n56), .ZN(n266) );
  ND2D1BWP30P140LVT U16 ( .A1(n275), .A2(i_data_bus[193]), .ZN(n268) );
  ND2D1BWP30P140LVT U17 ( .A1(n275), .A2(i_data_bus[197]), .ZN(n57) );
  NR3OPTPAD2BWP30P140LVT U18 ( .A1(n48), .A2(n47), .A3(n46), .ZN(n265) );
  NR2D1BWP30P140LVT U19 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .ZN(n44) );
  AOI21D1BWP30P140LVT U20 ( .A1(n132), .A2(i_data_bus[249]), .B(n160), .ZN(
        n163) );
  OR3D1BWP30P140LVT U21 ( .A1(n40), .A2(n50), .A3(n18), .Z(n161) );
  ND2OPTIBD1BWP30P140LVT U22 ( .A1(n26), .A2(n25), .ZN(n137) );
  INVD2BWP30P140LVT U23 ( .I(n137), .ZN(n132) );
  INVD3BWP30P140LVT U24 ( .I(n1), .ZN(n287) );
  INVD3BWP30P140LVT U25 ( .I(n1), .ZN(n226) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n16), .A2(n8), .Z(n5) );
  INVD1BWP30P140LVT U27 ( .I(i_cmd[3]), .ZN(n16) );
  INVD1BWP30P140LVT U28 ( .I(rst), .ZN(n6) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n6), .A2(i_en), .Z(n31) );
  INVD1BWP30P140LVT U30 ( .I(n31), .ZN(n7) );
  NR2D1BWP30P140LVT U31 ( .A1(i_cmd[0]), .A2(n7), .ZN(n8) );
  OR2D4BWP30P140LVT U32 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n30) );
  NR2D1BWP30P140LVT U33 ( .A1(i_cmd[4]), .A2(n30), .ZN(n9) );
  INVD2BWP30P140LVT U34 ( .I(i_cmd[6]), .ZN(n10) );
  INVD2BWP30P140LVT U35 ( .I(i_cmd[7]), .ZN(n24) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(n10), .A2(n24), .ZN(n14) );
  INVD1BWP30P140LVT U37 ( .I(n14), .ZN(n11) );
  ND3D1BWP30P140LVT U38 ( .A1(n11), .A2(i_valid[5]), .A3(i_cmd[5]), .ZN(n12)
         );
  NR2OPTPAD1BWP30P140LVT U39 ( .A1(n23), .A2(n12), .ZN(n13) );
  INVD2BWP30P140LVT U40 ( .I(n13), .ZN(n121) );
  NR2OPTPAD1BWP30P140LVT U41 ( .A1(n14), .A2(i_cmd[5]), .ZN(n32) );
  INR2D1BWP30P140LVT U42 ( .A1(n31), .B1(i_cmd[1]), .ZN(n15) );
  ND2OPTIBD1BWP30P140LVT U43 ( .A1(n32), .A2(n15), .ZN(n40) );
  INVD1BWP30P140LVT U44 ( .I(i_cmd[2]), .ZN(n45) );
  INVD1BWP30P140LVT U45 ( .I(i_cmd[0]), .ZN(n33) );
  INR3D0BWP30P140LVT U46 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n33), .ZN(n17)
         );
  INVD1BWP30P140LVT U47 ( .I(n17), .ZN(n18) );
  ND2D1BWP30P140LVT U48 ( .A1(n226), .A2(n161), .ZN(n28) );
  NR2D1BWP30P140LVT U49 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n20) );
  CKAN2D1BWP30P140LVT U50 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n19) );
  ND2OPTIBD1BWP30P140LVT U51 ( .A1(n20), .A2(n19), .ZN(n21) );
  OR2D2BWP30P140LVT U52 ( .A1(n23), .A2(n21), .Z(n22) );
  INVD4BWP30P140LVT U53 ( .I(n22), .ZN(n275) );
  INVD1BWP30P140LVT U54 ( .I(n23), .ZN(n26) );
  INR4D0BWP30P140LVT U55 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n24), .ZN(n25) );
  ND2D1BWP30P140LVT U56 ( .A1(n2), .A2(n137), .ZN(n27) );
  NR2D1BWP30P140LVT U57 ( .A1(n28), .A2(n27), .ZN(n54) );
  ND2D1BWP30P140LVT U58 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n29) );
  NR2D1BWP30P140LVT U59 ( .A1(n30), .A2(n29), .ZN(n36) );
  ND2OPTIBD2BWP30P140LVT U60 ( .A1(n32), .A2(n31), .ZN(n48) );
  INVD1BWP30P140LVT U61 ( .I(i_cmd[4]), .ZN(n34) );
  ND2OPTIBD1BWP30P140LVT U62 ( .A1(n34), .A2(n33), .ZN(n46) );
  INR2D1BWP30P140LVT U63 ( .A1(n36), .B1(n51), .ZN(n37) );
  INVD2BWP30P140LVT U64 ( .I(n37), .ZN(n157) );
  ND2OPTIBD1BWP30P140LVT U65 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n38) );
  NR2D1BWP30P140LVT U66 ( .A1(n38), .A2(i_cmd[0]), .ZN(n42) );
  INVD1BWP30P140LVT U67 ( .I(n50), .ZN(n39) );
  IND2D2BWP30P140LVT U68 ( .A1(n40), .B1(n39), .ZN(n41) );
  INR2D2BWP30P140LVT U69 ( .A1(n42), .B1(n41), .ZN(n43) );
  INVD2BWP30P140LVT U70 ( .I(n43), .ZN(n56) );
  NR2D1BWP30P140LVT U71 ( .A1(n147), .A2(n284), .ZN(n53) );
  IND3D1BWP30P140LVT U72 ( .A1(n45), .B1(i_valid[2]), .B2(n44), .ZN(n47) );
  ND2D1BWP30P140LVT U73 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n49) );
  NR2D1BWP30P140LVT U74 ( .A1(n50), .A2(n49), .ZN(n52) );
  INR2D2BWP30P140LVT U75 ( .A1(n52), .B1(n51), .ZN(n155) );
  INVD1BWP30P140LVT U76 ( .I(n155), .ZN(n64) );
  ND4D1BWP30P140LVT U77 ( .A1(n54), .A2(n53), .A3(n4), .A4(n64), .ZN(N402) );
  INVD2BWP30P140LVT U78 ( .I(n155), .ZN(n55) );
  INVD2BWP30P140LVT U79 ( .I(n55), .ZN(n264) );
  AOI22D1BWP30P140LVT U80 ( .A1(n265), .A2(i_data_bus[69]), .B1(n264), .B2(
        i_data_bus[37]), .ZN(n63) );
  INVD2BWP30P140LVT U81 ( .I(n157), .ZN(n267) );
  AOI22D1BWP30P140LVT U82 ( .A1(n267), .A2(i_data_bus[101]), .B1(n266), .B2(
        i_data_bus[133]), .ZN(n62) );
  INVD1BWP30P140LVT U83 ( .I(i_data_bus[165]), .ZN(n58) );
  OAI21D1BWP30P140LVT U84 ( .A1(n287), .A2(n58), .B(n57), .ZN(n59) );
  AOI21D1BWP30P140LVT U85 ( .A1(n132), .A2(i_data_bus[229]), .B(n59), .ZN(n61)
         );
  ND2D1BWP30P140LVT U86 ( .A1(n3), .A2(i_data_bus[5]), .ZN(n60) );
  ND4D1BWP30P140LVT U87 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(N374) );
  INVD1BWP30P140LVT U88 ( .I(n4), .ZN(n146) );
  INVD2BWP30P140LVT U89 ( .I(n64), .ZN(n145) );
  AOI22D1BWP30P140LVT U90 ( .A1(n146), .A2(i_data_bus[95]), .B1(n145), .B2(
        i_data_bus[63]), .ZN(n71) );
  AOI22D1BWP30P140LVT U91 ( .A1(n147), .A2(i_data_bus[127]), .B1(n284), .B2(
        i_data_bus[159]), .ZN(n70) );
  INVD1BWP30P140LVT U92 ( .I(i_data_bus[223]), .ZN(n66) );
  INVD1BWP30P140LVT U93 ( .I(i_data_bus[191]), .ZN(n65) );
  OAI22D1BWP30P140LVT U94 ( .A1(n2), .A2(n66), .B1(n287), .B2(n65), .ZN(n67)
         );
  AOI21D1BWP30P140LVT U95 ( .A1(n132), .A2(i_data_bus[255]), .B(n67), .ZN(n69)
         );
  ND2D1BWP30P140LVT U96 ( .A1(n3), .A2(i_data_bus[31]), .ZN(n68) );
  ND4D1BWP30P140LVT U97 ( .A1(n71), .A2(n70), .A3(n69), .A4(n68), .ZN(N400) );
  AOI22D1BWP30P140LVT U98 ( .A1(n146), .A2(i_data_bus[94]), .B1(n145), .B2(
        i_data_bus[62]), .ZN(n78) );
  AOI22D1BWP30P140LVT U99 ( .A1(n147), .A2(i_data_bus[126]), .B1(n284), .B2(
        i_data_bus[158]), .ZN(n77) );
  INVD1BWP30P140LVT U100 ( .I(i_data_bus[222]), .ZN(n73) );
  INVD1BWP30P140LVT U101 ( .I(i_data_bus[190]), .ZN(n72) );
  OAI22D1BWP30P140LVT U102 ( .A1(n2), .A2(n73), .B1(n226), .B2(n72), .ZN(n74)
         );
  AOI21D1BWP30P140LVT U103 ( .A1(n132), .A2(i_data_bus[254]), .B(n74), .ZN(n76) );
  ND2D1BWP30P140LVT U104 ( .A1(n3), .A2(i_data_bus[30]), .ZN(n75) );
  ND4D1BWP30P140LVT U105 ( .A1(n78), .A2(n77), .A3(n76), .A4(n75), .ZN(N399)
         );
  AOI22D1BWP30P140LVT U106 ( .A1(n265), .A2(i_data_bus[76]), .B1(n264), .B2(
        i_data_bus[44]), .ZN(n85) );
  AOI22D1BWP30P140LVT U107 ( .A1(n267), .A2(i_data_bus[108]), .B1(n266), .B2(
        i_data_bus[140]), .ZN(n84) );
  INVD1BWP30P140LVT U108 ( .I(i_data_bus[204]), .ZN(n80) );
  INVD1BWP30P140LVT U109 ( .I(i_data_bus[172]), .ZN(n79) );
  OAI22D1BWP30P140LVT U110 ( .A1(n289), .A2(n80), .B1(n287), .B2(n79), .ZN(n81) );
  AOI21D1BWP30P140LVT U111 ( .A1(n132), .A2(i_data_bus[236]), .B(n81), .ZN(n83) );
  ND2D1BWP30P140LVT U112 ( .A1(n3), .A2(i_data_bus[12]), .ZN(n82) );
  ND4D1BWP30P140LVT U113 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(N381)
         );
  AOI22D1BWP30P140LVT U114 ( .A1(n265), .A2(i_data_bus[75]), .B1(n264), .B2(
        i_data_bus[43]), .ZN(n92) );
  AOI22D1BWP30P140LVT U115 ( .A1(n267), .A2(i_data_bus[107]), .B1(n266), .B2(
        i_data_bus[139]), .ZN(n91) );
  INVD1BWP30P140LVT U116 ( .I(i_data_bus[203]), .ZN(n87) );
  INVD1BWP30P140LVT U117 ( .I(i_data_bus[171]), .ZN(n86) );
  OAI22D1BWP30P140LVT U118 ( .A1(n289), .A2(n87), .B1(n287), .B2(n86), .ZN(n88) );
  AOI21D1BWP30P140LVT U119 ( .A1(n132), .A2(i_data_bus[235]), .B(n88), .ZN(n90) );
  ND2D1BWP30P140LVT U120 ( .A1(n3), .A2(i_data_bus[11]), .ZN(n89) );
  ND4D1BWP30P140LVT U121 ( .A1(n92), .A2(n91), .A3(n90), .A4(n89), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U122 ( .A1(n265), .A2(i_data_bus[74]), .B1(n264), .B2(
        i_data_bus[42]), .ZN(n99) );
  AOI22D1BWP30P140LVT U123 ( .A1(n267), .A2(i_data_bus[106]), .B1(n266), .B2(
        i_data_bus[138]), .ZN(n98) );
  INVD1BWP30P140LVT U124 ( .I(i_data_bus[202]), .ZN(n94) );
  INVD1BWP30P140LVT U125 ( .I(i_data_bus[170]), .ZN(n93) );
  OAI22D1BWP30P140LVT U126 ( .A1(n289), .A2(n94), .B1(n287), .B2(n93), .ZN(n95) );
  AOI21D1BWP30P140LVT U127 ( .A1(n132), .A2(i_data_bus[234]), .B(n95), .ZN(n97) );
  ND2D1BWP30P140LVT U128 ( .A1(n3), .A2(i_data_bus[10]), .ZN(n96) );
  ND4D1BWP30P140LVT U129 ( .A1(n99), .A2(n98), .A3(n97), .A4(n96), .ZN(N379)
         );
  AOI22D1BWP30P140LVT U130 ( .A1(n265), .A2(i_data_bus[73]), .B1(n264), .B2(
        i_data_bus[41]), .ZN(n106) );
  AOI22D1BWP30P140LVT U131 ( .A1(n267), .A2(i_data_bus[105]), .B1(n266), .B2(
        i_data_bus[137]), .ZN(n105) );
  INVD1BWP30P140LVT U132 ( .I(i_data_bus[201]), .ZN(n101) );
  INVD1BWP30P140LVT U133 ( .I(i_data_bus[169]), .ZN(n100) );
  OAI22D1BWP30P140LVT U134 ( .A1(n289), .A2(n101), .B1(n287), .B2(n100), .ZN(
        n102) );
  AOI21D1BWP30P140LVT U135 ( .A1(n132), .A2(i_data_bus[233]), .B(n102), .ZN(
        n104) );
  ND2D1BWP30P140LVT U136 ( .A1(n3), .A2(i_data_bus[9]), .ZN(n103) );
  ND4D1BWP30P140LVT U137 ( .A1(n106), .A2(n105), .A3(n104), .A4(n103), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U138 ( .A1(n265), .A2(i_data_bus[71]), .B1(n264), .B2(
        i_data_bus[39]), .ZN(n113) );
  AOI22D1BWP30P140LVT U139 ( .A1(n267), .A2(i_data_bus[103]), .B1(n266), .B2(
        i_data_bus[135]), .ZN(n112) );
  INVD1BWP30P140LVT U140 ( .I(i_data_bus[199]), .ZN(n108) );
  INVD1BWP30P140LVT U141 ( .I(i_data_bus[167]), .ZN(n107) );
  OAI22D1BWP30P140LVT U142 ( .A1(n289), .A2(n108), .B1(n287), .B2(n107), .ZN(
        n109) );
  AOI21D1BWP30P140LVT U143 ( .A1(n132), .A2(i_data_bus[231]), .B(n109), .ZN(
        n111) );
  ND2D1BWP30P140LVT U144 ( .A1(n3), .A2(i_data_bus[7]), .ZN(n110) );
  ND4D1BWP30P140LVT U145 ( .A1(n113), .A2(n112), .A3(n111), .A4(n110), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U146 ( .A1(n265), .A2(i_data_bus[70]), .B1(n264), .B2(
        i_data_bus[38]), .ZN(n120) );
  AOI22D1BWP30P140LVT U147 ( .A1(n267), .A2(i_data_bus[102]), .B1(n266), .B2(
        i_data_bus[134]), .ZN(n119) );
  INVD1BWP30P140LVT U148 ( .I(i_data_bus[198]), .ZN(n115) );
  INVD1BWP30P140LVT U149 ( .I(i_data_bus[166]), .ZN(n114) );
  OAI22D1BWP30P140LVT U150 ( .A1(n289), .A2(n115), .B1(n287), .B2(n114), .ZN(
        n116) );
  AOI21D1BWP30P140LVT U151 ( .A1(n132), .A2(i_data_bus[230]), .B(n116), .ZN(
        n118) );
  ND2D1BWP30P140LVT U152 ( .A1(n3), .A2(i_data_bus[6]), .ZN(n117) );
  ND4D1BWP30P140LVT U153 ( .A1(n120), .A2(n119), .A3(n118), .A4(n117), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U154 ( .A1(n146), .A2(i_data_bus[93]), .B1(n145), .B2(
        i_data_bus[61]), .ZN(n128) );
  AOI22D1BWP30P140LVT U155 ( .A1(n147), .A2(i_data_bus[125]), .B1(n284), .B2(
        i_data_bus[157]), .ZN(n127) );
  INVD1BWP30P140LVT U156 ( .I(i_data_bus[221]), .ZN(n123) );
  INVD1BWP30P140LVT U157 ( .I(i_data_bus[189]), .ZN(n122) );
  OAI22D1BWP30P140LVT U158 ( .A1(n2), .A2(n123), .B1(n226), .B2(n122), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U159 ( .A1(n132), .A2(i_data_bus[253]), .B(n124), .ZN(
        n126) );
  ND2D1BWP30P140LVT U160 ( .A1(n3), .A2(i_data_bus[29]), .ZN(n125) );
  ND4D1BWP30P140LVT U161 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U162 ( .A1(n146), .A2(i_data_bus[92]), .B1(n145), .B2(
        i_data_bus[60]), .ZN(n136) );
  AOI22D1BWP30P140LVT U163 ( .A1(n147), .A2(i_data_bus[124]), .B1(n284), .B2(
        i_data_bus[156]), .ZN(n135) );
  INVD1BWP30P140LVT U164 ( .I(i_data_bus[220]), .ZN(n130) );
  INVD1BWP30P140LVT U165 ( .I(i_data_bus[188]), .ZN(n129) );
  OAI22D1BWP30P140LVT U166 ( .A1(n2), .A2(n130), .B1(n226), .B2(n129), .ZN(
        n131) );
  AOI21D1BWP30P140LVT U167 ( .A1(n132), .A2(i_data_bus[252]), .B(n131), .ZN(
        n134) );
  ND2D1BWP30P140LVT U168 ( .A1(n3), .A2(i_data_bus[28]), .ZN(n133) );
  ND4D1BWP30P140LVT U169 ( .A1(n136), .A2(n135), .A3(n134), .A4(n133), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U170 ( .A1(n146), .A2(i_data_bus[91]), .B1(n145), .B2(
        i_data_bus[59]), .ZN(n144) );
  AOI22D1BWP30P140LVT U171 ( .A1(n147), .A2(i_data_bus[123]), .B1(n284), .B2(
        i_data_bus[155]), .ZN(n143) );
  INVD1BWP30P140LVT U172 ( .I(i_data_bus[219]), .ZN(n139) );
  INVD1BWP30P140LVT U173 ( .I(i_data_bus[187]), .ZN(n138) );
  OAI22D1BWP30P140LVT U174 ( .A1(n2), .A2(n139), .B1(n226), .B2(n138), .ZN(
        n140) );
  AOI21D1BWP30P140LVT U175 ( .A1(n132), .A2(i_data_bus[251]), .B(n140), .ZN(
        n142) );
  ND2D1BWP30P140LVT U176 ( .A1(n3), .A2(i_data_bus[27]), .ZN(n141) );
  ND4D1BWP30P140LVT U177 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U178 ( .A1(n146), .A2(i_data_bus[90]), .B1(n145), .B2(
        i_data_bus[58]), .ZN(n154) );
  AOI22D1BWP30P140LVT U179 ( .A1(n147), .A2(i_data_bus[122]), .B1(n284), .B2(
        i_data_bus[154]), .ZN(n153) );
  INVD1BWP30P140LVT U180 ( .I(i_data_bus[218]), .ZN(n149) );
  INVD1BWP30P140LVT U181 ( .I(i_data_bus[186]), .ZN(n148) );
  OAI22D1BWP30P140LVT U182 ( .A1(n2), .A2(n149), .B1(n226), .B2(n148), .ZN(
        n150) );
  AOI21D1BWP30P140LVT U183 ( .A1(n132), .A2(i_data_bus[250]), .B(n150), .ZN(
        n152) );
  ND2D1BWP30P140LVT U184 ( .A1(n3), .A2(i_data_bus[26]), .ZN(n151) );
  ND4D1BWP30P140LVT U185 ( .A1(n154), .A2(n153), .A3(n152), .A4(n151), .ZN(
        N395) );
  INVD2BWP30P140LVT U186 ( .I(n4), .ZN(n283) );
  INVD2BWP30P140LVT U187 ( .I(n155), .ZN(n156) );
  INVD2BWP30P140LVT U188 ( .I(n156), .ZN(n282) );
  AOI22D1BWP30P140LVT U189 ( .A1(n283), .A2(i_data_bus[89]), .B1(n282), .B2(
        i_data_bus[57]), .ZN(n165) );
  INVD2BWP30P140LVT U190 ( .I(n157), .ZN(n285) );
  AOI22D1BWP30P140LVT U191 ( .A1(n285), .A2(i_data_bus[121]), .B1(n284), .B2(
        i_data_bus[153]), .ZN(n164) );
  INVD1BWP30P140LVT U192 ( .I(i_data_bus[217]), .ZN(n159) );
  INVD1BWP30P140LVT U193 ( .I(i_data_bus[185]), .ZN(n158) );
  ND2D1BWP30P140LVT U194 ( .A1(n3), .A2(i_data_bus[25]), .ZN(n162) );
  ND4D1BWP30P140LVT U195 ( .A1(n165), .A2(n164), .A3(n163), .A4(n162), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U196 ( .A1(n283), .A2(i_data_bus[88]), .B1(n282), .B2(
        i_data_bus[56]), .ZN(n172) );
  AOI22D1BWP30P140LVT U197 ( .A1(n285), .A2(i_data_bus[120]), .B1(n284), .B2(
        i_data_bus[152]), .ZN(n171) );
  INVD1BWP30P140LVT U198 ( .I(i_data_bus[216]), .ZN(n167) );
  INVD1BWP30P140LVT U199 ( .I(i_data_bus[184]), .ZN(n166) );
  OAI22D1BWP30P140LVT U200 ( .A1(n289), .A2(n167), .B1(n226), .B2(n166), .ZN(
        n168) );
  AOI21D1BWP30P140LVT U201 ( .A1(n132), .A2(i_data_bus[248]), .B(n168), .ZN(
        n170) );
  ND2D1BWP30P140LVT U202 ( .A1(n3), .A2(i_data_bus[24]), .ZN(n169) );
  ND4D1BWP30P140LVT U203 ( .A1(n172), .A2(n171), .A3(n170), .A4(n169), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U204 ( .A1(n283), .A2(i_data_bus[87]), .B1(n282), .B2(
        i_data_bus[55]), .ZN(n179) );
  AOI22D1BWP30P140LVT U205 ( .A1(n285), .A2(i_data_bus[119]), .B1(n284), .B2(
        i_data_bus[151]), .ZN(n178) );
  INVD1BWP30P140LVT U206 ( .I(i_data_bus[215]), .ZN(n174) );
  INVD1BWP30P140LVT U207 ( .I(i_data_bus[183]), .ZN(n173) );
  OAI22D1BWP30P140LVT U208 ( .A1(n289), .A2(n174), .B1(n226), .B2(n173), .ZN(
        n175) );
  AOI21D1BWP30P140LVT U209 ( .A1(n132), .A2(i_data_bus[247]), .B(n175), .ZN(
        n177) );
  ND2D1BWP30P140LVT U210 ( .A1(n3), .A2(i_data_bus[23]), .ZN(n176) );
  ND4D1BWP30P140LVT U211 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U212 ( .A1(n283), .A2(i_data_bus[86]), .B1(n282), .B2(
        i_data_bus[54]), .ZN(n186) );
  AOI22D1BWP30P140LVT U213 ( .A1(n285), .A2(i_data_bus[118]), .B1(n284), .B2(
        i_data_bus[150]), .ZN(n185) );
  INVD1BWP30P140LVT U214 ( .I(i_data_bus[214]), .ZN(n181) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[182]), .ZN(n180) );
  OAI22D1BWP30P140LVT U216 ( .A1(n289), .A2(n181), .B1(n226), .B2(n180), .ZN(
        n182) );
  AOI21D1BWP30P140LVT U217 ( .A1(n132), .A2(i_data_bus[246]), .B(n182), .ZN(
        n184) );
  ND2D1BWP30P140LVT U218 ( .A1(n3), .A2(i_data_bus[22]), .ZN(n183) );
  ND4D1BWP30P140LVT U219 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U220 ( .A1(n283), .A2(i_data_bus[85]), .B1(n282), .B2(
        i_data_bus[53]), .ZN(n193) );
  AOI22D1BWP30P140LVT U221 ( .A1(n285), .A2(i_data_bus[117]), .B1(n284), .B2(
        i_data_bus[149]), .ZN(n192) );
  INVD1BWP30P140LVT U222 ( .I(i_data_bus[213]), .ZN(n188) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[181]), .ZN(n187) );
  OAI22D1BWP30P140LVT U224 ( .A1(n289), .A2(n188), .B1(n226), .B2(n187), .ZN(
        n189) );
  AOI21D1BWP30P140LVT U225 ( .A1(n132), .A2(i_data_bus[245]), .B(n189), .ZN(
        n191) );
  ND2D1BWP30P140LVT U226 ( .A1(n3), .A2(i_data_bus[21]), .ZN(n190) );
  ND4D1BWP30P140LVT U227 ( .A1(n193), .A2(n192), .A3(n191), .A4(n190), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U228 ( .A1(n283), .A2(i_data_bus[84]), .B1(n282), .B2(
        i_data_bus[52]), .ZN(n200) );
  AOI22D1BWP30P140LVT U229 ( .A1(n285), .A2(i_data_bus[116]), .B1(n284), .B2(
        i_data_bus[148]), .ZN(n199) );
  INVD1BWP30P140LVT U230 ( .I(i_data_bus[212]), .ZN(n195) );
  INVD1BWP30P140LVT U231 ( .I(i_data_bus[180]), .ZN(n194) );
  OAI22D1BWP30P140LVT U232 ( .A1(n289), .A2(n195), .B1(n226), .B2(n194), .ZN(
        n196) );
  AOI21D1BWP30P140LVT U233 ( .A1(n132), .A2(i_data_bus[244]), .B(n196), .ZN(
        n198) );
  ND2D1BWP30P140LVT U234 ( .A1(n3), .A2(i_data_bus[20]), .ZN(n197) );
  ND4D1BWP30P140LVT U235 ( .A1(n200), .A2(n199), .A3(n198), .A4(n197), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U236 ( .A1(n283), .A2(i_data_bus[83]), .B1(n282), .B2(
        i_data_bus[51]), .ZN(n206) );
  AOI22D1BWP30P140LVT U237 ( .A1(n285), .A2(i_data_bus[115]), .B1(n284), .B2(
        i_data_bus[147]), .ZN(n205) );
  INVD1BWP30P140LVT U238 ( .I(i_data_bus[179]), .ZN(n201) );
  MOAI22D1BWP30P140LVT U239 ( .A1(n226), .A2(n201), .B1(n275), .B2(
        i_data_bus[211]), .ZN(n202) );
  AOI21D1BWP30P140LVT U240 ( .A1(n132), .A2(i_data_bus[243]), .B(n202), .ZN(
        n204) );
  ND2D1BWP30P140LVT U241 ( .A1(n3), .A2(i_data_bus[19]), .ZN(n203) );
  ND4D1BWP30P140LVT U242 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U243 ( .A1(n283), .A2(i_data_bus[82]), .B1(n282), .B2(
        i_data_bus[50]), .ZN(n212) );
  AOI22D1BWP30P140LVT U244 ( .A1(n285), .A2(i_data_bus[114]), .B1(n284), .B2(
        i_data_bus[146]), .ZN(n211) );
  INVD1BWP30P140LVT U245 ( .I(i_data_bus[178]), .ZN(n207) );
  MOAI22D1BWP30P140LVT U246 ( .A1(n226), .A2(n207), .B1(n275), .B2(
        i_data_bus[210]), .ZN(n208) );
  AOI21D1BWP30P140LVT U247 ( .A1(n132), .A2(i_data_bus[242]), .B(n208), .ZN(
        n210) );
  ND2D1BWP30P140LVT U248 ( .A1(n3), .A2(i_data_bus[18]), .ZN(n209) );
  ND4D1BWP30P140LVT U249 ( .A1(n212), .A2(n211), .A3(n210), .A4(n209), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U250 ( .A1(n283), .A2(i_data_bus[81]), .B1(n282), .B2(
        i_data_bus[49]), .ZN(n218) );
  AOI22D1BWP30P140LVT U251 ( .A1(n285), .A2(i_data_bus[113]), .B1(n284), .B2(
        i_data_bus[145]), .ZN(n217) );
  INVD1BWP30P140LVT U252 ( .I(i_data_bus[177]), .ZN(n213) );
  MOAI22D1BWP30P140LVT U253 ( .A1(n226), .A2(n213), .B1(n275), .B2(
        i_data_bus[209]), .ZN(n214) );
  AOI21D1BWP30P140LVT U254 ( .A1(n132), .A2(i_data_bus[241]), .B(n214), .ZN(
        n216) );
  ND2D1BWP30P140LVT U255 ( .A1(n3), .A2(i_data_bus[17]), .ZN(n215) );
  ND4D1BWP30P140LVT U256 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U257 ( .A1(n283), .A2(i_data_bus[80]), .B1(n282), .B2(
        i_data_bus[48]), .ZN(n224) );
  AOI22D1BWP30P140LVT U258 ( .A1(n285), .A2(i_data_bus[112]), .B1(n284), .B2(
        i_data_bus[144]), .ZN(n223) );
  INVD1BWP30P140LVT U259 ( .I(i_data_bus[176]), .ZN(n219) );
  MOAI22D1BWP30P140LVT U260 ( .A1(n226), .A2(n219), .B1(n275), .B2(
        i_data_bus[208]), .ZN(n220) );
  AOI21D1BWP30P140LVT U261 ( .A1(n132), .A2(i_data_bus[240]), .B(n220), .ZN(
        n222) );
  ND2D1BWP30P140LVT U262 ( .A1(n3), .A2(i_data_bus[16]), .ZN(n221) );
  ND4D1BWP30P140LVT U263 ( .A1(n224), .A2(n223), .A3(n222), .A4(n221), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U264 ( .A1(n283), .A2(i_data_bus[79]), .B1(n282), .B2(
        i_data_bus[47]), .ZN(n231) );
  AOI22D1BWP30P140LVT U265 ( .A1(n285), .A2(i_data_bus[111]), .B1(n284), .B2(
        i_data_bus[143]), .ZN(n230) );
  INVD1BWP30P140LVT U266 ( .I(i_data_bus[175]), .ZN(n225) );
  MOAI22D1BWP30P140LVT U267 ( .A1(n226), .A2(n225), .B1(n275), .B2(
        i_data_bus[207]), .ZN(n227) );
  AOI21D1BWP30P140LVT U268 ( .A1(n132), .A2(i_data_bus[239]), .B(n227), .ZN(
        n229) );
  ND2D1BWP30P140LVT U269 ( .A1(n3), .A2(i_data_bus[15]), .ZN(n228) );
  ND4D1BWP30P140LVT U270 ( .A1(n231), .A2(n230), .A3(n229), .A4(n228), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U271 ( .A1(n265), .A2(i_data_bus[68]), .B1(n264), .B2(
        i_data_bus[36]), .ZN(n238) );
  AOI22D1BWP30P140LVT U272 ( .A1(n267), .A2(i_data_bus[100]), .B1(n266), .B2(
        i_data_bus[132]), .ZN(n237) );
  INVD1BWP30P140LVT U273 ( .I(i_data_bus[196]), .ZN(n233) );
  INVD1BWP30P140LVT U274 ( .I(i_data_bus[164]), .ZN(n232) );
  OAI22D1BWP30P140LVT U275 ( .A1(n289), .A2(n233), .B1(n287), .B2(n232), .ZN(
        n234) );
  AOI21D1BWP30P140LVT U276 ( .A1(n132), .A2(i_data_bus[228]), .B(n234), .ZN(
        n236) );
  ND2D1BWP30P140LVT U277 ( .A1(n3), .A2(i_data_bus[4]), .ZN(n235) );
  ND4D1BWP30P140LVT U278 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U279 ( .A1(n265), .A2(i_data_bus[67]), .B1(n264), .B2(
        i_data_bus[35]), .ZN(n245) );
  AOI22D1BWP30P140LVT U280 ( .A1(n267), .A2(i_data_bus[99]), .B1(n266), .B2(
        i_data_bus[131]), .ZN(n244) );
  INVD1BWP30P140LVT U281 ( .I(i_data_bus[195]), .ZN(n240) );
  INVD1BWP30P140LVT U282 ( .I(i_data_bus[163]), .ZN(n239) );
  OAI22D1BWP30P140LVT U283 ( .A1(n289), .A2(n240), .B1(n287), .B2(n239), .ZN(
        n241) );
  AOI21D1BWP30P140LVT U284 ( .A1(n132), .A2(i_data_bus[227]), .B(n241), .ZN(
        n243) );
  ND2D1BWP30P140LVT U285 ( .A1(n3), .A2(i_data_bus[3]), .ZN(n242) );
  ND4D1BWP30P140LVT U286 ( .A1(n245), .A2(n244), .A3(n243), .A4(n242), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U287 ( .A1(n265), .A2(i_data_bus[66]), .B1(n264), .B2(
        i_data_bus[34]), .ZN(n251) );
  AOI22D1BWP30P140LVT U288 ( .A1(n267), .A2(i_data_bus[98]), .B1(n266), .B2(
        i_data_bus[130]), .ZN(n250) );
  INVD1BWP30P140LVT U289 ( .I(i_data_bus[162]), .ZN(n246) );
  MOAI22D1BWP30P140LVT U290 ( .A1(n287), .A2(n246), .B1(n275), .B2(
        i_data_bus[194]), .ZN(n247) );
  AOI21D1BWP30P140LVT U291 ( .A1(n132), .A2(i_data_bus[226]), .B(n247), .ZN(
        n249) );
  ND2D1BWP30P140LVT U292 ( .A1(n3), .A2(i_data_bus[2]), .ZN(n248) );
  ND4D1BWP30P140LVT U293 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U294 ( .A1(n265), .A2(i_data_bus[72]), .B1(n264), .B2(
        i_data_bus[40]), .ZN(n257) );
  AOI22D1BWP30P140LVT U295 ( .A1(n267), .A2(i_data_bus[104]), .B1(n266), .B2(
        i_data_bus[136]), .ZN(n256) );
  INVD1BWP30P140LVT U296 ( .I(i_data_bus[168]), .ZN(n252) );
  MOAI22D1BWP30P140LVT U297 ( .A1(n287), .A2(n252), .B1(n275), .B2(
        i_data_bus[200]), .ZN(n253) );
  AOI21D1BWP30P140LVT U298 ( .A1(n132), .A2(i_data_bus[232]), .B(n253), .ZN(
        n255) );
  ND2D1BWP30P140LVT U299 ( .A1(n3), .A2(i_data_bus[8]), .ZN(n254) );
  ND4D1BWP30P140LVT U300 ( .A1(n257), .A2(n256), .A3(n255), .A4(n254), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U301 ( .A1(n265), .A2(i_data_bus[64]), .B1(n264), .B2(
        i_data_bus[32]), .ZN(n263) );
  AOI22D1BWP30P140LVT U302 ( .A1(n267), .A2(i_data_bus[96]), .B1(n266), .B2(
        i_data_bus[128]), .ZN(n262) );
  INR2D1BWP30P140LVT U303 ( .A1(i_data_bus[192]), .B1(n289), .ZN(n259) );
  INR2D1BWP30P140LVT U304 ( .A1(i_data_bus[160]), .B1(n287), .ZN(n258) );
  AOI211D1BWP30P140LVT U305 ( .A1(i_data_bus[224]), .A2(n132), .B(n259), .C(
        n258), .ZN(n261) );
  ND2D1BWP30P140LVT U306 ( .A1(n3), .A2(i_data_bus[0]), .ZN(n260) );
  ND4D1BWP30P140LVT U307 ( .A1(n263), .A2(n262), .A3(n261), .A4(n260), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U308 ( .A1(n265), .A2(i_data_bus[65]), .B1(n264), .B2(
        i_data_bus[33]), .ZN(n274) );
  AOI22D1BWP30P140LVT U309 ( .A1(n267), .A2(i_data_bus[97]), .B1(n266), .B2(
        i_data_bus[129]), .ZN(n273) );
  INVD1BWP30P140LVT U310 ( .I(i_data_bus[161]), .ZN(n269) );
  OAI21D1BWP30P140LVT U311 ( .A1(n287), .A2(n269), .B(n268), .ZN(n270) );
  AOI21D1BWP30P140LVT U312 ( .A1(n132), .A2(i_data_bus[225]), .B(n270), .ZN(
        n272) );
  ND2D1BWP30P140LVT U313 ( .A1(n3), .A2(i_data_bus[1]), .ZN(n271) );
  ND4D1BWP30P140LVT U314 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U315 ( .A1(n283), .A2(i_data_bus[78]), .B1(n282), .B2(
        i_data_bus[46]), .ZN(n281) );
  AOI22D1BWP30P140LVT U316 ( .A1(n285), .A2(i_data_bus[110]), .B1(n284), .B2(
        i_data_bus[142]), .ZN(n280) );
  INVD1BWP30P140LVT U317 ( .I(i_data_bus[174]), .ZN(n276) );
  MOAI22D1BWP30P140LVT U318 ( .A1(n287), .A2(n276), .B1(n275), .B2(
        i_data_bus[206]), .ZN(n277) );
  AOI21D1BWP30P140LVT U319 ( .A1(n132), .A2(i_data_bus[238]), .B(n277), .ZN(
        n279) );
  ND2D1BWP30P140LVT U320 ( .A1(n3), .A2(i_data_bus[14]), .ZN(n278) );
  ND4D1BWP30P140LVT U321 ( .A1(n281), .A2(n280), .A3(n279), .A4(n278), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U322 ( .A1(n283), .A2(i_data_bus[77]), .B1(n282), .B2(
        i_data_bus[45]), .ZN(n294) );
  AOI22D1BWP30P140LVT U323 ( .A1(n285), .A2(i_data_bus[109]), .B1(n284), .B2(
        i_data_bus[141]), .ZN(n293) );
  INVD1BWP30P140LVT U324 ( .I(i_data_bus[205]), .ZN(n288) );
  INVD1BWP30P140LVT U325 ( .I(i_data_bus[173]), .ZN(n286) );
  OAI22D1BWP30P140LVT U326 ( .A1(n289), .A2(n288), .B1(n287), .B2(n286), .ZN(
        n290) );
  AOI21D1BWP30P140LVT U327 ( .A1(n132), .A2(i_data_bus[237]), .B(n290), .ZN(
        n292) );
  ND2D1BWP30P140LVT U328 ( .A1(n3), .A2(i_data_bus[13]), .ZN(n291) );
  ND4D1BWP30P140LVT U329 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_5 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n113), .ZN(n4) );
  INVD1BWP30P140LVT U4 ( .I(n21), .ZN(n63) );
  CKND2D3BWP30P140LVT U5 ( .A1(n12), .A2(n18), .ZN(n55) );
  CKND2D2BWP30P140LVT U6 ( .A1(n11), .A2(n23), .ZN(n37) );
  AOI22D1BWP30P140LVT U7 ( .A1(n265), .A2(i_data_bus[72]), .B1(n264), .B2(
        i_data_bus[40]), .ZN(n244) );
  AOI21D1BWP30P140LVT U8 ( .A1(n1), .A2(i_data_bus[243]), .B(n159), .ZN(n161)
         );
  AN2D2BWP30P140LVT U9 ( .A1(n32), .A2(n40), .Z(n1) );
  INVD1BWP30P140LVT U10 ( .I(n5), .ZN(n6) );
  ND2D1BWP30P140LVT U11 ( .A1(n241), .A2(n244), .ZN(n5) );
  INVD2BWP30P140LVT U12 ( .I(n82), .ZN(n2) );
  INVD6BWP30P140LVT U13 ( .I(n274), .ZN(n3) );
  NR2OPTPAD2BWP30P140LVT U14 ( .A1(n37), .A2(i_cmd[5]), .ZN(n18) );
  INVD2BWP30P140LVT U15 ( .I(n63), .ZN(n266) );
  INVD3BWP30P140LVT U16 ( .I(n63), .ZN(n283) );
  ND3D1BWP30P140LVT U17 ( .A1(n242), .A2(n243), .A3(n6), .ZN(N377) );
  INVD3BWP30P140LVT U18 ( .I(n42), .ZN(n285) );
  INVD2BWP30P140LVT U19 ( .I(i_cmd[4]), .ZN(n28) );
  OR2D1BWP30P140LVT U20 ( .A1(n55), .A2(n15), .Z(n113) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n18), .A2(n17), .Z(n7) );
  INVD1BWP30P140LVT U22 ( .I(rst), .ZN(n8) );
  ND2D1BWP30P140LVT U23 ( .A1(n8), .A2(i_en), .ZN(n25) );
  OR2D1BWP30P140LVT U24 ( .A1(i_cmd[0]), .A2(n25), .Z(n10) );
  INVD1BWP30P140LVT U25 ( .I(n28), .ZN(n9) );
  NR2OPTPAD1BWP30P140LVT U26 ( .A1(n10), .A2(n9), .ZN(n12) );
  INVD2BWP30P140LVT U27 ( .I(i_cmd[6]), .ZN(n11) );
  INVD2BWP30P140LVT U28 ( .I(i_cmd[7]), .ZN(n23) );
  INVD2BWP30P140LVT U29 ( .I(i_cmd[2]), .ZN(n51) );
  INVD2BWP30P140LVT U30 ( .I(i_cmd[1]), .ZN(n13) );
  ND2OPTIBD2BWP30P140LVT U31 ( .A1(n51), .A2(n13), .ZN(n24) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n14) );
  OR2D1BWP30P140LVT U33 ( .A1(n24), .A2(n14), .Z(n15) );
  ND2OPTIBD1BWP30P140LVT U34 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n16) );
  NR2D1BWP30P140LVT U35 ( .A1(n16), .A2(i_cmd[0]), .ZN(n20) );
  INVD1BWP30P140LVT U36 ( .I(n25), .ZN(n17) );
  OR2D1BWP30P140LVT U37 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n54) );
  NR2D1BWP30P140LVT U38 ( .A1(n54), .A2(i_cmd[1]), .ZN(n19) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(n7), .A2(n19), .ZN(n46) );
  INR2D1BWP30P140LVT U40 ( .A1(n20), .B1(n46), .ZN(n21) );
  AOI22D1BWP30P140LVT U41 ( .A1(n4), .A2(i_data_bus[96]), .B1(n266), .B2(
        i_data_bus[128]), .ZN(n62) );
  INVD1BWP30P140LVT U42 ( .I(i_valid[7]), .ZN(n22) );
  NR4D0BWP30P140LVT U43 ( .A1(n23), .A2(n22), .A3(i_cmd[6]), .A4(i_cmd[5]), 
        .ZN(n32) );
  INVD1BWP30P140LVT U44 ( .I(n24), .ZN(n27) );
  NR2OPTPAD1BWP30P140LVT U45 ( .A1(i_cmd[0]), .A2(n25), .ZN(n26) );
  ND2OPTIBD2BWP30P140LVT U46 ( .A1(n27), .A2(n26), .ZN(n31) );
  INVD1BWP30P140LVT U47 ( .I(i_cmd[3]), .ZN(n29) );
  ND2OPTIBD1BWP30P140LVT U48 ( .A1(n29), .A2(n28), .ZN(n30) );
  NR2D3BWP30P140LVT U49 ( .A1(n31), .A2(n30), .ZN(n40) );
  NR2D1BWP30P140LVT U50 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n34) );
  CKAN2D1BWP30P140LVT U51 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n33) );
  ND2D1BWP30P140LVT U52 ( .A1(n34), .A2(n33), .ZN(n35) );
  INVD1BWP30P140LVT U53 ( .I(n35), .ZN(n36) );
  CKAN2D4BWP30P140LVT U54 ( .A1(n36), .A2(n40), .Z(n274) );
  INR2D1BWP30P140LVT U55 ( .A1(i_data_bus[192]), .B1(n3), .ZN(n44) );
  INVD1BWP30P140LVT U56 ( .I(n37), .ZN(n39) );
  ND2OPTIBD1BWP30P140LVT U57 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n38) );
  INR2D1BWP30P140LVT U58 ( .A1(n39), .B1(n38), .ZN(n41) );
  ND2OPTIBD2BWP30P140LVT U59 ( .A1(n41), .A2(n40), .ZN(n82) );
  INVD2BWP30P140LVT U60 ( .I(n82), .ZN(n42) );
  INR2D1BWP30P140LVT U61 ( .A1(i_data_bus[160]), .B1(n285), .ZN(n43) );
  AOI211D1BWP30P140LVT U62 ( .A1(i_data_bus[224]), .A2(n1), .B(n44), .C(n43), 
        .ZN(n61) );
  INVD1BWP30P140LVT U63 ( .I(i_cmd[0]), .ZN(n45) );
  INR3D0BWP30P140LVT U64 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n45), .ZN(n47)
         );
  INR2D1BWP30P140LVT U65 ( .A1(n47), .B1(n46), .ZN(n48) );
  INVD2BWP30P140LVT U66 ( .I(n48), .ZN(n117) );
  INVD3BWP30P140LVT U67 ( .I(n117), .ZN(n269) );
  ND2D1BWP30P140LVT U68 ( .A1(n269), .A2(i_data_bus[0]), .ZN(n58) );
  OR2D1BWP30P140LVT U69 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .Z(n50) );
  INVD1BWP30P140LVT U70 ( .I(i_valid[2]), .ZN(n49) );
  OR3D1BWP30P140LVT U71 ( .A1(n51), .A2(n50), .A3(n49), .Z(n52) );
  OR2D4BWP30P140LVT U72 ( .A1(n52), .A2(n55), .Z(n72) );
  INVD3BWP30P140LVT U73 ( .I(n72), .ZN(n265) );
  ND2D1BWP30P140LVT U74 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n53) );
  NR2D1BWP30P140LVT U75 ( .A1(n54), .A2(n53), .ZN(n56) );
  INR2D6BWP30P140LVT U76 ( .A1(n56), .B1(n55), .ZN(n264) );
  AOI22D1BWP30P140LVT U77 ( .A1(n265), .A2(i_data_bus[64]), .B1(n264), .B2(
        i_data_bus[32]), .ZN(n57) );
  ND2D1BWP30P140LVT U78 ( .A1(n58), .A2(n57), .ZN(n59) );
  INVD1BWP30P140LVT U79 ( .I(n59), .ZN(n60) );
  ND3D1BWP30P140LVT U80 ( .A1(n62), .A2(n61), .A3(n60), .ZN(N369) );
  INVD2BWP30P140LVT U81 ( .I(n72), .ZN(n282) );
  AOI22D1BWP30P140LVT U82 ( .A1(n282), .A2(i_data_bus[94]), .B1(n264), .B2(
        i_data_bus[62]), .ZN(n70) );
  AOI22D1BWP30P140LVT U83 ( .A1(n4), .A2(i_data_bus[126]), .B1(n283), .B2(
        i_data_bus[158]), .ZN(n69) );
  INVD1BWP30P140LVT U84 ( .I(i_data_bus[222]), .ZN(n65) );
  INVD1BWP30P140LVT U85 ( .I(i_data_bus[190]), .ZN(n64) );
  OAI22D1BWP30P140LVT U86 ( .A1(n3), .A2(n65), .B1(n82), .B2(n64), .ZN(n66) );
  AOI21D1BWP30P140LVT U87 ( .A1(n1), .A2(i_data_bus[254]), .B(n66), .ZN(n68)
         );
  INVD1BWP30P140LVT U88 ( .I(n117), .ZN(n107) );
  ND2D1BWP30P140LVT U89 ( .A1(n107), .A2(i_data_bus[30]), .ZN(n67) );
  ND4D1BWP30P140LVT U90 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(N399) );
  NR4D0BWP30P140LVT U91 ( .A1(n107), .A2(n274), .A3(n2), .A4(n1), .ZN(n74) );
  NR2D1BWP30P140LVT U92 ( .A1(n4), .A2(n283), .ZN(n73) );
  INVD1BWP30P140LVT U93 ( .I(n264), .ZN(n71) );
  ND4D1BWP30P140LVT U94 ( .A1(n74), .A2(n73), .A3(n72), .A4(n71), .ZN(N402) );
  AOI22D1BWP30P140LVT U95 ( .A1(n282), .A2(i_data_bus[95]), .B1(n264), .B2(
        i_data_bus[63]), .ZN(n81) );
  AOI22D1BWP30P140LVT U96 ( .A1(n4), .A2(i_data_bus[127]), .B1(n283), .B2(
        i_data_bus[159]), .ZN(n80) );
  INVD1BWP30P140LVT U97 ( .I(i_data_bus[223]), .ZN(n76) );
  INVD1BWP30P140LVT U98 ( .I(i_data_bus[191]), .ZN(n75) );
  OAI22D1BWP30P140LVT U99 ( .A1(n3), .A2(n76), .B1(n82), .B2(n75), .ZN(n77) );
  AOI21D1BWP30P140LVT U100 ( .A1(n1), .A2(i_data_bus[255]), .B(n77), .ZN(n79)
         );
  ND2D1BWP30P140LVT U101 ( .A1(n107), .A2(i_data_bus[31]), .ZN(n78) );
  ND4D1BWP30P140LVT U102 ( .A1(n81), .A2(n80), .A3(n79), .A4(n78), .ZN(N400)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n282), .A2(i_data_bus[93]), .B1(n264), .B2(
        i_data_bus[61]), .ZN(n89) );
  AOI22D1BWP30P140LVT U104 ( .A1(n4), .A2(i_data_bus[125]), .B1(n283), .B2(
        i_data_bus[157]), .ZN(n88) );
  INVD1BWP30P140LVT U105 ( .I(i_data_bus[221]), .ZN(n84) );
  INVD3BWP30P140LVT U106 ( .I(n2), .ZN(n183) );
  INVD1BWP30P140LVT U107 ( .I(i_data_bus[189]), .ZN(n83) );
  OAI22D1BWP30P140LVT U108 ( .A1(n3), .A2(n84), .B1(n183), .B2(n83), .ZN(n85)
         );
  AOI21D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[253]), .B(n85), .ZN(n87)
         );
  ND2D1BWP30P140LVT U110 ( .A1(n107), .A2(i_data_bus[29]), .ZN(n86) );
  ND4D1BWP30P140LVT U111 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(N398)
         );
  AOI22D1BWP30P140LVT U112 ( .A1(n282), .A2(i_data_bus[92]), .B1(n264), .B2(
        i_data_bus[60]), .ZN(n96) );
  AOI22D1BWP30P140LVT U113 ( .A1(n4), .A2(i_data_bus[124]), .B1(n283), .B2(
        i_data_bus[156]), .ZN(n95) );
  INVD1BWP30P140LVT U114 ( .I(i_data_bus[220]), .ZN(n91) );
  INVD1BWP30P140LVT U115 ( .I(i_data_bus[188]), .ZN(n90) );
  OAI22D1BWP30P140LVT U116 ( .A1(n3), .A2(n91), .B1(n183), .B2(n90), .ZN(n92)
         );
  AOI21D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[252]), .B(n92), .ZN(n94)
         );
  ND2D1BWP30P140LVT U118 ( .A1(n107), .A2(i_data_bus[28]), .ZN(n93) );
  ND4D1BWP30P140LVT U119 ( .A1(n96), .A2(n95), .A3(n94), .A4(n93), .ZN(N397)
         );
  AOI22D1BWP30P140LVT U120 ( .A1(n282), .A2(i_data_bus[91]), .B1(n264), .B2(
        i_data_bus[59]), .ZN(n103) );
  AOI22D1BWP30P140LVT U121 ( .A1(n4), .A2(i_data_bus[123]), .B1(n283), .B2(
        i_data_bus[155]), .ZN(n102) );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[219]), .ZN(n98) );
  INVD1BWP30P140LVT U123 ( .I(i_data_bus[187]), .ZN(n97) );
  OAI22D1BWP30P140LVT U124 ( .A1(n3), .A2(n98), .B1(n183), .B2(n97), .ZN(n99)
         );
  AOI21D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[251]), .B(n99), .ZN(n101)
         );
  ND2D1BWP30P140LVT U126 ( .A1(n107), .A2(i_data_bus[27]), .ZN(n100) );
  ND4D1BWP30P140LVT U127 ( .A1(n103), .A2(n102), .A3(n101), .A4(n100), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U128 ( .A1(n282), .A2(i_data_bus[90]), .B1(n264), .B2(
        i_data_bus[58]), .ZN(n111) );
  AOI22D1BWP30P140LVT U129 ( .A1(n4), .A2(i_data_bus[122]), .B1(n283), .B2(
        i_data_bus[154]), .ZN(n110) );
  INVD1BWP30P140LVT U130 ( .I(i_data_bus[218]), .ZN(n105) );
  INVD1BWP30P140LVT U131 ( .I(i_data_bus[186]), .ZN(n104) );
  OAI22D1BWP30P140LVT U132 ( .A1(n3), .A2(n105), .B1(n183), .B2(n104), .ZN(
        n106) );
  AOI21D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[250]), .B(n106), .ZN(n109) );
  ND2D1BWP30P140LVT U134 ( .A1(n107), .A2(i_data_bus[26]), .ZN(n108) );
  ND4D1BWP30P140LVT U135 ( .A1(n111), .A2(n110), .A3(n109), .A4(n108), .ZN(
        N395) );
  INVD2BWP30P140LVT U136 ( .I(n264), .ZN(n112) );
  INVD2BWP30P140LVT U137 ( .I(n112), .ZN(n281) );
  AOI22D1BWP30P140LVT U138 ( .A1(n282), .A2(i_data_bus[89]), .B1(n281), .B2(
        i_data_bus[57]), .ZN(n121) );
  AOI22D1BWP30P140LVT U139 ( .A1(n4), .A2(i_data_bus[121]), .B1(n283), .B2(
        i_data_bus[153]), .ZN(n120) );
  INVD1BWP30P140LVT U140 ( .I(i_data_bus[217]), .ZN(n115) );
  INVD1BWP30P140LVT U141 ( .I(i_data_bus[185]), .ZN(n114) );
  OAI22D1BWP30P140LVT U142 ( .A1(n3), .A2(n115), .B1(n183), .B2(n114), .ZN(
        n116) );
  AOI21D1BWP30P140LVT U143 ( .A1(n1), .A2(i_data_bus[249]), .B(n116), .ZN(n119) );
  INVD2BWP30P140LVT U144 ( .I(n117), .ZN(n288) );
  ND2D1BWP30P140LVT U145 ( .A1(n288), .A2(i_data_bus[25]), .ZN(n118) );
  ND4D1BWP30P140LVT U146 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U147 ( .A1(n282), .A2(i_data_bus[88]), .B1(n281), .B2(
        i_data_bus[56]), .ZN(n128) );
  AOI22D1BWP30P140LVT U148 ( .A1(n4), .A2(i_data_bus[120]), .B1(n283), .B2(
        i_data_bus[152]), .ZN(n127) );
  INVD1BWP30P140LVT U149 ( .I(i_data_bus[216]), .ZN(n123) );
  INVD1BWP30P140LVT U150 ( .I(i_data_bus[184]), .ZN(n122) );
  OAI22D1BWP30P140LVT U151 ( .A1(n3), .A2(n123), .B1(n183), .B2(n122), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U152 ( .A1(n1), .A2(i_data_bus[248]), .B(n124), .ZN(n126) );
  ND2D1BWP30P140LVT U153 ( .A1(n288), .A2(i_data_bus[24]), .ZN(n125) );
  ND4D1BWP30P140LVT U154 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U155 ( .A1(n282), .A2(i_data_bus[87]), .B1(n281), .B2(
        i_data_bus[55]), .ZN(n135) );
  AOI22D1BWP30P140LVT U156 ( .A1(n4), .A2(i_data_bus[119]), .B1(n283), .B2(
        i_data_bus[151]), .ZN(n134) );
  INVD1BWP30P140LVT U157 ( .I(i_data_bus[215]), .ZN(n130) );
  INVD1BWP30P140LVT U158 ( .I(i_data_bus[183]), .ZN(n129) );
  OAI22D1BWP30P140LVT U159 ( .A1(n3), .A2(n130), .B1(n183), .B2(n129), .ZN(
        n131) );
  AOI21D1BWP30P140LVT U160 ( .A1(n1), .A2(i_data_bus[247]), .B(n131), .ZN(n133) );
  ND2D1BWP30P140LVT U161 ( .A1(n288), .A2(i_data_bus[23]), .ZN(n132) );
  ND4D1BWP30P140LVT U162 ( .A1(n135), .A2(n134), .A3(n133), .A4(n132), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U163 ( .A1(n282), .A2(i_data_bus[86]), .B1(n281), .B2(
        i_data_bus[54]), .ZN(n142) );
  AOI22D1BWP30P140LVT U164 ( .A1(n4), .A2(i_data_bus[118]), .B1(n283), .B2(
        i_data_bus[150]), .ZN(n141) );
  INVD1BWP30P140LVT U165 ( .I(i_data_bus[214]), .ZN(n137) );
  INVD1BWP30P140LVT U166 ( .I(i_data_bus[182]), .ZN(n136) );
  OAI22D1BWP30P140LVT U167 ( .A1(n3), .A2(n137), .B1(n183), .B2(n136), .ZN(
        n138) );
  AOI21D1BWP30P140LVT U168 ( .A1(n1), .A2(i_data_bus[246]), .B(n138), .ZN(n140) );
  ND2D1BWP30P140LVT U169 ( .A1(n288), .A2(i_data_bus[22]), .ZN(n139) );
  ND4D1BWP30P140LVT U170 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U171 ( .A1(n282), .A2(i_data_bus[85]), .B1(n281), .B2(
        i_data_bus[53]), .ZN(n149) );
  AOI22D1BWP30P140LVT U172 ( .A1(n4), .A2(i_data_bus[117]), .B1(n283), .B2(
        i_data_bus[149]), .ZN(n148) );
  INVD1BWP30P140LVT U173 ( .I(i_data_bus[213]), .ZN(n144) );
  INVD1BWP30P140LVT U174 ( .I(i_data_bus[181]), .ZN(n143) );
  OAI22D1BWP30P140LVT U175 ( .A1(n3), .A2(n144), .B1(n183), .B2(n143), .ZN(
        n145) );
  AOI21D1BWP30P140LVT U176 ( .A1(n1), .A2(i_data_bus[245]), .B(n145), .ZN(n147) );
  ND2D1BWP30P140LVT U177 ( .A1(n288), .A2(i_data_bus[21]), .ZN(n146) );
  ND4D1BWP30P140LVT U178 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U179 ( .A1(n282), .A2(i_data_bus[84]), .B1(n281), .B2(
        i_data_bus[52]), .ZN(n156) );
  AOI22D1BWP30P140LVT U180 ( .A1(n4), .A2(i_data_bus[116]), .B1(n283), .B2(
        i_data_bus[148]), .ZN(n155) );
  INVD1BWP30P140LVT U181 ( .I(i_data_bus[212]), .ZN(n151) );
  INVD1BWP30P140LVT U182 ( .I(i_data_bus[180]), .ZN(n150) );
  OAI22D1BWP30P140LVT U183 ( .A1(n3), .A2(n151), .B1(n183), .B2(n150), .ZN(
        n152) );
  AOI21D1BWP30P140LVT U184 ( .A1(n1), .A2(i_data_bus[244]), .B(n152), .ZN(n154) );
  ND2D1BWP30P140LVT U185 ( .A1(n288), .A2(i_data_bus[20]), .ZN(n153) );
  ND4D1BWP30P140LVT U186 ( .A1(n156), .A2(n155), .A3(n154), .A4(n153), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U187 ( .A1(n282), .A2(i_data_bus[83]), .B1(n281), .B2(
        i_data_bus[51]), .ZN(n163) );
  AOI22D1BWP30P140LVT U188 ( .A1(n4), .A2(i_data_bus[115]), .B1(n283), .B2(
        i_data_bus[147]), .ZN(n162) );
  INVD1BWP30P140LVT U189 ( .I(i_data_bus[211]), .ZN(n158) );
  INVD1BWP30P140LVT U190 ( .I(i_data_bus[179]), .ZN(n157) );
  OAI22D1BWP30P140LVT U191 ( .A1(n3), .A2(n158), .B1(n183), .B2(n157), .ZN(
        n159) );
  ND2D1BWP30P140LVT U192 ( .A1(n288), .A2(i_data_bus[19]), .ZN(n160) );
  ND4D1BWP30P140LVT U193 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U194 ( .A1(n282), .A2(i_data_bus[82]), .B1(n281), .B2(
        i_data_bus[50]), .ZN(n169) );
  AOI22D1BWP30P140LVT U195 ( .A1(n4), .A2(i_data_bus[114]), .B1(n283), .B2(
        i_data_bus[146]), .ZN(n168) );
  INVD1BWP30P140LVT U196 ( .I(i_data_bus[178]), .ZN(n164) );
  MOAI22D1BWP30P140LVT U197 ( .A1(n183), .A2(n164), .B1(n274), .B2(
        i_data_bus[210]), .ZN(n165) );
  AOI21D1BWP30P140LVT U198 ( .A1(n1), .A2(i_data_bus[242]), .B(n165), .ZN(n167) );
  ND2D1BWP30P140LVT U199 ( .A1(n288), .A2(i_data_bus[18]), .ZN(n166) );
  ND4D1BWP30P140LVT U200 ( .A1(n169), .A2(n168), .A3(n167), .A4(n166), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U201 ( .A1(n282), .A2(i_data_bus[81]), .B1(n281), .B2(
        i_data_bus[49]), .ZN(n175) );
  AOI22D1BWP30P140LVT U202 ( .A1(n4), .A2(i_data_bus[113]), .B1(n283), .B2(
        i_data_bus[145]), .ZN(n174) );
  INVD1BWP30P140LVT U203 ( .I(i_data_bus[177]), .ZN(n170) );
  MOAI22D1BWP30P140LVT U204 ( .A1(n183), .A2(n170), .B1(n274), .B2(
        i_data_bus[209]), .ZN(n171) );
  AOI21D1BWP30P140LVT U205 ( .A1(n1), .A2(i_data_bus[241]), .B(n171), .ZN(n173) );
  ND2D1BWP30P140LVT U206 ( .A1(n288), .A2(i_data_bus[17]), .ZN(n172) );
  ND4D1BWP30P140LVT U207 ( .A1(n175), .A2(n174), .A3(n173), .A4(n172), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U208 ( .A1(n282), .A2(i_data_bus[80]), .B1(n281), .B2(
        i_data_bus[48]), .ZN(n181) );
  AOI22D1BWP30P140LVT U209 ( .A1(n4), .A2(i_data_bus[112]), .B1(n283), .B2(
        i_data_bus[144]), .ZN(n180) );
  INVD1BWP30P140LVT U210 ( .I(i_data_bus[176]), .ZN(n176) );
  MOAI22D1BWP30P140LVT U211 ( .A1(n183), .A2(n176), .B1(n274), .B2(
        i_data_bus[208]), .ZN(n177) );
  AOI21D1BWP30P140LVT U212 ( .A1(n1), .A2(i_data_bus[240]), .B(n177), .ZN(n179) );
  ND2D1BWP30P140LVT U213 ( .A1(n288), .A2(i_data_bus[16]), .ZN(n178) );
  ND4D1BWP30P140LVT U214 ( .A1(n181), .A2(n180), .A3(n179), .A4(n178), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U215 ( .A1(n282), .A2(i_data_bus[79]), .B1(n281), .B2(
        i_data_bus[47]), .ZN(n188) );
  AOI22D1BWP30P140LVT U216 ( .A1(n4), .A2(i_data_bus[111]), .B1(n283), .B2(
        i_data_bus[143]), .ZN(n187) );
  INVD1BWP30P140LVT U217 ( .I(i_data_bus[175]), .ZN(n182) );
  MOAI22D1BWP30P140LVT U218 ( .A1(n285), .A2(n182), .B1(n274), .B2(
        i_data_bus[207]), .ZN(n184) );
  AOI21D1BWP30P140LVT U219 ( .A1(n1), .A2(i_data_bus[239]), .B(n184), .ZN(n186) );
  ND2D1BWP30P140LVT U220 ( .A1(n288), .A2(i_data_bus[15]), .ZN(n185) );
  ND4D1BWP30P140LVT U221 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U222 ( .A1(n265), .A2(i_data_bus[76]), .B1(n264), .B2(
        i_data_bus[44]), .ZN(n195) );
  AOI22D1BWP30P140LVT U223 ( .A1(n4), .A2(i_data_bus[108]), .B1(n266), .B2(
        i_data_bus[140]), .ZN(n194) );
  INVD1BWP30P140LVT U224 ( .I(i_data_bus[204]), .ZN(n190) );
  INVD1BWP30P140LVT U225 ( .I(i_data_bus[172]), .ZN(n189) );
  OAI22D1BWP30P140LVT U226 ( .A1(n3), .A2(n190), .B1(n285), .B2(n189), .ZN(
        n191) );
  AOI21D1BWP30P140LVT U227 ( .A1(n1), .A2(i_data_bus[236]), .B(n191), .ZN(n193) );
  ND2D1BWP30P140LVT U228 ( .A1(n269), .A2(i_data_bus[12]), .ZN(n192) );
  ND4D1BWP30P140LVT U229 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .ZN(
        N381) );
  AOI22D1BWP30P140LVT U230 ( .A1(n265), .A2(i_data_bus[75]), .B1(n264), .B2(
        i_data_bus[43]), .ZN(n202) );
  AOI22D1BWP30P140LVT U231 ( .A1(n4), .A2(i_data_bus[107]), .B1(n266), .B2(
        i_data_bus[139]), .ZN(n201) );
  INVD1BWP30P140LVT U232 ( .I(i_data_bus[203]), .ZN(n197) );
  INVD1BWP30P140LVT U233 ( .I(i_data_bus[171]), .ZN(n196) );
  OAI22D1BWP30P140LVT U234 ( .A1(n3), .A2(n197), .B1(n285), .B2(n196), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U235 ( .A1(n1), .A2(i_data_bus[235]), .B(n198), .ZN(n200) );
  ND2D1BWP30P140LVT U236 ( .A1(n269), .A2(i_data_bus[11]), .ZN(n199) );
  ND4D1BWP30P140LVT U237 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(
        N380) );
  AOI22D1BWP30P140LVT U238 ( .A1(n265), .A2(i_data_bus[74]), .B1(n264), .B2(
        i_data_bus[42]), .ZN(n209) );
  AOI22D1BWP30P140LVT U239 ( .A1(n4), .A2(i_data_bus[106]), .B1(n266), .B2(
        i_data_bus[138]), .ZN(n208) );
  INVD1BWP30P140LVT U240 ( .I(i_data_bus[202]), .ZN(n204) );
  INVD1BWP30P140LVT U241 ( .I(i_data_bus[170]), .ZN(n203) );
  OAI22D1BWP30P140LVT U242 ( .A1(n3), .A2(n204), .B1(n285), .B2(n203), .ZN(
        n205) );
  AOI21D1BWP30P140LVT U243 ( .A1(n1), .A2(i_data_bus[234]), .B(n205), .ZN(n207) );
  ND2D1BWP30P140LVT U244 ( .A1(n269), .A2(i_data_bus[10]), .ZN(n206) );
  ND4D1BWP30P140LVT U245 ( .A1(n209), .A2(n208), .A3(n207), .A4(n206), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U246 ( .A1(n265), .A2(i_data_bus[73]), .B1(n264), .B2(
        i_data_bus[41]), .ZN(n216) );
  AOI22D1BWP30P140LVT U247 ( .A1(n4), .A2(i_data_bus[105]), .B1(n266), .B2(
        i_data_bus[137]), .ZN(n215) );
  INVD1BWP30P140LVT U248 ( .I(i_data_bus[201]), .ZN(n211) );
  INVD1BWP30P140LVT U249 ( .I(i_data_bus[169]), .ZN(n210) );
  OAI22D1BWP30P140LVT U250 ( .A1(n3), .A2(n211), .B1(n285), .B2(n210), .ZN(
        n212) );
  AOI21D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[233]), .B(n212), .ZN(n214) );
  ND2D1BWP30P140LVT U252 ( .A1(n269), .A2(i_data_bus[9]), .ZN(n213) );
  ND4D1BWP30P140LVT U253 ( .A1(n216), .A2(n215), .A3(n214), .A4(n213), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U254 ( .A1(n265), .A2(i_data_bus[71]), .B1(n264), .B2(
        i_data_bus[39]), .ZN(n223) );
  AOI22D1BWP30P140LVT U255 ( .A1(n4), .A2(i_data_bus[103]), .B1(n266), .B2(
        i_data_bus[135]), .ZN(n222) );
  INVD1BWP30P140LVT U256 ( .I(i_data_bus[199]), .ZN(n218) );
  INVD1BWP30P140LVT U257 ( .I(i_data_bus[167]), .ZN(n217) );
  OAI22D1BWP30P140LVT U258 ( .A1(n3), .A2(n218), .B1(n285), .B2(n217), .ZN(
        n219) );
  AOI21D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[231]), .B(n219), .ZN(n221) );
  ND2D1BWP30P140LVT U260 ( .A1(n269), .A2(i_data_bus[7]), .ZN(n220) );
  ND4D1BWP30P140LVT U261 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U262 ( .A1(n265), .A2(i_data_bus[70]), .B1(n264), .B2(
        i_data_bus[38]), .ZN(n230) );
  AOI22D1BWP30P140LVT U263 ( .A1(n4), .A2(i_data_bus[102]), .B1(n266), .B2(
        i_data_bus[134]), .ZN(n229) );
  INVD1BWP30P140LVT U264 ( .I(i_data_bus[198]), .ZN(n225) );
  INVD1BWP30P140LVT U265 ( .I(i_data_bus[166]), .ZN(n224) );
  OAI22D1BWP30P140LVT U266 ( .A1(n3), .A2(n225), .B1(n285), .B2(n224), .ZN(
        n226) );
  AOI21D1BWP30P140LVT U267 ( .A1(n1), .A2(i_data_bus[230]), .B(n226), .ZN(n228) );
  ND2D1BWP30P140LVT U268 ( .A1(n269), .A2(i_data_bus[6]), .ZN(n227) );
  ND4D1BWP30P140LVT U269 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U270 ( .A1(n265), .A2(i_data_bus[69]), .B1(n264), .B2(
        i_data_bus[37]), .ZN(n237) );
  AOI22D1BWP30P140LVT U271 ( .A1(n4), .A2(i_data_bus[101]), .B1(n266), .B2(
        i_data_bus[133]), .ZN(n236) );
  INVD1BWP30P140LVT U272 ( .I(i_data_bus[197]), .ZN(n232) );
  INVD1BWP30P140LVT U273 ( .I(i_data_bus[165]), .ZN(n231) );
  OAI22D1BWP30P140LVT U274 ( .A1(n3), .A2(n232), .B1(n285), .B2(n231), .ZN(
        n233) );
  AOI21D1BWP30P140LVT U275 ( .A1(n1), .A2(i_data_bus[229]), .B(n233), .ZN(n235) );
  ND2D1BWP30P140LVT U276 ( .A1(n269), .A2(i_data_bus[5]), .ZN(n234) );
  ND4D1BWP30P140LVT U277 ( .A1(n237), .A2(n236), .A3(n235), .A4(n234), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U278 ( .A1(n4), .A2(i_data_bus[104]), .B1(n266), .B2(
        i_data_bus[136]), .ZN(n243) );
  INVD1BWP30P140LVT U279 ( .I(i_data_bus[168]), .ZN(n239) );
  INVD1BWP30P140LVT U280 ( .I(i_data_bus[200]), .ZN(n238) );
  OAI22D1BWP30P140LVT U281 ( .A1(n285), .A2(n239), .B1(n3), .B2(n238), .ZN(
        n240) );
  AOI21OPTREPBD1BWP30P140LVT U282 ( .A1(n1), .A2(i_data_bus[232]), .B(n240), 
        .ZN(n242) );
  ND2D1BWP30P140LVT U283 ( .A1(n269), .A2(i_data_bus[8]), .ZN(n241) );
  AOI22D1BWP30P140LVT U284 ( .A1(n265), .A2(i_data_bus[68]), .B1(n264), .B2(
        i_data_bus[36]), .ZN(n251) );
  AOI22D1BWP30P140LVT U285 ( .A1(n4), .A2(i_data_bus[100]), .B1(n266), .B2(
        i_data_bus[132]), .ZN(n250) );
  INVD1BWP30P140LVT U286 ( .I(i_data_bus[196]), .ZN(n246) );
  INVD1BWP30P140LVT U287 ( .I(i_data_bus[164]), .ZN(n245) );
  OAI22D1BWP30P140LVT U288 ( .A1(n3), .A2(n246), .B1(n285), .B2(n245), .ZN(
        n247) );
  AOI21D1BWP30P140LVT U289 ( .A1(n1), .A2(i_data_bus[228]), .B(n247), .ZN(n249) );
  ND2D1BWP30P140LVT U290 ( .A1(n269), .A2(i_data_bus[4]), .ZN(n248) );
  ND4D1BWP30P140LVT U291 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U292 ( .A1(n265), .A2(i_data_bus[67]), .B1(n264), .B2(
        i_data_bus[35]), .ZN(n257) );
  AOI22D1BWP30P140LVT U293 ( .A1(n4), .A2(i_data_bus[99]), .B1(n266), .B2(
        i_data_bus[131]), .ZN(n256) );
  INVD1BWP30P140LVT U294 ( .I(i_data_bus[163]), .ZN(n252) );
  MOAI22D1BWP30P140LVT U295 ( .A1(n285), .A2(n252), .B1(n274), .B2(
        i_data_bus[195]), .ZN(n253) );
  AOI21D1BWP30P140LVT U296 ( .A1(n1), .A2(i_data_bus[227]), .B(n253), .ZN(n255) );
  ND2D1BWP30P140LVT U297 ( .A1(n269), .A2(i_data_bus[3]), .ZN(n254) );
  ND4D1BWP30P140LVT U298 ( .A1(n257), .A2(n256), .A3(n255), .A4(n254), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U299 ( .A1(n265), .A2(i_data_bus[66]), .B1(n264), .B2(
        i_data_bus[34]), .ZN(n263) );
  AOI22D1BWP30P140LVT U300 ( .A1(n4), .A2(i_data_bus[98]), .B1(n266), .B2(
        i_data_bus[130]), .ZN(n262) );
  INVD1BWP30P140LVT U301 ( .I(i_data_bus[162]), .ZN(n258) );
  MOAI22D1BWP30P140LVT U302 ( .A1(n285), .A2(n258), .B1(n274), .B2(
        i_data_bus[194]), .ZN(n259) );
  AOI21D1BWP30P140LVT U303 ( .A1(n1), .A2(i_data_bus[226]), .B(n259), .ZN(n261) );
  ND2D1BWP30P140LVT U304 ( .A1(n269), .A2(i_data_bus[2]), .ZN(n260) );
  ND4D1BWP30P140LVT U305 ( .A1(n263), .A2(n262), .A3(n261), .A4(n260), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U306 ( .A1(n265), .A2(i_data_bus[65]), .B1(n264), .B2(
        i_data_bus[33]), .ZN(n273) );
  AOI22D1BWP30P140LVT U307 ( .A1(n4), .A2(i_data_bus[97]), .B1(n266), .B2(
        i_data_bus[129]), .ZN(n272) );
  INVD1BWP30P140LVT U308 ( .I(i_data_bus[161]), .ZN(n267) );
  MOAI22D1BWP30P140LVT U309 ( .A1(n285), .A2(n267), .B1(n274), .B2(
        i_data_bus[193]), .ZN(n268) );
  AOI21D1BWP30P140LVT U310 ( .A1(n1), .A2(i_data_bus[225]), .B(n268), .ZN(n271) );
  ND2D1BWP30P140LVT U311 ( .A1(n269), .A2(i_data_bus[1]), .ZN(n270) );
  ND4D1BWP30P140LVT U312 ( .A1(n273), .A2(n272), .A3(n271), .A4(n270), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U313 ( .A1(n282), .A2(i_data_bus[78]), .B1(n281), .B2(
        i_data_bus[46]), .ZN(n280) );
  AOI22D1BWP30P140LVT U314 ( .A1(n4), .A2(i_data_bus[110]), .B1(n283), .B2(
        i_data_bus[142]), .ZN(n279) );
  INVD1BWP30P140LVT U315 ( .I(i_data_bus[174]), .ZN(n275) );
  MOAI22D1BWP30P140LVT U316 ( .A1(n285), .A2(n275), .B1(n274), .B2(
        i_data_bus[206]), .ZN(n276) );
  AOI21D1BWP30P140LVT U317 ( .A1(n1), .A2(i_data_bus[238]), .B(n276), .ZN(n278) );
  ND2D1BWP30P140LVT U318 ( .A1(n288), .A2(i_data_bus[14]), .ZN(n277) );
  ND4D1BWP30P140LVT U319 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U320 ( .A1(n282), .A2(i_data_bus[77]), .B1(n281), .B2(
        i_data_bus[45]), .ZN(n292) );
  AOI22D1BWP30P140LVT U321 ( .A1(n4), .A2(i_data_bus[109]), .B1(n283), .B2(
        i_data_bus[141]), .ZN(n291) );
  INVD1BWP30P140LVT U322 ( .I(i_data_bus[205]), .ZN(n286) );
  INVD1BWP30P140LVT U323 ( .I(i_data_bus[173]), .ZN(n284) );
  OAI22D1BWP30P140LVT U324 ( .A1(n3), .A2(n286), .B1(n285), .B2(n284), .ZN(
        n287) );
  AOI21D1BWP30P140LVT U325 ( .A1(n1), .A2(i_data_bus[237]), .B(n287), .ZN(n290) );
  ND2D1BWP30P140LVT U326 ( .A1(n288), .A2(i_data_bus[13]), .ZN(n289) );
  ND4D1BWP30P140LVT U327 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_6 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  AOI21D1BWP30P140LVT U3 ( .A1(n73), .A2(i_data_bus[238]), .B(n274), .ZN(n277)
         );
  INVD3BWP30P140LVT U4 ( .I(n46), .ZN(n1) );
  INR2D1BWP30P140LVT U5 ( .A1(n5), .B1(n18), .ZN(n31) );
  OR2D1BWP30P140LVT U6 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n18) );
  AOI21D1BWP30P140LVT U7 ( .A1(n73), .A2(i_data_bus[237]), .B(n286), .ZN(n290)
         );
  INVD4BWP30P140LVT U8 ( .I(n131), .ZN(n2) );
  INVD1BWP30P140LVT U9 ( .I(n130), .ZN(n3) );
  INVD4BWP30P140LVT U10 ( .I(n134), .ZN(n283) );
  INR2D4BWP30P140LVT U11 ( .A1(n43), .B1(n42), .ZN(n130) );
  NR2D1BWP30P140LVT U12 ( .A1(n41), .A2(n40), .ZN(n43) );
  ND2D1BWP30P140LVT U13 ( .A1(n12), .A2(n11), .ZN(n22) );
  INVD1BWP30P140LVT U14 ( .I(n24), .ZN(n78) );
  INVD1BWP30P140LVT U15 ( .I(n78), .ZN(n275) );
  INVD1BWP30P140LVT U16 ( .I(n78), .ZN(n287) );
  ND2D1BWP30P140LVT U17 ( .A1(n14), .A2(n13), .ZN(n15) );
  AOI21D1BWP30P140LVT U18 ( .A1(n73), .A2(i_data_bus[225]), .B(n229), .ZN(n231) );
  AOI21D1BWP30P140LVT U19 ( .A1(n287), .A2(i_data_bus[239]), .B(n258), .ZN(
        n260) );
  INVD1BWP30P140LVT U20 ( .I(n9), .ZN(n138) );
  INVD1BWP30P140LVT U21 ( .I(n33), .ZN(n131) );
  INR2D1BWP30P140LVT U22 ( .A1(n39), .B1(n42), .ZN(n129) );
  CKBD1BWP30P140LVT U23 ( .I(n133), .Z(n55) );
  INVD1BWP30P140LVT U24 ( .I(i_cmd[0]), .ZN(n28) );
  INR3D0BWP30P140LVT U25 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n28), .ZN(n8)
         );
  INVD1BWP30P140LVT U26 ( .I(rst), .ZN(n4) );
  ND2D1BWP30P140LVT U27 ( .A1(n4), .A2(i_en), .ZN(n10) );
  NR2D1BWP30P140LVT U28 ( .A1(i_cmd[5]), .A2(n10), .ZN(n5) );
  INVD1BWP30P140LVT U29 ( .I(i_cmd[3]), .ZN(n6) );
  INVD1BWP30P140LVT U30 ( .I(i_cmd[2]), .ZN(n38) );
  ND2OPTIBD1BWP30P140LVT U31 ( .A1(n6), .A2(n38), .ZN(n41) );
  NR2D1BWP30P140LVT U32 ( .A1(n41), .A2(i_cmd[1]), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U33 ( .A1(n31), .A2(n7), .ZN(n35) );
  INR2D1BWP30P140LVT U34 ( .A1(n8), .B1(n35), .ZN(n9) );
  NR4D1BWP30P140LVT U35 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .A3(i_cmd[1]), .A4(n10), .ZN(n12) );
  NR2D1BWP30P140LVT U36 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n11) );
  NR2D1BWP30P140LVT U37 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n14) );
  CKAN2D1BWP30P140LVT U38 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n13) );
  OR2D2BWP30P140LVT U39 ( .A1(n22), .A2(n15), .Z(n285) );
  INVD1BWP30P140LVT U40 ( .I(n285), .ZN(n25) );
  INVD1BWP30P140LVT U41 ( .I(i_valid[5]), .ZN(n16) );
  IND2D1BWP30P140LVT U42 ( .A1(n16), .B1(i_cmd[5]), .ZN(n17) );
  NR2D1BWP30P140LVT U43 ( .A1(n18), .A2(n17), .ZN(n19) );
  INR2D1BWP30P140LVT U44 ( .A1(n19), .B1(n22), .ZN(n20) );
  INVD2BWP30P140LVT U45 ( .I(n20), .ZN(n133) );
  INVD1BWP30P140LVT U46 ( .I(i_cmd[7]), .ZN(n21) );
  INR4D0BWP30P140LVT U47 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n21), .ZN(n23) );
  INR2D1BWP30P140LVT U48 ( .A1(n23), .B1(n22), .ZN(n24) );
  NR4D0BWP30P140LVT U49 ( .A1(n267), .A2(n25), .A3(n134), .A4(n287), .ZN(n45)
         );
  OR2D1BWP30P140LVT U50 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n27) );
  ND2D1BWP30P140LVT U51 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n26) );
  NR2D1BWP30P140LVT U52 ( .A1(n27), .A2(n26), .ZN(n32) );
  INVD1BWP30P140LVT U53 ( .I(i_cmd[4]), .ZN(n29) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n29), .A2(n28), .Z(n30) );
  ND2OPTIBD2BWP30P140LVT U55 ( .A1(n31), .A2(n30), .ZN(n42) );
  INR2D1BWP30P140LVT U56 ( .A1(n32), .B1(n42), .ZN(n33) );
  ND2OPTIBD1BWP30P140LVT U57 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n34) );
  NR2D1BWP30P140LVT U58 ( .A1(n34), .A2(i_cmd[0]), .ZN(n36) );
  INR2D1BWP30P140LVT U59 ( .A1(n36), .B1(n35), .ZN(n37) );
  INVD1BWP30P140LVT U60 ( .I(n37), .ZN(n132) );
  INVD3BWP30P140LVT U61 ( .I(n132), .ZN(n281) );
  NR2D1BWP30P140LVT U62 ( .A1(n33), .A2(n281), .ZN(n44) );
  INR4D0BWP30P140LVT U63 ( .A1(i_valid[2]), .B1(i_cmd[1]), .B2(i_cmd[3]), .B3(
        n38), .ZN(n39) );
  INVD1BWP30P140LVT U64 ( .I(n129), .ZN(n46) );
  ND2D1BWP30P140LVT U65 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n40) );
  ND4D1BWP30P140LVT U66 ( .A1(n45), .A2(n44), .A3(n46), .A4(n3), .ZN(N402) );
  AOI22D1BWP30P140LVT U67 ( .A1(n1), .A2(i_data_bus[94]), .B1(n130), .B2(
        i_data_bus[62]), .ZN(n53) );
  AOI22D1BWP30P140LVT U68 ( .A1(n2), .A2(i_data_bus[126]), .B1(n281), .B2(
        i_data_bus[158]), .ZN(n52) );
  INVD1BWP30P140LVT U69 ( .I(n78), .ZN(n73) );
  INVD1BWP30P140LVT U70 ( .I(i_data_bus[222]), .ZN(n48) );
  INVD1BWP30P140LVT U71 ( .I(i_data_bus[190]), .ZN(n47) );
  OAI22D1BWP30P140LVT U72 ( .A1(n285), .A2(n48), .B1(n55), .B2(n47), .ZN(n49)
         );
  AOI21D1BWP30P140LVT U73 ( .A1(n287), .A2(i_data_bus[254]), .B(n49), .ZN(n51)
         );
  ND2D1BWP30P140LVT U74 ( .A1(n288), .A2(i_data_bus[30]), .ZN(n50) );
  ND4D1BWP30P140LVT U75 ( .A1(n53), .A2(n52), .A3(n51), .A4(n50), .ZN(N399) );
  AOI22D1BWP30P140LVT U76 ( .A1(n1), .A2(i_data_bus[95]), .B1(n130), .B2(
        i_data_bus[63]), .ZN(n61) );
  AOI22D1BWP30P140LVT U77 ( .A1(n2), .A2(i_data_bus[127]), .B1(n281), .B2(
        i_data_bus[159]), .ZN(n60) );
  INVD1BWP30P140LVT U78 ( .I(i_data_bus[223]), .ZN(n56) );
  INVD1BWP30P140LVT U79 ( .I(i_data_bus[191]), .ZN(n54) );
  OAI22D1BWP30P140LVT U80 ( .A1(n285), .A2(n56), .B1(n55), .B2(n54), .ZN(n57)
         );
  AOI21D1BWP30P140LVT U81 ( .A1(n287), .A2(i_data_bus[255]), .B(n57), .ZN(n59)
         );
  ND2D1BWP30P140LVT U82 ( .A1(n267), .A2(i_data_bus[31]), .ZN(n58) );
  ND4D1BWP30P140LVT U83 ( .A1(n61), .A2(n60), .A3(n59), .A4(n58), .ZN(N400) );
  AOI22D1BWP30P140LVT U84 ( .A1(n1), .A2(i_data_bus[93]), .B1(n130), .B2(
        i_data_bus[61]), .ZN(n69) );
  AOI22D1BWP30P140LVT U85 ( .A1(n2), .A2(i_data_bus[125]), .B1(n281), .B2(
        i_data_bus[157]), .ZN(n68) );
  INVD1BWP30P140LVT U86 ( .I(i_data_bus[221]), .ZN(n64) );
  INVD2BWP30P140LVT U87 ( .I(n133), .ZN(n62) );
  INVD3BWP30P140LVT U88 ( .I(n62), .ZN(n256) );
  INVD1BWP30P140LVT U89 ( .I(i_data_bus[189]), .ZN(n63) );
  OAI22D1BWP30P140LVT U90 ( .A1(n285), .A2(n64), .B1(n256), .B2(n63), .ZN(n65)
         );
  AOI21D1BWP30P140LVT U91 ( .A1(n275), .A2(i_data_bus[253]), .B(n65), .ZN(n67)
         );
  ND2D1BWP30P140LVT U92 ( .A1(n288), .A2(i_data_bus[29]), .ZN(n66) );
  ND4D1BWP30P140LVT U93 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(N398) );
  AOI22D1BWP30P140LVT U94 ( .A1(n1), .A2(i_data_bus[92]), .B1(n130), .B2(
        i_data_bus[60]), .ZN(n77) );
  AOI22D1BWP30P140LVT U95 ( .A1(n2), .A2(i_data_bus[124]), .B1(n281), .B2(
        i_data_bus[156]), .ZN(n76) );
  INVD1BWP30P140LVT U96 ( .I(i_data_bus[220]), .ZN(n71) );
  INVD1BWP30P140LVT U97 ( .I(i_data_bus[188]), .ZN(n70) );
  OAI22D1BWP30P140LVT U98 ( .A1(n285), .A2(n71), .B1(n256), .B2(n70), .ZN(n72)
         );
  AOI21D1BWP30P140LVT U99 ( .A1(n73), .A2(i_data_bus[252]), .B(n72), .ZN(n75)
         );
  ND2D1BWP30P140LVT U100 ( .A1(n267), .A2(i_data_bus[28]), .ZN(n74) );
  ND4D1BWP30P140LVT U101 ( .A1(n77), .A2(n76), .A3(n75), .A4(n74), .ZN(N397)
         );
  AOI22D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[91]), .B1(n130), .B2(
        i_data_bus[59]), .ZN(n85) );
  AOI22D1BWP30P140LVT U103 ( .A1(n2), .A2(i_data_bus[123]), .B1(n281), .B2(
        i_data_bus[155]), .ZN(n84) );
  INVD1BWP30P140LVT U104 ( .I(i_data_bus[219]), .ZN(n80) );
  INVD1BWP30P140LVT U105 ( .I(i_data_bus[187]), .ZN(n79) );
  OAI22D1BWP30P140LVT U106 ( .A1(n285), .A2(n80), .B1(n256), .B2(n79), .ZN(n81) );
  AOI21D1BWP30P140LVT U107 ( .A1(n275), .A2(i_data_bus[251]), .B(n81), .ZN(n83) );
  ND2D1BWP30P140LVT U108 ( .A1(n288), .A2(i_data_bus[27]), .ZN(n82) );
  ND4D1BWP30P140LVT U109 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(N396)
         );
  AOI22D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[90]), .B1(n130), .B2(
        i_data_bus[58]), .ZN(n92) );
  AOI22D1BWP30P140LVT U111 ( .A1(n2), .A2(i_data_bus[122]), .B1(n281), .B2(
        i_data_bus[154]), .ZN(n91) );
  INVD1BWP30P140LVT U112 ( .I(i_data_bus[218]), .ZN(n87) );
  INVD1BWP30P140LVT U113 ( .I(i_data_bus[186]), .ZN(n86) );
  OAI22D1BWP30P140LVT U114 ( .A1(n285), .A2(n87), .B1(n256), .B2(n86), .ZN(n88) );
  AOI21D1BWP30P140LVT U115 ( .A1(n73), .A2(i_data_bus[250]), .B(n88), .ZN(n90)
         );
  ND2D1BWP30P140LVT U116 ( .A1(n9), .A2(i_data_bus[26]), .ZN(n89) );
  ND4D1BWP30P140LVT U117 ( .A1(n92), .A2(n91), .A3(n90), .A4(n89), .ZN(N395)
         );
  INVD1BWP30P140LVT U118 ( .I(n130), .ZN(n93) );
  INVD2BWP30P140LVT U119 ( .I(n93), .ZN(n280) );
  AOI22D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[89]), .B1(n280), .B2(
        i_data_bus[57]), .ZN(n100) );
  AOI22D1BWP30P140LVT U121 ( .A1(n2), .A2(i_data_bus[121]), .B1(n281), .B2(
        i_data_bus[153]), .ZN(n99) );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[217]), .ZN(n95) );
  INVD1BWP30P140LVT U123 ( .I(i_data_bus[185]), .ZN(n94) );
  OAI22D1BWP30P140LVT U124 ( .A1(n285), .A2(n95), .B1(n256), .B2(n94), .ZN(n96) );
  AOI21D1BWP30P140LVT U125 ( .A1(n287), .A2(i_data_bus[249]), .B(n96), .ZN(n98) );
  INVD2BWP30P140LVT U126 ( .I(n138), .ZN(n288) );
  ND2D1BWP30P140LVT U127 ( .A1(n288), .A2(i_data_bus[25]), .ZN(n97) );
  ND4D1BWP30P140LVT U128 ( .A1(n100), .A2(n99), .A3(n98), .A4(n97), .ZN(N394)
         );
  AOI22D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[88]), .B1(n280), .B2(
        i_data_bus[56]), .ZN(n107) );
  AOI22D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[120]), .B1(n281), .B2(
        i_data_bus[152]), .ZN(n106) );
  INVD1BWP30P140LVT U131 ( .I(i_data_bus[216]), .ZN(n102) );
  INVD1BWP30P140LVT U132 ( .I(i_data_bus[184]), .ZN(n101) );
  OAI22D1BWP30P140LVT U133 ( .A1(n285), .A2(n102), .B1(n256), .B2(n101), .ZN(
        n103) );
  AOI21D1BWP30P140LVT U134 ( .A1(n275), .A2(i_data_bus[248]), .B(n103), .ZN(
        n105) );
  ND2D1BWP30P140LVT U135 ( .A1(n288), .A2(i_data_bus[24]), .ZN(n104) );
  ND4D1BWP30P140LVT U136 ( .A1(n107), .A2(n106), .A3(n105), .A4(n104), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U137 ( .A1(n1), .A2(i_data_bus[87]), .B1(n280), .B2(
        i_data_bus[55]), .ZN(n114) );
  AOI22D1BWP30P140LVT U138 ( .A1(n2), .A2(i_data_bus[119]), .B1(n281), .B2(
        i_data_bus[151]), .ZN(n113) );
  INVD1BWP30P140LVT U139 ( .I(i_data_bus[215]), .ZN(n109) );
  INVD1BWP30P140LVT U140 ( .I(i_data_bus[183]), .ZN(n108) );
  OAI22D1BWP30P140LVT U141 ( .A1(n285), .A2(n109), .B1(n256), .B2(n108), .ZN(
        n110) );
  AOI21D1BWP30P140LVT U142 ( .A1(n73), .A2(i_data_bus[247]), .B(n110), .ZN(
        n112) );
  ND2D1BWP30P140LVT U143 ( .A1(n288), .A2(i_data_bus[23]), .ZN(n111) );
  ND4D1BWP30P140LVT U144 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U145 ( .A1(n1), .A2(i_data_bus[86]), .B1(n280), .B2(
        i_data_bus[54]), .ZN(n121) );
  AOI22D1BWP30P140LVT U146 ( .A1(n2), .A2(i_data_bus[118]), .B1(n281), .B2(
        i_data_bus[150]), .ZN(n120) );
  INVD1BWP30P140LVT U147 ( .I(i_data_bus[214]), .ZN(n116) );
  INVD1BWP30P140LVT U148 ( .I(i_data_bus[182]), .ZN(n115) );
  OAI22D1BWP30P140LVT U149 ( .A1(n285), .A2(n116), .B1(n256), .B2(n115), .ZN(
        n117) );
  AOI21D1BWP30P140LVT U150 ( .A1(n287), .A2(i_data_bus[246]), .B(n117), .ZN(
        n119) );
  ND2D1BWP30P140LVT U151 ( .A1(n288), .A2(i_data_bus[22]), .ZN(n118) );
  ND4D1BWP30P140LVT U152 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U153 ( .A1(n1), .A2(i_data_bus[85]), .B1(n280), .B2(
        i_data_bus[53]), .ZN(n128) );
  AOI22D1BWP30P140LVT U154 ( .A1(n2), .A2(i_data_bus[117]), .B1(n281), .B2(
        i_data_bus[149]), .ZN(n127) );
  INVD1BWP30P140LVT U155 ( .I(i_data_bus[213]), .ZN(n123) );
  INVD1BWP30P140LVT U156 ( .I(i_data_bus[181]), .ZN(n122) );
  OAI22D1BWP30P140LVT U157 ( .A1(n285), .A2(n123), .B1(n256), .B2(n122), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U158 ( .A1(n275), .A2(i_data_bus[245]), .B(n124), .ZN(
        n126) );
  ND2D1BWP30P140LVT U159 ( .A1(n288), .A2(i_data_bus[21]), .ZN(n125) );
  ND4D1BWP30P140LVT U160 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(
        N390) );
  INVD2BWP30P140LVT U161 ( .I(n3), .ZN(n263) );
  AOI22D1BWP30P140LVT U162 ( .A1(n1), .A2(i_data_bus[72]), .B1(n263), .B2(
        i_data_bus[40]), .ZN(n142) );
  INVD2BWP30P140LVT U163 ( .I(n132), .ZN(n264) );
  AOI22D1BWP30P140LVT U164 ( .A1(n2), .A2(i_data_bus[104]), .B1(n264), .B2(
        i_data_bus[136]), .ZN(n141) );
  INVD1BWP30P140LVT U165 ( .I(i_data_bus[200]), .ZN(n136) );
  INVD2BWP30P140LVT U166 ( .I(n133), .ZN(n134) );
  INVD1BWP30P140LVT U167 ( .I(i_data_bus[168]), .ZN(n135) );
  OAI22D1BWP30P140LVT U168 ( .A1(n285), .A2(n136), .B1(n283), .B2(n135), .ZN(
        n137) );
  AOI21D1BWP30P140LVT U169 ( .A1(n73), .A2(i_data_bus[232]), .B(n137), .ZN(
        n140) );
  INVD2BWP30P140LVT U170 ( .I(n138), .ZN(n267) );
  ND2D1BWP30P140LVT U171 ( .A1(n267), .A2(i_data_bus[8]), .ZN(n139) );
  ND4D1BWP30P140LVT U172 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U173 ( .A1(n1), .A2(i_data_bus[76]), .B1(n263), .B2(
        i_data_bus[44]), .ZN(n149) );
  AOI22D1BWP30P140LVT U174 ( .A1(n2), .A2(i_data_bus[108]), .B1(n264), .B2(
        i_data_bus[140]), .ZN(n148) );
  INVD1BWP30P140LVT U175 ( .I(i_data_bus[204]), .ZN(n144) );
  INVD1BWP30P140LVT U176 ( .I(i_data_bus[172]), .ZN(n143) );
  OAI22D1BWP30P140LVT U177 ( .A1(n285), .A2(n144), .B1(n283), .B2(n143), .ZN(
        n145) );
  AOI21D1BWP30P140LVT U178 ( .A1(n275), .A2(i_data_bus[236]), .B(n145), .ZN(
        n147) );
  ND2D1BWP30P140LVT U179 ( .A1(n267), .A2(i_data_bus[12]), .ZN(n146) );
  ND4D1BWP30P140LVT U180 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(
        N381) );
  AOI22D1BWP30P140LVT U181 ( .A1(n1), .A2(i_data_bus[75]), .B1(n263), .B2(
        i_data_bus[43]), .ZN(n156) );
  AOI22D1BWP30P140LVT U182 ( .A1(n2), .A2(i_data_bus[107]), .B1(n264), .B2(
        i_data_bus[139]), .ZN(n155) );
  INVD1BWP30P140LVT U183 ( .I(i_data_bus[203]), .ZN(n151) );
  INVD1BWP30P140LVT U184 ( .I(i_data_bus[171]), .ZN(n150) );
  OAI22D1BWP30P140LVT U185 ( .A1(n285), .A2(n151), .B1(n283), .B2(n150), .ZN(
        n152) );
  AOI21D1BWP30P140LVT U186 ( .A1(n73), .A2(i_data_bus[235]), .B(n152), .ZN(
        n154) );
  ND2D1BWP30P140LVT U187 ( .A1(n267), .A2(i_data_bus[11]), .ZN(n153) );
  ND4D1BWP30P140LVT U188 ( .A1(n156), .A2(n155), .A3(n154), .A4(n153), .ZN(
        N380) );
  AOI22D1BWP30P140LVT U189 ( .A1(n1), .A2(i_data_bus[74]), .B1(n263), .B2(
        i_data_bus[42]), .ZN(n163) );
  AOI22D1BWP30P140LVT U190 ( .A1(n2), .A2(i_data_bus[106]), .B1(n264), .B2(
        i_data_bus[138]), .ZN(n162) );
  INVD1BWP30P140LVT U191 ( .I(i_data_bus[202]), .ZN(n158) );
  INVD1BWP30P140LVT U192 ( .I(i_data_bus[170]), .ZN(n157) );
  OAI22D1BWP30P140LVT U193 ( .A1(n285), .A2(n158), .B1(n283), .B2(n157), .ZN(
        n159) );
  AOI21D1BWP30P140LVT U194 ( .A1(n287), .A2(i_data_bus[234]), .B(n159), .ZN(
        n161) );
  ND2D1BWP30P140LVT U195 ( .A1(n267), .A2(i_data_bus[10]), .ZN(n160) );
  ND4D1BWP30P140LVT U196 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U197 ( .A1(n1), .A2(i_data_bus[73]), .B1(n263), .B2(
        i_data_bus[41]), .ZN(n170) );
  AOI22D1BWP30P140LVT U198 ( .A1(n2), .A2(i_data_bus[105]), .B1(n264), .B2(
        i_data_bus[137]), .ZN(n169) );
  INVD1BWP30P140LVT U199 ( .I(i_data_bus[201]), .ZN(n165) );
  INVD1BWP30P140LVT U200 ( .I(i_data_bus[169]), .ZN(n164) );
  OAI22D1BWP30P140LVT U201 ( .A1(n285), .A2(n165), .B1(n283), .B2(n164), .ZN(
        n166) );
  AOI21D1BWP30P140LVT U202 ( .A1(n275), .A2(i_data_bus[233]), .B(n166), .ZN(
        n168) );
  ND2D1BWP30P140LVT U203 ( .A1(n267), .A2(i_data_bus[9]), .ZN(n167) );
  ND4D1BWP30P140LVT U204 ( .A1(n170), .A2(n169), .A3(n168), .A4(n167), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U205 ( .A1(n1), .A2(i_data_bus[71]), .B1(n263), .B2(
        i_data_bus[39]), .ZN(n177) );
  AOI22D1BWP30P140LVT U206 ( .A1(n2), .A2(i_data_bus[103]), .B1(n264), .B2(
        i_data_bus[135]), .ZN(n176) );
  INVD1BWP30P140LVT U207 ( .I(i_data_bus[199]), .ZN(n172) );
  INVD1BWP30P140LVT U208 ( .I(i_data_bus[167]), .ZN(n171) );
  OAI22D1BWP30P140LVT U209 ( .A1(n285), .A2(n172), .B1(n283), .B2(n171), .ZN(
        n173) );
  AOI21D1BWP30P140LVT U210 ( .A1(n73), .A2(i_data_bus[231]), .B(n173), .ZN(
        n175) );
  ND2D1BWP30P140LVT U211 ( .A1(n267), .A2(i_data_bus[7]), .ZN(n174) );
  ND4D1BWP30P140LVT U212 ( .A1(n177), .A2(n176), .A3(n175), .A4(n174), .ZN(
        N376) );
  AOI22D1BWP30P140LVT U213 ( .A1(n1), .A2(i_data_bus[70]), .B1(n263), .B2(
        i_data_bus[38]), .ZN(n184) );
  AOI22D1BWP30P140LVT U214 ( .A1(n2), .A2(i_data_bus[102]), .B1(n264), .B2(
        i_data_bus[134]), .ZN(n183) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[198]), .ZN(n179) );
  INVD1BWP30P140LVT U216 ( .I(i_data_bus[166]), .ZN(n178) );
  OAI22D1BWP30P140LVT U217 ( .A1(n285), .A2(n179), .B1(n283), .B2(n178), .ZN(
        n180) );
  AOI21D1BWP30P140LVT U218 ( .A1(n287), .A2(i_data_bus[230]), .B(n180), .ZN(
        n182) );
  ND2D1BWP30P140LVT U219 ( .A1(n267), .A2(i_data_bus[6]), .ZN(n181) );
  ND4D1BWP30P140LVT U220 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U221 ( .A1(n1), .A2(i_data_bus[69]), .B1(n263), .B2(
        i_data_bus[37]), .ZN(n191) );
  AOI22D1BWP30P140LVT U222 ( .A1(n2), .A2(i_data_bus[101]), .B1(n264), .B2(
        i_data_bus[133]), .ZN(n190) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[197]), .ZN(n186) );
  INVD1BWP30P140LVT U224 ( .I(i_data_bus[165]), .ZN(n185) );
  OAI22D1BWP30P140LVT U225 ( .A1(n285), .A2(n186), .B1(n283), .B2(n185), .ZN(
        n187) );
  AOI21D1BWP30P140LVT U226 ( .A1(n275), .A2(i_data_bus[229]), .B(n187), .ZN(
        n189) );
  ND2D1BWP30P140LVT U227 ( .A1(n267), .A2(i_data_bus[5]), .ZN(n188) );
  ND4D1BWP30P140LVT U228 ( .A1(n191), .A2(n190), .A3(n189), .A4(n188), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U229 ( .A1(n1), .A2(i_data_bus[84]), .B1(n280), .B2(
        i_data_bus[52]), .ZN(n198) );
  AOI22D1BWP30P140LVT U230 ( .A1(n2), .A2(i_data_bus[116]), .B1(n281), .B2(
        i_data_bus[148]), .ZN(n197) );
  INVD1BWP30P140LVT U231 ( .I(i_data_bus[212]), .ZN(n193) );
  INVD1BWP30P140LVT U232 ( .I(i_data_bus[180]), .ZN(n192) );
  OAI22D1BWP30P140LVT U233 ( .A1(n285), .A2(n193), .B1(n256), .B2(n192), .ZN(
        n194) );
  AOI21D1BWP30P140LVT U234 ( .A1(n287), .A2(i_data_bus[244]), .B(n194), .ZN(
        n196) );
  ND2D1BWP30P140LVT U235 ( .A1(n288), .A2(i_data_bus[20]), .ZN(n195) );
  ND4D1BWP30P140LVT U236 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U237 ( .A1(n1), .A2(i_data_bus[83]), .B1(n280), .B2(
        i_data_bus[51]), .ZN(n205) );
  AOI22D1BWP30P140LVT U238 ( .A1(n2), .A2(i_data_bus[115]), .B1(n281), .B2(
        i_data_bus[147]), .ZN(n204) );
  INVD1BWP30P140LVT U239 ( .I(i_data_bus[211]), .ZN(n200) );
  INVD1BWP30P140LVT U240 ( .I(i_data_bus[179]), .ZN(n199) );
  OAI22D1BWP30P140LVT U241 ( .A1(n285), .A2(n200), .B1(n256), .B2(n199), .ZN(
        n201) );
  AOI21D1BWP30P140LVT U242 ( .A1(n275), .A2(i_data_bus[243]), .B(n201), .ZN(
        n203) );
  ND2D1BWP30P140LVT U243 ( .A1(n288), .A2(i_data_bus[19]), .ZN(n202) );
  ND4D1BWP30P140LVT U244 ( .A1(n205), .A2(n204), .A3(n203), .A4(n202), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U245 ( .A1(n1), .A2(i_data_bus[68]), .B1(n263), .B2(
        i_data_bus[36]), .ZN(n212) );
  AOI22D1BWP30P140LVT U246 ( .A1(n2), .A2(i_data_bus[100]), .B1(n264), .B2(
        i_data_bus[132]), .ZN(n211) );
  INVD1BWP30P140LVT U247 ( .I(i_data_bus[196]), .ZN(n207) );
  INVD1BWP30P140LVT U248 ( .I(i_data_bus[164]), .ZN(n206) );
  OAI22D1BWP30P140LVT U249 ( .A1(n285), .A2(n207), .B1(n283), .B2(n206), .ZN(
        n208) );
  AOI21D1BWP30P140LVT U250 ( .A1(n73), .A2(i_data_bus[228]), .B(n208), .ZN(
        n210) );
  ND2D1BWP30P140LVT U251 ( .A1(n267), .A2(i_data_bus[4]), .ZN(n209) );
  ND4D1BWP30P140LVT U252 ( .A1(n212), .A2(n211), .A3(n210), .A4(n209), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[67]), .B1(n263), .B2(
        i_data_bus[35]), .ZN(n219) );
  AOI22D1BWP30P140LVT U254 ( .A1(n2), .A2(i_data_bus[99]), .B1(n264), .B2(
        i_data_bus[131]), .ZN(n218) );
  INVD1BWP30P140LVT U255 ( .I(i_data_bus[195]), .ZN(n214) );
  INVD1BWP30P140LVT U256 ( .I(i_data_bus[163]), .ZN(n213) );
  OAI22D1BWP30P140LVT U257 ( .A1(n285), .A2(n214), .B1(n283), .B2(n213), .ZN(
        n215) );
  AOI21D1BWP30P140LVT U258 ( .A1(n287), .A2(i_data_bus[227]), .B(n215), .ZN(
        n217) );
  ND2D1BWP30P140LVT U259 ( .A1(n267), .A2(i_data_bus[3]), .ZN(n216) );
  ND4D1BWP30P140LVT U260 ( .A1(n219), .A2(n218), .A3(n217), .A4(n216), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[66]), .B1(n263), .B2(
        i_data_bus[34]), .ZN(n226) );
  AOI22D1BWP30P140LVT U262 ( .A1(n2), .A2(i_data_bus[98]), .B1(n264), .B2(
        i_data_bus[130]), .ZN(n225) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[194]), .ZN(n221) );
  INVD1BWP30P140LVT U264 ( .I(i_data_bus[162]), .ZN(n220) );
  OAI22D1BWP30P140LVT U265 ( .A1(n285), .A2(n221), .B1(n283), .B2(n220), .ZN(
        n222) );
  AOI21D1BWP30P140LVT U266 ( .A1(n275), .A2(i_data_bus[226]), .B(n222), .ZN(
        n224) );
  ND2D1BWP30P140LVT U267 ( .A1(n267), .A2(i_data_bus[2]), .ZN(n223) );
  ND4D1BWP30P140LVT U268 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U269 ( .A1(n1), .A2(i_data_bus[65]), .B1(n263), .B2(
        i_data_bus[33]), .ZN(n233) );
  AOI22D1BWP30P140LVT U270 ( .A1(n2), .A2(i_data_bus[97]), .B1(n264), .B2(
        i_data_bus[129]), .ZN(n232) );
  INVD1BWP30P140LVT U271 ( .I(i_data_bus[193]), .ZN(n228) );
  INVD1BWP30P140LVT U272 ( .I(i_data_bus[161]), .ZN(n227) );
  OAI22D1BWP30P140LVT U273 ( .A1(n285), .A2(n228), .B1(n283), .B2(n227), .ZN(
        n229) );
  ND2D1BWP30P140LVT U274 ( .A1(n267), .A2(i_data_bus[1]), .ZN(n230) );
  ND4D1BWP30P140LVT U275 ( .A1(n233), .A2(n232), .A3(n231), .A4(n230), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U276 ( .A1(n1), .A2(i_data_bus[82]), .B1(n280), .B2(
        i_data_bus[50]), .ZN(n240) );
  AOI22D1BWP30P140LVT U277 ( .A1(n2), .A2(i_data_bus[114]), .B1(n281), .B2(
        i_data_bus[146]), .ZN(n239) );
  INVD1BWP30P140LVT U278 ( .I(i_data_bus[210]), .ZN(n235) );
  INVD1BWP30P140LVT U279 ( .I(i_data_bus[178]), .ZN(n234) );
  OAI22D1BWP30P140LVT U280 ( .A1(n285), .A2(n235), .B1(n256), .B2(n234), .ZN(
        n236) );
  AOI21D1BWP30P140LVT U281 ( .A1(n73), .A2(i_data_bus[242]), .B(n236), .ZN(
        n238) );
  ND2D1BWP30P140LVT U282 ( .A1(n288), .A2(i_data_bus[18]), .ZN(n237) );
  ND4D1BWP30P140LVT U283 ( .A1(n240), .A2(n239), .A3(n238), .A4(n237), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U284 ( .A1(n1), .A2(i_data_bus[81]), .B1(n280), .B2(
        i_data_bus[49]), .ZN(n247) );
  AOI22D1BWP30P140LVT U285 ( .A1(n2), .A2(i_data_bus[113]), .B1(n281), .B2(
        i_data_bus[145]), .ZN(n246) );
  INVD1BWP30P140LVT U286 ( .I(i_data_bus[209]), .ZN(n242) );
  INVD1BWP30P140LVT U287 ( .I(i_data_bus[177]), .ZN(n241) );
  OAI22D1BWP30P140LVT U288 ( .A1(n285), .A2(n242), .B1(n256), .B2(n241), .ZN(
        n243) );
  AOI21D1BWP30P140LVT U289 ( .A1(n287), .A2(i_data_bus[241]), .B(n243), .ZN(
        n245) );
  ND2D1BWP30P140LVT U290 ( .A1(n288), .A2(i_data_bus[17]), .ZN(n244) );
  ND4D1BWP30P140LVT U291 ( .A1(n247), .A2(n246), .A3(n245), .A4(n244), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U292 ( .A1(n1), .A2(i_data_bus[80]), .B1(n280), .B2(
        i_data_bus[48]), .ZN(n254) );
  AOI22D1BWP30P140LVT U293 ( .A1(n2), .A2(i_data_bus[112]), .B1(n281), .B2(
        i_data_bus[144]), .ZN(n253) );
  INVD1BWP30P140LVT U294 ( .I(i_data_bus[208]), .ZN(n249) );
  INVD1BWP30P140LVT U295 ( .I(i_data_bus[176]), .ZN(n248) );
  OAI22D1BWP30P140LVT U296 ( .A1(n285), .A2(n249), .B1(n256), .B2(n248), .ZN(
        n250) );
  AOI21D1BWP30P140LVT U297 ( .A1(n275), .A2(i_data_bus[240]), .B(n250), .ZN(
        n252) );
  ND2D1BWP30P140LVT U298 ( .A1(n288), .A2(i_data_bus[16]), .ZN(n251) );
  ND4D1BWP30P140LVT U299 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U300 ( .A1(n1), .A2(i_data_bus[79]), .B1(n280), .B2(
        i_data_bus[47]), .ZN(n262) );
  AOI22D1BWP30P140LVT U301 ( .A1(n2), .A2(i_data_bus[111]), .B1(n281), .B2(
        i_data_bus[143]), .ZN(n261) );
  INVD1BWP30P140LVT U302 ( .I(i_data_bus[207]), .ZN(n257) );
  INVD1BWP30P140LVT U303 ( .I(i_data_bus[175]), .ZN(n255) );
  OAI22D1BWP30P140LVT U304 ( .A1(n285), .A2(n257), .B1(n256), .B2(n255), .ZN(
        n258) );
  ND2D1BWP30P140LVT U305 ( .A1(n288), .A2(i_data_bus[15]), .ZN(n259) );
  ND4D1BWP30P140LVT U306 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U307 ( .A1(n1), .A2(i_data_bus[64]), .B1(n263), .B2(
        i_data_bus[32]), .ZN(n271) );
  AOI22D1BWP30P140LVT U308 ( .A1(n2), .A2(i_data_bus[96]), .B1(n264), .B2(
        i_data_bus[128]), .ZN(n270) );
  INR2D1BWP30P140LVT U309 ( .A1(i_data_bus[192]), .B1(n285), .ZN(n266) );
  INR2D1BWP30P140LVT U310 ( .A1(i_data_bus[160]), .B1(n283), .ZN(n265) );
  AOI211D1BWP30P140LVT U311 ( .A1(i_data_bus[224]), .A2(n275), .B(n266), .C(
        n265), .ZN(n269) );
  ND2D1BWP30P140LVT U312 ( .A1(n267), .A2(i_data_bus[0]), .ZN(n268) );
  ND4D1BWP30P140LVT U313 ( .A1(n271), .A2(n270), .A3(n269), .A4(n268), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U314 ( .A1(n1), .A2(i_data_bus[78]), .B1(n280), .B2(
        i_data_bus[46]), .ZN(n279) );
  AOI22D1BWP30P140LVT U315 ( .A1(n2), .A2(i_data_bus[110]), .B1(n281), .B2(
        i_data_bus[142]), .ZN(n278) );
  INVD1BWP30P140LVT U316 ( .I(i_data_bus[206]), .ZN(n273) );
  INVD1BWP30P140LVT U317 ( .I(i_data_bus[174]), .ZN(n272) );
  OAI22D1BWP30P140LVT U318 ( .A1(n285), .A2(n273), .B1(n283), .B2(n272), .ZN(
        n274) );
  ND2D1BWP30P140LVT U319 ( .A1(n288), .A2(i_data_bus[14]), .ZN(n276) );
  ND4D1BWP30P140LVT U320 ( .A1(n279), .A2(n278), .A3(n277), .A4(n276), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U321 ( .A1(n1), .A2(i_data_bus[77]), .B1(n280), .B2(
        i_data_bus[45]), .ZN(n292) );
  AOI22D1BWP30P140LVT U322 ( .A1(n2), .A2(i_data_bus[109]), .B1(n281), .B2(
        i_data_bus[141]), .ZN(n291) );
  INVD1BWP30P140LVT U323 ( .I(i_data_bus[205]), .ZN(n284) );
  INVD1BWP30P140LVT U324 ( .I(i_data_bus[173]), .ZN(n282) );
  OAI22D1BWP30P140LVT U325 ( .A1(n285), .A2(n284), .B1(n283), .B2(n282), .ZN(
        n286) );
  ND2D1BWP30P140LVT U326 ( .A1(n288), .A2(i_data_bus[13]), .ZN(n289) );
  ND4D1BWP30P140LVT U327 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_7 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n24), .ZN(n287) );
  BUFFD4BWP30P140LVT U4 ( .I(n58), .Z(n276) );
  INVD1BWP30P140LVT U5 ( .I(n12), .ZN(n110) );
  INR2D1BWP30P140LVT U6 ( .A1(n11), .B1(n10), .ZN(n12) );
  CKND2D3BWP30P140LVT U7 ( .A1(n30), .A2(n29), .ZN(n46) );
  CKND2D3BWP30P140LVT U8 ( .A1(n9), .A2(n15), .ZN(n97) );
  AO22D1BWP30P140LVT U9 ( .A1(n155), .A2(i_data_bus[71]), .B1(n284), .B2(
        i_data_bus[39]), .Z(n2) );
  INVD3BWP30P140LVT U10 ( .I(n64), .ZN(n1) );
  IND4D1BWP30P140LVT U11 ( .A1(n2), .B1(n188), .B2(n187), .B3(n186), .ZN(N376)
         );
  INVD3BWP30P140LVT U12 ( .I(n65), .ZN(n285) );
  BUFFD4BWP30P140LVT U13 ( .I(n97), .Z(n289) );
  ND2OPTIBD2BWP30P140LVT U14 ( .A1(n23), .A2(n22), .ZN(n58) );
  ND2D1BWP30P140LVT U15 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n20) );
  INVD1BWP30P140LVT U16 ( .I(n41), .ZN(n65) );
  ND2D1BWP30P140LVT U17 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n34) );
  NR2D1BWP30P140LVT U18 ( .A1(n28), .A2(i_cmd[4]), .ZN(n30) );
  AO22D1BWP30P140LVT U19 ( .A1(n155), .A2(i_data_bus[70]), .B1(n284), .B2(
        i_data_bus[38]), .Z(n3) );
  OAI22D1BWP30P140LVT U20 ( .A1(n289), .A2(n184), .B1(n287), .B2(n183), .ZN(
        n185) );
  IND4D1BWP30P140LVT U21 ( .A1(n3), .B1(n182), .B2(n181), .B3(n180), .ZN(N375)
         );
  INR2D6BWP30P140LVT U22 ( .A1(n47), .B1(n46), .ZN(n284) );
  OR2D1BWP30P140LVT U23 ( .A1(n46), .A2(n33), .Z(n64) );
  INVD1BWP30P140LVT U24 ( .I(n51), .ZN(n69) );
  INVD2BWP30P140LVT U25 ( .I(n110), .ZN(n291) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n61), .A2(n60), .Z(n4) );
  INVD2BWP30P140LVT U27 ( .I(i_cmd[7]), .ZN(n17) );
  INR4D0BWP30P140LVT U28 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n17), .ZN(n11) );
  INVD1BWP30P140LVT U29 ( .I(i_cmd[1]), .ZN(n5) );
  INVD2BWP30P140LVT U30 ( .I(i_cmd[2]), .ZN(n42) );
  ND2OPTIBD1BWP30P140LVT U31 ( .A1(n5), .A2(n42), .ZN(n32) );
  OR2D1BWP30P140LVT U32 ( .A1(n32), .A2(i_cmd[4]), .Z(n19) );
  INVD1BWP30P140LVT U33 ( .I(rst), .ZN(n6) );
  ND2D1BWP30P140LVT U34 ( .A1(n6), .A2(i_en), .ZN(n35) );
  NR2D1BWP30P140LVT U35 ( .A1(i_cmd[0]), .A2(n35), .ZN(n8) );
  INVD1BWP30P140LVT U36 ( .I(i_cmd[3]), .ZN(n7) );
  ND2OPTIBD1BWP30P140LVT U37 ( .A1(n8), .A2(n7), .ZN(n21) );
  NR2OPTPAD1BWP30P140LVT U38 ( .A1(n19), .A2(n21), .ZN(n9) );
  INVD2BWP30P140LVT U39 ( .I(n9), .ZN(n10) );
  INVD2BWP30P140LVT U40 ( .I(n110), .ZN(n279) );
  NR2D1BWP30P140LVT U41 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n14) );
  CKAN2D1BWP30P140LVT U42 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n13) );
  AN2D2BWP30P140LVT U43 ( .A1(n14), .A2(n13), .Z(n15) );
  INVD1BWP30P140LVT U44 ( .I(i_data_bus[206]), .ZN(n26) );
  INVD1BWP30P140LVT U45 ( .I(i_cmd[6]), .ZN(n18) );
  ND2OPTIBD2BWP30P140LVT U46 ( .A1(n18), .A2(n17), .ZN(n37) );
  NR2D1BWP30P140LVT U47 ( .A1(n37), .A2(n19), .ZN(n23) );
  NR2D1BWP30P140LVT U48 ( .A1(n21), .A2(n20), .ZN(n22) );
  INVD2BWP30P140LVT U49 ( .I(n58), .ZN(n24) );
  INVD1BWP30P140LVT U50 ( .I(i_data_bus[174]), .ZN(n25) );
  OAI22D1BWP30P140LVT U51 ( .A1(n158), .A2(n26), .B1(n287), .B2(n25), .ZN(n27)
         );
  AOI21D1BWP30P140LVT U52 ( .A1(n279), .A2(i_data_bus[238]), .B(n27), .ZN(n57)
         );
  OR2D1BWP30P140LVT U53 ( .A1(i_cmd[0]), .A2(n35), .Z(n28) );
  NR2OPTPAD1BWP30P140LVT U54 ( .A1(i_cmd[5]), .A2(n37), .ZN(n29) );
  ND2OPTIBD1BWP30P140LVT U55 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n31) );
  OR2D1BWP30P140LVT U56 ( .A1(n32), .A2(n31), .Z(n33) );
  NR2D1BWP30P140LVT U57 ( .A1(n34), .A2(i_cmd[0]), .ZN(n40) );
  OR2D1BWP30P140LVT U58 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n45) );
  INVD1BWP30P140LVT U59 ( .I(n45), .ZN(n39) );
  OR2D1BWP30P140LVT U60 ( .A1(i_cmd[1]), .A2(n35), .Z(n36) );
  NR3D0P7BWP30P140LVT U61 ( .A1(n37), .A2(i_cmd[5]), .A3(n36), .ZN(n38) );
  ND2OPTIBD1BWP30P140LVT U62 ( .A1(n39), .A2(n38), .ZN(n49) );
  INR2D1BWP30P140LVT U63 ( .A1(n40), .B1(n49), .ZN(n41) );
  AOI22D1BWP30P140LVT U64 ( .A1(n1), .A2(i_data_bus[110]), .B1(n285), .B2(
        i_data_bus[142]), .ZN(n56) );
  INR4D1BWP30P140LVT U65 ( .A1(i_valid[2]), .B1(i_cmd[1]), .B2(i_cmd[3]), .B3(
        n42), .ZN(n43) );
  INR2D4BWP30P140LVT U66 ( .A1(n43), .B1(n46), .ZN(n155) );
  ND2D1BWP30P140LVT U67 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n44) );
  NR2OPTPAD1BWP30P140LVT U68 ( .A1(n45), .A2(n44), .ZN(n47) );
  AOI22D1BWP30P140LVT U69 ( .A1(n155), .A2(i_data_bus[78]), .B1(n284), .B2(
        i_data_bus[46]), .ZN(n53) );
  INVD1BWP30P140LVT U70 ( .I(i_cmd[0]), .ZN(n48) );
  INR3D0BWP30P140LVT U71 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n48), .ZN(n50)
         );
  INR2D1BWP30P140LVT U72 ( .A1(n50), .B1(n49), .ZN(n51) );
  INVD2BWP30P140LVT U73 ( .I(n69), .ZN(n292) );
  ND2D1BWP30P140LVT U74 ( .A1(n292), .A2(i_data_bus[14]), .ZN(n52) );
  ND2D1BWP30P140LVT U75 ( .A1(n53), .A2(n52), .ZN(n54) );
  INVD1BWP30P140LVT U76 ( .I(n54), .ZN(n55) );
  ND3D1BWP30P140LVT U77 ( .A1(n57), .A2(n56), .A3(n55), .ZN(N383) );
  INVD2BWP30P140LVT U78 ( .I(n97), .ZN(n111) );
  INVD1BWP30P140LVT U79 ( .I(n276), .ZN(n59) );
  NR4D0BWP30P140LVT U80 ( .A1(n207), .A2(n111), .A3(n59), .A4(n291), .ZN(n63)
         );
  NR2D1BWP30P140LVT U81 ( .A1(n1), .A2(n285), .ZN(n62) );
  INVD1BWP30P140LVT U82 ( .I(n155), .ZN(n61) );
  INVD1BWP30P140LVT U83 ( .I(n284), .ZN(n60) );
  ND3D1BWP30P140LVT U84 ( .A1(n63), .A2(n62), .A3(n4), .ZN(N402) );
  AOI22D1BWP30P140LVT U85 ( .A1(n155), .A2(i_data_bus[65]), .B1(n284), .B2(
        i_data_bus[33]), .ZN(n73) );
  INVD2BWP30P140LVT U86 ( .I(n65), .ZN(n203) );
  AOI22D1BWP30P140LVT U87 ( .A1(n1), .A2(i_data_bus[97]), .B1(n203), .B2(
        i_data_bus[129]), .ZN(n72) );
  INVD1BWP30P140LVT U88 ( .I(i_data_bus[193]), .ZN(n67) );
  INVD1BWP30P140LVT U89 ( .I(i_data_bus[161]), .ZN(n66) );
  OAI22D1BWP30P140LVT U90 ( .A1(n97), .A2(n67), .B1(n287), .B2(n66), .ZN(n68)
         );
  AOI21D1BWP30P140LVT U91 ( .A1(n291), .A2(i_data_bus[225]), .B(n68), .ZN(n71)
         );
  INVD2BWP30P140LVT U92 ( .I(n69), .ZN(n207) );
  ND2D1BWP30P140LVT U93 ( .A1(n207), .A2(i_data_bus[1]), .ZN(n70) );
  ND4D1BWP30P140LVT U94 ( .A1(n73), .A2(n72), .A3(n71), .A4(n70), .ZN(N370) );
  AOI22D1BWP30P140LVT U95 ( .A1(n155), .A2(i_data_bus[68]), .B1(n284), .B2(
        i_data_bus[36]), .ZN(n80) );
  AOI22D1BWP30P140LVT U96 ( .A1(n1), .A2(i_data_bus[100]), .B1(n203), .B2(
        i_data_bus[132]), .ZN(n79) );
  INVD1BWP30P140LVT U97 ( .I(i_data_bus[196]), .ZN(n75) );
  INVD1BWP30P140LVT U98 ( .I(i_data_bus[164]), .ZN(n74) );
  OAI22D1BWP30P140LVT U99 ( .A1(n97), .A2(n75), .B1(n287), .B2(n74), .ZN(n76)
         );
  AOI21D1BWP30P140LVT U100 ( .A1(n291), .A2(i_data_bus[228]), .B(n76), .ZN(n78) );
  ND2D1BWP30P140LVT U101 ( .A1(n207), .A2(i_data_bus[4]), .ZN(n77) );
  ND4D1BWP30P140LVT U102 ( .A1(n80), .A2(n79), .A3(n78), .A4(n77), .ZN(N373)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n155), .A2(i_data_bus[67]), .B1(n284), .B2(
        i_data_bus[35]), .ZN(n87) );
  AOI22D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[99]), .B1(n203), .B2(
        i_data_bus[131]), .ZN(n86) );
  INVD1BWP30P140LVT U105 ( .I(i_data_bus[195]), .ZN(n82) );
  INVD1BWP30P140LVT U106 ( .I(i_data_bus[163]), .ZN(n81) );
  OAI22D1BWP30P140LVT U107 ( .A1(n97), .A2(n82), .B1(n287), .B2(n81), .ZN(n83)
         );
  AOI21D1BWP30P140LVT U108 ( .A1(n291), .A2(i_data_bus[227]), .B(n83), .ZN(n85) );
  ND2D1BWP30P140LVT U109 ( .A1(n207), .A2(i_data_bus[3]), .ZN(n84) );
  ND4D1BWP30P140LVT U110 ( .A1(n87), .A2(n86), .A3(n85), .A4(n84), .ZN(N372)
         );
  AOI22D1BWP30P140LVT U111 ( .A1(n155), .A2(i_data_bus[69]), .B1(n284), .B2(
        i_data_bus[37]), .ZN(n94) );
  AOI22D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[101]), .B1(n203), .B2(
        i_data_bus[133]), .ZN(n93) );
  INVD1BWP30P140LVT U113 ( .I(i_data_bus[197]), .ZN(n89) );
  INVD1BWP30P140LVT U114 ( .I(i_data_bus[165]), .ZN(n88) );
  OAI22D1BWP30P140LVT U115 ( .A1(n97), .A2(n89), .B1(n287), .B2(n88), .ZN(n90)
         );
  AOI21D1BWP30P140LVT U116 ( .A1(n291), .A2(i_data_bus[229]), .B(n90), .ZN(n92) );
  ND2D1BWP30P140LVT U117 ( .A1(n207), .A2(i_data_bus[5]), .ZN(n91) );
  ND4D1BWP30P140LVT U118 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U119 ( .A1(n155), .A2(i_data_bus[66]), .B1(n284), .B2(
        i_data_bus[34]), .ZN(n102) );
  AOI22D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[98]), .B1(n203), .B2(
        i_data_bus[130]), .ZN(n101) );
  INVD1BWP30P140LVT U121 ( .I(i_data_bus[194]), .ZN(n96) );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[162]), .ZN(n95) );
  OAI22D1BWP30P140LVT U123 ( .A1(n97), .A2(n96), .B1(n287), .B2(n95), .ZN(n98)
         );
  AOI21D1BWP30P140LVT U124 ( .A1(n291), .A2(i_data_bus[226]), .B(n98), .ZN(
        n100) );
  ND2D1BWP30P140LVT U125 ( .A1(n207), .A2(i_data_bus[2]), .ZN(n99) );
  ND4D1BWP30P140LVT U126 ( .A1(n102), .A2(n101), .A3(n100), .A4(n99), .ZN(N371) );
  AOI22D1BWP30P140LVT U127 ( .A1(n155), .A2(i_data_bus[76]), .B1(n284), .B2(
        i_data_bus[44]), .ZN(n109) );
  AOI22D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[108]), .B1(n203), .B2(
        i_data_bus[140]), .ZN(n108) );
  INVD1BWP30P140LVT U129 ( .I(i_data_bus[172]), .ZN(n104) );
  ND2D1BWP30P140LVT U130 ( .A1(n111), .A2(i_data_bus[204]), .ZN(n103) );
  OAI21D1BWP30P140LVT U131 ( .A1(n287), .A2(n104), .B(n103), .ZN(n105) );
  AOI21D1BWP30P140LVT U132 ( .A1(n291), .A2(i_data_bus[236]), .B(n105), .ZN(
        n107) );
  ND2D1BWP30P140LVT U133 ( .A1(n207), .A2(i_data_bus[12]), .ZN(n106) );
  ND4D1BWP30P140LVT U134 ( .A1(n109), .A2(n108), .A3(n107), .A4(n106), .ZN(
        N381) );
  AOI22D1BWP30P140LVT U135 ( .A1(n155), .A2(i_data_bus[93]), .B1(n284), .B2(
        i_data_bus[61]), .ZN(n118) );
  AOI22D1BWP30P140LVT U136 ( .A1(n1), .A2(i_data_bus[125]), .B1(n285), .B2(
        i_data_bus[157]), .ZN(n117) );
  INVD2BWP30P140LVT U137 ( .I(n111), .ZN(n158) );
  INVD1BWP30P140LVT U138 ( .I(i_data_bus[221]), .ZN(n113) );
  INVD1BWP30P140LVT U139 ( .I(i_data_bus[189]), .ZN(n112) );
  OAI22D1BWP30P140LVT U140 ( .A1(n158), .A2(n113), .B1(n276), .B2(n112), .ZN(
        n114) );
  AOI21D1BWP30P140LVT U141 ( .A1(n291), .A2(i_data_bus[253]), .B(n114), .ZN(
        n116) );
  ND2D1BWP30P140LVT U142 ( .A1(n207), .A2(i_data_bus[29]), .ZN(n115) );
  ND4D1BWP30P140LVT U143 ( .A1(n118), .A2(n117), .A3(n116), .A4(n115), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U144 ( .A1(n155), .A2(i_data_bus[92]), .B1(n284), .B2(
        i_data_bus[60]), .ZN(n125) );
  AOI22D1BWP30P140LVT U145 ( .A1(n1), .A2(i_data_bus[124]), .B1(n285), .B2(
        i_data_bus[156]), .ZN(n124) );
  INVD1BWP30P140LVT U146 ( .I(i_data_bus[220]), .ZN(n120) );
  INVD1BWP30P140LVT U147 ( .I(i_data_bus[188]), .ZN(n119) );
  OAI22D1BWP30P140LVT U148 ( .A1(n158), .A2(n120), .B1(n276), .B2(n119), .ZN(
        n121) );
  AOI21D1BWP30P140LVT U149 ( .A1(n291), .A2(i_data_bus[252]), .B(n121), .ZN(
        n123) );
  ND2D1BWP30P140LVT U150 ( .A1(n207), .A2(i_data_bus[28]), .ZN(n122) );
  ND4D1BWP30P140LVT U151 ( .A1(n125), .A2(n124), .A3(n123), .A4(n122), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U152 ( .A1(n155), .A2(i_data_bus[94]), .B1(n284), .B2(
        i_data_bus[62]), .ZN(n132) );
  AOI22D1BWP30P140LVT U153 ( .A1(n1), .A2(i_data_bus[126]), .B1(n285), .B2(
        i_data_bus[158]), .ZN(n131) );
  INVD1BWP30P140LVT U154 ( .I(i_data_bus[222]), .ZN(n127) );
  INVD1BWP30P140LVT U155 ( .I(i_data_bus[190]), .ZN(n126) );
  OAI22D1BWP30P140LVT U156 ( .A1(n158), .A2(n127), .B1(n276), .B2(n126), .ZN(
        n128) );
  AOI21D1BWP30P140LVT U157 ( .A1(n291), .A2(i_data_bus[254]), .B(n128), .ZN(
        n130) );
  ND2D1BWP30P140LVT U158 ( .A1(n207), .A2(i_data_bus[30]), .ZN(n129) );
  ND4D1BWP30P140LVT U159 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U160 ( .A1(n155), .A2(i_data_bus[91]), .B1(n284), .B2(
        i_data_bus[59]), .ZN(n139) );
  AOI22D1BWP30P140LVT U161 ( .A1(n1), .A2(i_data_bus[123]), .B1(n285), .B2(
        i_data_bus[155]), .ZN(n138) );
  INVD1BWP30P140LVT U162 ( .I(i_data_bus[219]), .ZN(n134) );
  INVD1BWP30P140LVT U163 ( .I(i_data_bus[187]), .ZN(n133) );
  OAI22D1BWP30P140LVT U164 ( .A1(n158), .A2(n134), .B1(n276), .B2(n133), .ZN(
        n135) );
  AOI21D1BWP30P140LVT U165 ( .A1(n279), .A2(i_data_bus[251]), .B(n135), .ZN(
        n137) );
  ND2D1BWP30P140LVT U166 ( .A1(n207), .A2(i_data_bus[27]), .ZN(n136) );
  ND4D1BWP30P140LVT U167 ( .A1(n139), .A2(n138), .A3(n137), .A4(n136), .ZN(
        N396) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n155), .A2(i_data_bus[89]), .Z(n140) );
  AOI21D1BWP30P140LVT U169 ( .A1(n284), .A2(i_data_bus[57]), .B(n140), .ZN(
        n147) );
  AOI22D1BWP30P140LVT U170 ( .A1(n1), .A2(i_data_bus[121]), .B1(n285), .B2(
        i_data_bus[153]), .ZN(n146) );
  INVD1BWP30P140LVT U171 ( .I(i_data_bus[217]), .ZN(n142) );
  INVD1BWP30P140LVT U172 ( .I(i_data_bus[185]), .ZN(n141) );
  OAI22D1BWP30P140LVT U173 ( .A1(n158), .A2(n142), .B1(n276), .B2(n141), .ZN(
        n143) );
  AOI21D1BWP30P140LVT U174 ( .A1(n279), .A2(i_data_bus[249]), .B(n143), .ZN(
        n145) );
  ND2D1BWP30P140LVT U175 ( .A1(n292), .A2(i_data_bus[25]), .ZN(n144) );
  ND4D1BWP30P140LVT U176 ( .A1(n147), .A2(n146), .A3(n145), .A4(n144), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U177 ( .A1(n155), .A2(i_data_bus[90]), .B1(n284), .B2(
        i_data_bus[58]), .ZN(n154) );
  AOI22D1BWP30P140LVT U178 ( .A1(n1), .A2(i_data_bus[122]), .B1(n285), .B2(
        i_data_bus[154]), .ZN(n153) );
  INVD1BWP30P140LVT U179 ( .I(i_data_bus[218]), .ZN(n149) );
  INVD1BWP30P140LVT U180 ( .I(i_data_bus[186]), .ZN(n148) );
  OAI22D1BWP30P140LVT U181 ( .A1(n158), .A2(n149), .B1(n276), .B2(n148), .ZN(
        n150) );
  AOI21D1BWP30P140LVT U182 ( .A1(n279), .A2(i_data_bus[250]), .B(n150), .ZN(
        n152) );
  ND2D1BWP30P140LVT U183 ( .A1(n207), .A2(i_data_bus[26]), .ZN(n151) );
  ND4D1BWP30P140LVT U184 ( .A1(n154), .A2(n153), .A3(n152), .A4(n151), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U185 ( .A1(n155), .A2(i_data_bus[95]), .B1(n284), .B2(
        i_data_bus[63]), .ZN(n163) );
  AOI22D1BWP30P140LVT U186 ( .A1(n1), .A2(i_data_bus[127]), .B1(n285), .B2(
        i_data_bus[159]), .ZN(n162) );
  INVD1BWP30P140LVT U187 ( .I(i_data_bus[223]), .ZN(n157) );
  INVD1BWP30P140LVT U188 ( .I(i_data_bus[191]), .ZN(n156) );
  OAI22D1BWP30P140LVT U189 ( .A1(n158), .A2(n157), .B1(n276), .B2(n156), .ZN(
        n159) );
  AOI21D1BWP30P140LVT U190 ( .A1(n291), .A2(i_data_bus[255]), .B(n159), .ZN(
        n161) );
  ND2D1BWP30P140LVT U191 ( .A1(n207), .A2(i_data_bus[31]), .ZN(n160) );
  ND4D1BWP30P140LVT U192 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U193 ( .A1(n155), .A2(i_data_bus[64]), .B1(n284), .B2(
        i_data_bus[32]), .ZN(n169) );
  AOI22D1BWP30P140LVT U194 ( .A1(n1), .A2(i_data_bus[96]), .B1(n203), .B2(
        i_data_bus[128]), .ZN(n168) );
  INR2D1BWP30P140LVT U195 ( .A1(i_data_bus[192]), .B1(n289), .ZN(n165) );
  INR2D1BWP30P140LVT U196 ( .A1(i_data_bus[160]), .B1(n287), .ZN(n164) );
  AOI211D1BWP30P140LVT U197 ( .A1(i_data_bus[224]), .A2(n291), .B(n165), .C(
        n164), .ZN(n167) );
  ND2D1BWP30P140LVT U198 ( .A1(n207), .A2(i_data_bus[0]), .ZN(n166) );
  ND4D1BWP30P140LVT U199 ( .A1(n169), .A2(n168), .A3(n167), .A4(n166), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U200 ( .A1(n155), .A2(i_data_bus[72]), .B1(n284), .B2(
        i_data_bus[40]), .ZN(n176) );
  AOI22D1BWP30P140LVT U201 ( .A1(n1), .A2(i_data_bus[104]), .B1(n203), .B2(
        i_data_bus[136]), .ZN(n175) );
  INVD1BWP30P140LVT U202 ( .I(i_data_bus[200]), .ZN(n171) );
  INVD1BWP30P140LVT U203 ( .I(i_data_bus[168]), .ZN(n170) );
  OAI22D1BWP30P140LVT U204 ( .A1(n289), .A2(n171), .B1(n287), .B2(n170), .ZN(
        n172) );
  AOI21D1BWP30P140LVT U205 ( .A1(n279), .A2(i_data_bus[232]), .B(n172), .ZN(
        n174) );
  ND2D1BWP30P140LVT U206 ( .A1(n207), .A2(i_data_bus[8]), .ZN(n173) );
  ND4D1BWP30P140LVT U207 ( .A1(n176), .A2(n175), .A3(n174), .A4(n173), .ZN(
        N377) );
  AOI22D1BWP30P140LVT U208 ( .A1(n1), .A2(i_data_bus[102]), .B1(n203), .B2(
        i_data_bus[134]), .ZN(n182) );
  INVD1BWP30P140LVT U209 ( .I(i_data_bus[198]), .ZN(n178) );
  INVD1BWP30P140LVT U210 ( .I(i_data_bus[166]), .ZN(n177) );
  OAI22D1BWP30P140LVT U211 ( .A1(n289), .A2(n178), .B1(n287), .B2(n177), .ZN(
        n179) );
  AOI21D1BWP30P140LVT U212 ( .A1(n291), .A2(i_data_bus[230]), .B(n179), .ZN(
        n181) );
  ND2D1BWP30P140LVT U213 ( .A1(n207), .A2(i_data_bus[6]), .ZN(n180) );
  AOI22D1BWP30P140LVT U214 ( .A1(n1), .A2(i_data_bus[103]), .B1(n203), .B2(
        i_data_bus[135]), .ZN(n188) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[199]), .ZN(n184) );
  INVD1BWP30P140LVT U216 ( .I(i_data_bus[167]), .ZN(n183) );
  AOI21D1BWP30P140LVT U217 ( .A1(n291), .A2(i_data_bus[231]), .B(n185), .ZN(
        n187) );
  ND2D1BWP30P140LVT U218 ( .A1(n207), .A2(i_data_bus[7]), .ZN(n186) );
  AOI22D1BWP30P140LVT U219 ( .A1(n155), .A2(i_data_bus[73]), .B1(n284), .B2(
        i_data_bus[41]), .ZN(n195) );
  AOI22D1BWP30P140LVT U220 ( .A1(n1), .A2(i_data_bus[105]), .B1(n203), .B2(
        i_data_bus[137]), .ZN(n194) );
  INVD1BWP30P140LVT U221 ( .I(i_data_bus[201]), .ZN(n190) );
  INVD1BWP30P140LVT U222 ( .I(i_data_bus[169]), .ZN(n189) );
  OAI22D1BWP30P140LVT U223 ( .A1(n289), .A2(n190), .B1(n287), .B2(n189), .ZN(
        n191) );
  AOI21D1BWP30P140LVT U224 ( .A1(n291), .A2(i_data_bus[233]), .B(n191), .ZN(
        n193) );
  ND2D1BWP30P140LVT U225 ( .A1(n207), .A2(i_data_bus[9]), .ZN(n192) );
  ND4D1BWP30P140LVT U226 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U227 ( .A1(n155), .A2(i_data_bus[74]), .B1(n284), .B2(
        i_data_bus[42]), .ZN(n202) );
  AOI22D1BWP30P140LVT U228 ( .A1(n1), .A2(i_data_bus[106]), .B1(n203), .B2(
        i_data_bus[138]), .ZN(n201) );
  INVD1BWP30P140LVT U229 ( .I(i_data_bus[202]), .ZN(n197) );
  INVD1BWP30P140LVT U230 ( .I(i_data_bus[170]), .ZN(n196) );
  OAI22D1BWP30P140LVT U231 ( .A1(n289), .A2(n197), .B1(n287), .B2(n196), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U232 ( .A1(n291), .A2(i_data_bus[234]), .B(n198), .ZN(
        n200) );
  ND2D1BWP30P140LVT U233 ( .A1(n207), .A2(i_data_bus[10]), .ZN(n199) );
  ND4D1BWP30P140LVT U234 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(
        N379) );
  AOI22D1BWP30P140LVT U235 ( .A1(n155), .A2(i_data_bus[75]), .B1(n284), .B2(
        i_data_bus[43]), .ZN(n211) );
  AOI22D1BWP30P140LVT U236 ( .A1(n1), .A2(i_data_bus[107]), .B1(n203), .B2(
        i_data_bus[139]), .ZN(n210) );
  INVD1BWP30P140LVT U237 ( .I(i_data_bus[203]), .ZN(n205) );
  INVD1BWP30P140LVT U238 ( .I(i_data_bus[171]), .ZN(n204) );
  OAI22D1BWP30P140LVT U239 ( .A1(n289), .A2(n205), .B1(n287), .B2(n204), .ZN(
        n206) );
  AOI21D1BWP30P140LVT U240 ( .A1(n291), .A2(i_data_bus[235]), .B(n206), .ZN(
        n209) );
  ND2D1BWP30P140LVT U241 ( .A1(n207), .A2(i_data_bus[11]), .ZN(n208) );
  ND4D1BWP30P140LVT U242 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .ZN(
        N380) );
  AOI22D1BWP30P140LVT U243 ( .A1(n155), .A2(i_data_bus[80]), .B1(n284), .B2(
        i_data_bus[48]), .ZN(n218) );
  AOI22D1BWP30P140LVT U244 ( .A1(n1), .A2(i_data_bus[112]), .B1(n285), .B2(
        i_data_bus[144]), .ZN(n217) );
  INVD1BWP30P140LVT U245 ( .I(i_data_bus[208]), .ZN(n213) );
  INVD1BWP30P140LVT U246 ( .I(i_data_bus[176]), .ZN(n212) );
  OAI22D1BWP30P140LVT U247 ( .A1(n289), .A2(n213), .B1(n276), .B2(n212), .ZN(
        n214) );
  AOI21D1BWP30P140LVT U248 ( .A1(n279), .A2(i_data_bus[240]), .B(n214), .ZN(
        n216) );
  ND2D1BWP30P140LVT U249 ( .A1(n292), .A2(i_data_bus[16]), .ZN(n215) );
  ND4D1BWP30P140LVT U250 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U251 ( .A1(n155), .A2(i_data_bus[87]), .B1(n284), .B2(
        i_data_bus[55]), .ZN(n225) );
  AOI22D1BWP30P140LVT U252 ( .A1(n1), .A2(i_data_bus[119]), .B1(n285), .B2(
        i_data_bus[151]), .ZN(n224) );
  INVD1BWP30P140LVT U253 ( .I(i_data_bus[215]), .ZN(n220) );
  INVD1BWP30P140LVT U254 ( .I(i_data_bus[183]), .ZN(n219) );
  OAI22D1BWP30P140LVT U255 ( .A1(n289), .A2(n220), .B1(n276), .B2(n219), .ZN(
        n221) );
  AOI21D1BWP30P140LVT U256 ( .A1(n279), .A2(i_data_bus[247]), .B(n221), .ZN(
        n223) );
  ND2D1BWP30P140LVT U257 ( .A1(n292), .A2(i_data_bus[23]), .ZN(n222) );
  ND4D1BWP30P140LVT U258 ( .A1(n225), .A2(n224), .A3(n223), .A4(n222), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U259 ( .A1(n155), .A2(i_data_bus[85]), .B1(n284), .B2(
        i_data_bus[53]), .ZN(n232) );
  AOI22D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[117]), .B1(n285), .B2(
        i_data_bus[149]), .ZN(n231) );
  INVD1BWP30P140LVT U261 ( .I(i_data_bus[213]), .ZN(n227) );
  INVD1BWP30P140LVT U262 ( .I(i_data_bus[181]), .ZN(n226) );
  OAI22D1BWP30P140LVT U263 ( .A1(n289), .A2(n227), .B1(n276), .B2(n226), .ZN(
        n228) );
  AOI21D1BWP30P140LVT U264 ( .A1(n279), .A2(i_data_bus[245]), .B(n228), .ZN(
        n230) );
  ND2D1BWP30P140LVT U265 ( .A1(n292), .A2(i_data_bus[21]), .ZN(n229) );
  ND4D1BWP30P140LVT U266 ( .A1(n232), .A2(n231), .A3(n230), .A4(n229), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U267 ( .A1(n155), .A2(i_data_bus[88]), .B1(n284), .B2(
        i_data_bus[56]), .ZN(n239) );
  AOI22D1BWP30P140LVT U268 ( .A1(n1), .A2(i_data_bus[120]), .B1(n285), .B2(
        i_data_bus[152]), .ZN(n238) );
  INVD1BWP30P140LVT U269 ( .I(i_data_bus[216]), .ZN(n234) );
  INVD1BWP30P140LVT U270 ( .I(i_data_bus[184]), .ZN(n233) );
  OAI22D1BWP30P140LVT U271 ( .A1(n289), .A2(n234), .B1(n276), .B2(n233), .ZN(
        n235) );
  AOI21D1BWP30P140LVT U272 ( .A1(n279), .A2(i_data_bus[248]), .B(n235), .ZN(
        n237) );
  ND2D1BWP30P140LVT U273 ( .A1(n292), .A2(i_data_bus[24]), .ZN(n236) );
  ND4D1BWP30P140LVT U274 ( .A1(n239), .A2(n238), .A3(n237), .A4(n236), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U275 ( .A1(n155), .A2(i_data_bus[83]), .B1(n284), .B2(
        i_data_bus[51]), .ZN(n246) );
  AOI22D1BWP30P140LVT U276 ( .A1(n1), .A2(i_data_bus[115]), .B1(n285), .B2(
        i_data_bus[147]), .ZN(n245) );
  INVD1BWP30P140LVT U277 ( .I(i_data_bus[211]), .ZN(n241) );
  INVD1BWP30P140LVT U278 ( .I(i_data_bus[179]), .ZN(n240) );
  OAI22D1BWP30P140LVT U279 ( .A1(n289), .A2(n241), .B1(n276), .B2(n240), .ZN(
        n242) );
  AOI21D1BWP30P140LVT U280 ( .A1(n279), .A2(i_data_bus[243]), .B(n242), .ZN(
        n244) );
  ND2D1BWP30P140LVT U281 ( .A1(n292), .A2(i_data_bus[19]), .ZN(n243) );
  ND4D1BWP30P140LVT U282 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U283 ( .A1(n155), .A2(i_data_bus[84]), .B1(n284), .B2(
        i_data_bus[52]), .ZN(n253) );
  AOI22D1BWP30P140LVT U284 ( .A1(n1), .A2(i_data_bus[116]), .B1(n285), .B2(
        i_data_bus[148]), .ZN(n252) );
  INVD1BWP30P140LVT U285 ( .I(i_data_bus[212]), .ZN(n248) );
  INVD1BWP30P140LVT U286 ( .I(i_data_bus[180]), .ZN(n247) );
  OAI22D1BWP30P140LVT U287 ( .A1(n289), .A2(n248), .B1(n276), .B2(n247), .ZN(
        n249) );
  AOI21D1BWP30P140LVT U288 ( .A1(n279), .A2(i_data_bus[244]), .B(n249), .ZN(
        n251) );
  ND2D1BWP30P140LVT U289 ( .A1(n292), .A2(i_data_bus[20]), .ZN(n250) );
  ND4D1BWP30P140LVT U290 ( .A1(n253), .A2(n252), .A3(n251), .A4(n250), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U291 ( .A1(n155), .A2(i_data_bus[81]), .B1(n284), .B2(
        i_data_bus[49]), .ZN(n260) );
  AOI22D1BWP30P140LVT U292 ( .A1(n1), .A2(i_data_bus[113]), .B1(n285), .B2(
        i_data_bus[145]), .ZN(n259) );
  INVD1BWP30P140LVT U293 ( .I(i_data_bus[209]), .ZN(n255) );
  INVD1BWP30P140LVT U294 ( .I(i_data_bus[177]), .ZN(n254) );
  OAI22D1BWP30P140LVT U295 ( .A1(n289), .A2(n255), .B1(n276), .B2(n254), .ZN(
        n256) );
  AOI21D1BWP30P140LVT U296 ( .A1(n279), .A2(i_data_bus[241]), .B(n256), .ZN(
        n258) );
  ND2D1BWP30P140LVT U297 ( .A1(n292), .A2(i_data_bus[17]), .ZN(n257) );
  ND4D1BWP30P140LVT U298 ( .A1(n260), .A2(n259), .A3(n258), .A4(n257), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U299 ( .A1(n155), .A2(i_data_bus[82]), .B1(n284), .B2(
        i_data_bus[50]), .ZN(n267) );
  AOI22D1BWP30P140LVT U300 ( .A1(n1), .A2(i_data_bus[114]), .B1(n285), .B2(
        i_data_bus[146]), .ZN(n266) );
  INVD1BWP30P140LVT U301 ( .I(i_data_bus[210]), .ZN(n262) );
  INVD1BWP30P140LVT U302 ( .I(i_data_bus[178]), .ZN(n261) );
  OAI22D1BWP30P140LVT U303 ( .A1(n289), .A2(n262), .B1(n276), .B2(n261), .ZN(
        n263) );
  AOI21D1BWP30P140LVT U304 ( .A1(n279), .A2(i_data_bus[242]), .B(n263), .ZN(
        n265) );
  ND2D1BWP30P140LVT U305 ( .A1(n292), .A2(i_data_bus[18]), .ZN(n264) );
  ND4D1BWP30P140LVT U306 ( .A1(n267), .A2(n266), .A3(n265), .A4(n264), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U307 ( .A1(n155), .A2(i_data_bus[86]), .B1(n284), .B2(
        i_data_bus[54]), .ZN(n274) );
  AOI22D1BWP30P140LVT U308 ( .A1(n1), .A2(i_data_bus[118]), .B1(n285), .B2(
        i_data_bus[150]), .ZN(n273) );
  INVD1BWP30P140LVT U309 ( .I(i_data_bus[214]), .ZN(n269) );
  INVD1BWP30P140LVT U310 ( .I(i_data_bus[182]), .ZN(n268) );
  OAI22D1BWP30P140LVT U311 ( .A1(n289), .A2(n269), .B1(n276), .B2(n268), .ZN(
        n270) );
  AOI21D1BWP30P140LVT U312 ( .A1(n279), .A2(i_data_bus[246]), .B(n270), .ZN(
        n272) );
  ND2D1BWP30P140LVT U313 ( .A1(n292), .A2(i_data_bus[22]), .ZN(n271) );
  ND4D1BWP30P140LVT U314 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U315 ( .A1(n155), .A2(i_data_bus[79]), .B1(n284), .B2(
        i_data_bus[47]), .ZN(n283) );
  AOI22D1BWP30P140LVT U316 ( .A1(n1), .A2(i_data_bus[111]), .B1(n285), .B2(
        i_data_bus[143]), .ZN(n282) );
  INVD1BWP30P140LVT U317 ( .I(i_data_bus[207]), .ZN(n277) );
  INVD1BWP30P140LVT U318 ( .I(i_data_bus[175]), .ZN(n275) );
  OAI22D1BWP30P140LVT U319 ( .A1(n289), .A2(n277), .B1(n276), .B2(n275), .ZN(
        n278) );
  AOI21D1BWP30P140LVT U320 ( .A1(n279), .A2(i_data_bus[239]), .B(n278), .ZN(
        n281) );
  ND2D1BWP30P140LVT U321 ( .A1(n292), .A2(i_data_bus[15]), .ZN(n280) );
  ND4D1BWP30P140LVT U322 ( .A1(n283), .A2(n282), .A3(n281), .A4(n280), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U323 ( .A1(n155), .A2(i_data_bus[77]), .B1(n284), .B2(
        i_data_bus[45]), .ZN(n296) );
  AOI22D1BWP30P140LVT U324 ( .A1(n1), .A2(i_data_bus[109]), .B1(n285), .B2(
        i_data_bus[141]), .ZN(n295) );
  INVD1BWP30P140LVT U325 ( .I(i_data_bus[205]), .ZN(n288) );
  INVD1BWP30P140LVT U326 ( .I(i_data_bus[173]), .ZN(n286) );
  OAI22D1BWP30P140LVT U327 ( .A1(n289), .A2(n288), .B1(n287), .B2(n286), .ZN(
        n290) );
  AOI21D1BWP30P140LVT U328 ( .A1(n291), .A2(i_data_bus[237]), .B(n290), .ZN(
        n294) );
  ND2D1BWP30P140LVT U329 ( .A1(n292), .A2(i_data_bus[13]), .ZN(n293) );
  ND4D1BWP30P140LVT U330 ( .A1(n296), .A2(n295), .A3(n294), .A4(n293), .ZN(
        N382) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_8 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input clk, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279;

  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(clk), .Q(o_valid[0]) );
  INVD3BWP30P140LVT U3 ( .I(n61), .ZN(n268) );
  INVD2BWP30P140LVT U4 ( .I(n14), .ZN(n259) );
  ND2OPTIBD2BWP30P140LVT U5 ( .A1(n17), .A2(n19), .ZN(n105) );
  NR2OPTPAD2BWP30P140LVT U6 ( .A1(n11), .A2(n28), .ZN(n19) );
  OR2D1BWP30P140LVT U7 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n28) );
  INVD1BWP30P140LVT U8 ( .I(n105), .ZN(n1) );
  INVD1BWP30P140LVT U9 ( .I(n243), .ZN(n2) );
  INVD3BWP30P140LVT U10 ( .I(n134), .ZN(n3) );
  NR2OPTPAD2BWP30P140LVT U11 ( .A1(n16), .A2(i_cmd[5]), .ZN(n26) );
  INVD2BWP30P140LVT U12 ( .I(n259), .ZN(n137) );
  INVD1BWP30P140LVT U13 ( .I(n48), .ZN(n56) );
  AOI21D1BWP30P140LVT U14 ( .A1(n274), .A2(i_data_bus[227]), .B(n231), .ZN(
        n233) );
  AOI21D1BWP30P140LVT U15 ( .A1(n274), .A2(i_data_bus[228]), .B(n224), .ZN(
        n226) );
  AOI21D1BWP30P140LVT U16 ( .A1(n274), .A2(i_data_bus[237]), .B(n273), .ZN(
        n277) );
  OR2D1BWP30P140LVT U17 ( .A1(n40), .A2(n29), .Z(n134) );
  INVD1BWP30P140LVT U18 ( .I(n22), .ZN(n70) );
  INR2D4BWP30P140LVT U19 ( .A1(n41), .B1(n40), .ZN(n242) );
  INVD1BWP30P140LVT U20 ( .I(i_cmd[0]), .ZN(n4) );
  INR3D0BWP30P140LVT U21 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n4), .ZN(n8) );
  OR2D4BWP30P140LVT U22 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .Z(n16) );
  INVD1BWP30P140LVT U23 ( .I(rst), .ZN(n5) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n5), .A2(i_en), .Z(n9) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n26), .A2(n9), .Z(n7) );
  OR2D1BWP30P140LVT U26 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n39) );
  NR2D1BWP30P140LVT U27 ( .A1(n39), .A2(i_cmd[1]), .ZN(n6) );
  ND2OPTIBD1BWP30P140LVT U28 ( .A1(n7), .A2(n6), .ZN(n31) );
  INR2D1BWP30P140LVT U29 ( .A1(n8), .B1(n31), .ZN(n48) );
  INVD1BWP30P140LVT U30 ( .I(n9), .ZN(n23) );
  NR4D1BWP30P140LVT U31 ( .A1(i_cmd[3]), .A2(i_cmd[0]), .A3(i_cmd[4]), .A4(n23), .ZN(n10) );
  INVD2BWP30P140LVT U32 ( .I(n10), .ZN(n11) );
  NR2D1BWP30P140LVT U33 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n13) );
  CKAN2D1BWP30P140LVT U34 ( .A1(i_cmd[6]), .A2(i_valid[6]), .Z(n12) );
  ND3D2BWP30P140LVT U35 ( .A1(n19), .A2(n13), .A3(n12), .ZN(n14) );
  ND2D1BWP30P140LVT U36 ( .A1(i_cmd[5]), .A2(i_valid[5]), .ZN(n15) );
  NR2D1BWP30P140LVT U37 ( .A1(n16), .A2(n15), .ZN(n17) );
  INVD1BWP30P140LVT U38 ( .I(i_cmd[7]), .ZN(n18) );
  INR4D0BWP30P140LVT U39 ( .A1(i_valid[7]), .B1(i_cmd[6]), .B2(i_cmd[5]), .B3(
        n18), .ZN(n21) );
  INVD1BWP30P140LVT U40 ( .I(n19), .ZN(n20) );
  INR2D1BWP30P140LVT U41 ( .A1(n21), .B1(n20), .ZN(n22) );
  INVD2BWP30P140LVT U42 ( .I(n70), .ZN(n274) );
  NR4D0BWP30P140LVT U43 ( .A1(n48), .A2(n259), .A3(n1), .A4(n274), .ZN(n44) );
  INVD1BWP30P140LVT U44 ( .I(i_cmd[4]), .ZN(n25) );
  NR2D1BWP30P140LVT U45 ( .A1(i_cmd[0]), .A2(n23), .ZN(n24) );
  ND3OPTPAD2BWP30P140LVT U46 ( .A1(n26), .A2(n25), .A3(n24), .ZN(n40) );
  ND2D1BWP30P140LVT U47 ( .A1(i_cmd[3]), .A2(i_valid[3]), .ZN(n27) );
  OR2D1BWP30P140LVT U48 ( .A1(n28), .A2(n27), .Z(n29) );
  ND2D1BWP30P140LVT U49 ( .A1(i_cmd[4]), .A2(i_valid[4]), .ZN(n30) );
  NR2D1BWP30P140LVT U50 ( .A1(n30), .A2(i_cmd[0]), .ZN(n32) );
  INR2D1BWP30P140LVT U51 ( .A1(n32), .B1(n31), .ZN(n33) );
  INVD2BWP30P140LVT U52 ( .I(n33), .ZN(n61) );
  NR2D1BWP30P140LVT U53 ( .A1(n3), .A2(n268), .ZN(n43) );
  INVD1BWP30P140LVT U54 ( .I(i_cmd[2]), .ZN(n36) );
  OR2D1BWP30P140LVT U55 ( .A1(i_cmd[3]), .A2(i_cmd[1]), .Z(n35) );
  INVD1BWP30P140LVT U56 ( .I(i_valid[2]), .ZN(n34) );
  NR3D0P7BWP30P140LVT U57 ( .A1(n36), .A2(n35), .A3(n34), .ZN(n37) );
  INR2D4BWP30P140LVT U58 ( .A1(n37), .B1(n40), .ZN(n243) );
  ND2D1BWP30P140LVT U59 ( .A1(i_cmd[1]), .A2(i_valid[1]), .ZN(n38) );
  NR2D1BWP30P140LVT U60 ( .A1(n39), .A2(n38), .ZN(n41) );
  INVD1BWP30P140LVT U61 ( .I(n242), .ZN(n42) );
  ND4D1BWP30P140LVT U62 ( .A1(n44), .A2(n43), .A3(n2), .A4(n42), .ZN(N402) );
  AOI22D1BWP30P140LVT U63 ( .A1(n243), .A2(i_data_bus[95]), .B1(n242), .B2(
        i_data_bus[63]), .ZN(n52) );
  AOI22D1BWP30P140LVT U64 ( .A1(n3), .A2(i_data_bus[127]), .B1(n268), .B2(
        i_data_bus[159]), .ZN(n51) );
  INVD1BWP30P140LVT U65 ( .I(i_data_bus[223]), .ZN(n46) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[191]), .ZN(n45) );
  OAI22D1BWP30P140LVT U67 ( .A1(n137), .A2(n46), .B1(n105), .B2(n45), .ZN(n47)
         );
  AOI21D1BWP30P140LVT U68 ( .A1(n274), .A2(i_data_bus[255]), .B(n47), .ZN(n50)
         );
  INVD2BWP30P140LVT U69 ( .I(n56), .ZN(n275) );
  ND2D1BWP30P140LVT U70 ( .A1(n275), .A2(i_data_bus[31]), .ZN(n49) );
  ND4D1BWP30P140LVT U71 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(N400) );
  AOI22D1BWP30P140LVT U72 ( .A1(n243), .A2(i_data_bus[94]), .B1(n242), .B2(
        i_data_bus[62]), .ZN(n60) );
  AOI22D1BWP30P140LVT U73 ( .A1(n3), .A2(i_data_bus[126]), .B1(n268), .B2(
        i_data_bus[158]), .ZN(n59) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[222]), .ZN(n54) );
  INVD1BWP30P140LVT U75 ( .I(i_data_bus[190]), .ZN(n53) );
  OAI22D1BWP30P140LVT U76 ( .A1(n137), .A2(n54), .B1(n105), .B2(n53), .ZN(n55)
         );
  AOI21D1BWP30P140LVT U77 ( .A1(n262), .A2(i_data_bus[254]), .B(n55), .ZN(n58)
         );
  INVD2BWP30P140LVT U78 ( .I(n56), .ZN(n247) );
  ND2D1BWP30P140LVT U79 ( .A1(n247), .A2(i_data_bus[30]), .ZN(n57) );
  ND4D1BWP30P140LVT U80 ( .A1(n60), .A2(n59), .A3(n58), .A4(n57), .ZN(N399) );
  AOI22D1BWP30P140LVT U81 ( .A1(n243), .A2(i_data_bus[71]), .B1(n242), .B2(
        i_data_bus[39]), .ZN(n69) );
  INVD2BWP30P140LVT U82 ( .I(n61), .ZN(n244) );
  AOI22D1BWP30P140LVT U83 ( .A1(n3), .A2(i_data_bus[103]), .B1(n244), .B2(
        i_data_bus[135]), .ZN(n68) );
  INVD1BWP30P140LVT U84 ( .I(n105), .ZN(n62) );
  INVD2BWP30P140LVT U85 ( .I(n62), .ZN(n270) );
  INVD1BWP30P140LVT U86 ( .I(i_data_bus[167]), .ZN(n64) );
  INVD1BWP30P140LVT U87 ( .I(i_data_bus[199]), .ZN(n63) );
  OAI22D1BWP30P140LVT U88 ( .A1(n270), .A2(n64), .B1(n137), .B2(n63), .ZN(n65)
         );
  AOI21D1BWP30P140LVT U89 ( .A1(n274), .A2(i_data_bus[231]), .B(n65), .ZN(n67)
         );
  ND2D1BWP30P140LVT U90 ( .A1(n247), .A2(i_data_bus[7]), .ZN(n66) );
  ND4D1BWP30P140LVT U91 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(N376) );
  AOI22D1BWP30P140LVT U92 ( .A1(n243), .A2(i_data_bus[72]), .B1(n242), .B2(
        i_data_bus[40]), .ZN(n76) );
  AOI22D1BWP30P140LVT U93 ( .A1(n3), .A2(i_data_bus[104]), .B1(n244), .B2(
        i_data_bus[136]), .ZN(n75) );
  INVD2BWP30P140LVT U94 ( .I(n70), .ZN(n262) );
  INVD1BWP30P140LVT U95 ( .I(i_data_bus[168]), .ZN(n71) );
  MOAI22D1BWP30P140LVT U96 ( .A1(n270), .A2(n71), .B1(n259), .B2(
        i_data_bus[200]), .ZN(n72) );
  AOI21D1BWP30P140LVT U97 ( .A1(n262), .A2(i_data_bus[232]), .B(n72), .ZN(n74)
         );
  ND2D1BWP30P140LVT U98 ( .A1(n247), .A2(i_data_bus[8]), .ZN(n73) );
  ND4D1BWP30P140LVT U99 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(N377) );
  AOI22D1BWP30P140LVT U100 ( .A1(n243), .A2(i_data_bus[76]), .B1(n242), .B2(
        i_data_bus[44]), .ZN(n83) );
  AOI22D1BWP30P140LVT U101 ( .A1(n3), .A2(i_data_bus[108]), .B1(n244), .B2(
        i_data_bus[140]), .ZN(n82) );
  INVD2BWP30P140LVT U102 ( .I(n259), .ZN(n272) );
  INVD1BWP30P140LVT U103 ( .I(i_data_bus[204]), .ZN(n78) );
  INVD1BWP30P140LVT U104 ( .I(i_data_bus[172]), .ZN(n77) );
  OAI22D1BWP30P140LVT U105 ( .A1(n272), .A2(n78), .B1(n270), .B2(n77), .ZN(n79) );
  AOI21D1BWP30P140LVT U106 ( .A1(n274), .A2(i_data_bus[236]), .B(n79), .ZN(n81) );
  ND2D1BWP30P140LVT U107 ( .A1(n247), .A2(i_data_bus[12]), .ZN(n80) );
  ND4D1BWP30P140LVT U108 ( .A1(n83), .A2(n82), .A3(n81), .A4(n80), .ZN(N381)
         );
  AOI22D1BWP30P140LVT U109 ( .A1(n243), .A2(i_data_bus[75]), .B1(n242), .B2(
        i_data_bus[43]), .ZN(n90) );
  AOI22D1BWP30P140LVT U110 ( .A1(n3), .A2(i_data_bus[107]), .B1(n244), .B2(
        i_data_bus[139]), .ZN(n89) );
  INVD1BWP30P140LVT U111 ( .I(i_data_bus[203]), .ZN(n85) );
  INVD1BWP30P140LVT U112 ( .I(i_data_bus[171]), .ZN(n84) );
  OAI22D1BWP30P140LVT U113 ( .A1(n272), .A2(n85), .B1(n270), .B2(n84), .ZN(n86) );
  AOI21D1BWP30P140LVT U114 ( .A1(n274), .A2(i_data_bus[235]), .B(n86), .ZN(n88) );
  ND2D1BWP30P140LVT U115 ( .A1(n247), .A2(i_data_bus[11]), .ZN(n87) );
  ND4D1BWP30P140LVT U116 ( .A1(n90), .A2(n89), .A3(n88), .A4(n87), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U117 ( .A1(n243), .A2(i_data_bus[74]), .B1(n242), .B2(
        i_data_bus[42]), .ZN(n97) );
  AOI22D1BWP30P140LVT U118 ( .A1(n3), .A2(i_data_bus[106]), .B1(n244), .B2(
        i_data_bus[138]), .ZN(n96) );
  INVD1BWP30P140LVT U119 ( .I(i_data_bus[202]), .ZN(n92) );
  INVD1BWP30P140LVT U120 ( .I(i_data_bus[170]), .ZN(n91) );
  OAI22D1BWP30P140LVT U121 ( .A1(n272), .A2(n92), .B1(n270), .B2(n91), .ZN(n93) );
  AOI21D1BWP30P140LVT U122 ( .A1(n274), .A2(i_data_bus[234]), .B(n93), .ZN(n95) );
  ND2D1BWP30P140LVT U123 ( .A1(n247), .A2(i_data_bus[10]), .ZN(n94) );
  ND4D1BWP30P140LVT U124 ( .A1(n97), .A2(n96), .A3(n95), .A4(n94), .ZN(N379)
         );
  AOI22D1BWP30P140LVT U125 ( .A1(n243), .A2(i_data_bus[73]), .B1(n242), .B2(
        i_data_bus[41]), .ZN(n104) );
  AOI22D1BWP30P140LVT U126 ( .A1(n3), .A2(i_data_bus[105]), .B1(n244), .B2(
        i_data_bus[137]), .ZN(n103) );
  INVD1BWP30P140LVT U127 ( .I(i_data_bus[201]), .ZN(n99) );
  INVD1BWP30P140LVT U128 ( .I(i_data_bus[169]), .ZN(n98) );
  OAI22D1BWP30P140LVT U129 ( .A1(n272), .A2(n99), .B1(n270), .B2(n98), .ZN(
        n100) );
  AOI21D1BWP30P140LVT U130 ( .A1(n274), .A2(i_data_bus[233]), .B(n100), .ZN(
        n102) );
  ND2D1BWP30P140LVT U131 ( .A1(n247), .A2(i_data_bus[9]), .ZN(n101) );
  ND4D1BWP30P140LVT U132 ( .A1(n104), .A2(n103), .A3(n102), .A4(n101), .ZN(
        N378) );
  AOI22D1BWP30P140LVT U133 ( .A1(n243), .A2(i_data_bus[93]), .B1(n242), .B2(
        i_data_bus[61]), .ZN(n112) );
  AOI22D1BWP30P140LVT U134 ( .A1(n3), .A2(i_data_bus[125]), .B1(n268), .B2(
        i_data_bus[157]), .ZN(n111) );
  INVD1BWP30P140LVT U135 ( .I(i_data_bus[221]), .ZN(n107) );
  INVD2BWP30P140LVT U136 ( .I(n1), .ZN(n253) );
  INVD1BWP30P140LVT U137 ( .I(i_data_bus[189]), .ZN(n106) );
  OAI22D1BWP30P140LVT U138 ( .A1(n137), .A2(n107), .B1(n253), .B2(n106), .ZN(
        n108) );
  AOI21D1BWP30P140LVT U139 ( .A1(n262), .A2(i_data_bus[253]), .B(n108), .ZN(
        n110) );
  ND2D1BWP30P140LVT U140 ( .A1(n247), .A2(i_data_bus[29]), .ZN(n109) );
  ND4D1BWP30P140LVT U141 ( .A1(n112), .A2(n111), .A3(n110), .A4(n109), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U142 ( .A1(n243), .A2(i_data_bus[92]), .B1(n242), .B2(
        i_data_bus[60]), .ZN(n119) );
  AOI22D1BWP30P140LVT U143 ( .A1(n3), .A2(i_data_bus[124]), .B1(n268), .B2(
        i_data_bus[156]), .ZN(n118) );
  INVD1BWP30P140LVT U144 ( .I(i_data_bus[220]), .ZN(n114) );
  INVD1BWP30P140LVT U145 ( .I(i_data_bus[188]), .ZN(n113) );
  OAI22D1BWP30P140LVT U146 ( .A1(n137), .A2(n114), .B1(n253), .B2(n113), .ZN(
        n115) );
  AOI21D1BWP30P140LVT U147 ( .A1(n262), .A2(i_data_bus[252]), .B(n115), .ZN(
        n117) );
  ND2D1BWP30P140LVT U148 ( .A1(n275), .A2(i_data_bus[28]), .ZN(n116) );
  ND4D1BWP30P140LVT U149 ( .A1(n119), .A2(n118), .A3(n117), .A4(n116), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U150 ( .A1(n243), .A2(i_data_bus[91]), .B1(n242), .B2(
        i_data_bus[59]), .ZN(n126) );
  AOI22D1BWP30P140LVT U151 ( .A1(n3), .A2(i_data_bus[123]), .B1(n268), .B2(
        i_data_bus[155]), .ZN(n125) );
  INVD1BWP30P140LVT U152 ( .I(i_data_bus[219]), .ZN(n121) );
  INVD1BWP30P140LVT U153 ( .I(i_data_bus[187]), .ZN(n120) );
  OAI22D1BWP30P140LVT U154 ( .A1(n137), .A2(n121), .B1(n253), .B2(n120), .ZN(
        n122) );
  AOI21D1BWP30P140LVT U155 ( .A1(n262), .A2(i_data_bus[251]), .B(n122), .ZN(
        n124) );
  ND2D1BWP30P140LVT U156 ( .A1(n247), .A2(i_data_bus[27]), .ZN(n123) );
  ND4D1BWP30P140LVT U157 ( .A1(n126), .A2(n125), .A3(n124), .A4(n123), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U158 ( .A1(n243), .A2(i_data_bus[90]), .B1(n242), .B2(
        i_data_bus[58]), .ZN(n133) );
  AOI22D1BWP30P140LVT U159 ( .A1(n3), .A2(i_data_bus[122]), .B1(n268), .B2(
        i_data_bus[154]), .ZN(n132) );
  INVD1BWP30P140LVT U160 ( .I(i_data_bus[218]), .ZN(n128) );
  INVD1BWP30P140LVT U161 ( .I(i_data_bus[186]), .ZN(n127) );
  OAI22D1BWP30P140LVT U162 ( .A1(n137), .A2(n128), .B1(n253), .B2(n127), .ZN(
        n129) );
  AOI21D1BWP30P140LVT U163 ( .A1(n262), .A2(i_data_bus[250]), .B(n129), .ZN(
        n131) );
  ND2D1BWP30P140LVT U164 ( .A1(n275), .A2(i_data_bus[26]), .ZN(n130) );
  ND4D1BWP30P140LVT U165 ( .A1(n133), .A2(n132), .A3(n131), .A4(n130), .ZN(
        N395) );
  INVD2BWP30P140LVT U166 ( .I(n2), .ZN(n267) );
  AOI22D1BWP30P140LVT U167 ( .A1(n267), .A2(i_data_bus[89]), .B1(n242), .B2(
        i_data_bus[57]), .ZN(n142) );
  AOI22D1BWP30P140LVT U168 ( .A1(n3), .A2(i_data_bus[121]), .B1(n268), .B2(
        i_data_bus[153]), .ZN(n141) );
  INVD1BWP30P140LVT U169 ( .I(i_data_bus[217]), .ZN(n136) );
  INVD1BWP30P140LVT U170 ( .I(i_data_bus[185]), .ZN(n135) );
  OAI22D1BWP30P140LVT U171 ( .A1(n137), .A2(n136), .B1(n253), .B2(n135), .ZN(
        n138) );
  AOI21D1BWP30P140LVT U172 ( .A1(n262), .A2(i_data_bus[249]), .B(n138), .ZN(
        n140) );
  ND2D1BWP30P140LVT U173 ( .A1(n275), .A2(i_data_bus[25]), .ZN(n139) );
  ND4D1BWP30P140LVT U174 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U175 ( .A1(n267), .A2(i_data_bus[88]), .B1(n242), .B2(
        i_data_bus[56]), .ZN(n149) );
  AOI22D1BWP30P140LVT U176 ( .A1(n3), .A2(i_data_bus[120]), .B1(n268), .B2(
        i_data_bus[152]), .ZN(n148) );
  INVD1BWP30P140LVT U177 ( .I(i_data_bus[216]), .ZN(n144) );
  INVD1BWP30P140LVT U178 ( .I(i_data_bus[184]), .ZN(n143) );
  OAI22D1BWP30P140LVT U179 ( .A1(n272), .A2(n144), .B1(n253), .B2(n143), .ZN(
        n145) );
  AOI21D1BWP30P140LVT U180 ( .A1(n262), .A2(i_data_bus[248]), .B(n145), .ZN(
        n147) );
  ND2D1BWP30P140LVT U181 ( .A1(n275), .A2(i_data_bus[24]), .ZN(n146) );
  ND4D1BWP30P140LVT U182 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U183 ( .A1(n267), .A2(i_data_bus[87]), .B1(n242), .B2(
        i_data_bus[55]), .ZN(n156) );
  AOI22D1BWP30P140LVT U184 ( .A1(n3), .A2(i_data_bus[119]), .B1(n268), .B2(
        i_data_bus[151]), .ZN(n155) );
  INVD1BWP30P140LVT U185 ( .I(i_data_bus[215]), .ZN(n151) );
  INVD1BWP30P140LVT U186 ( .I(i_data_bus[183]), .ZN(n150) );
  OAI22D1BWP30P140LVT U187 ( .A1(n272), .A2(n151), .B1(n253), .B2(n150), .ZN(
        n152) );
  AOI21D1BWP30P140LVT U188 ( .A1(n262), .A2(i_data_bus[247]), .B(n152), .ZN(
        n154) );
  ND2D1BWP30P140LVT U189 ( .A1(n275), .A2(i_data_bus[23]), .ZN(n153) );
  ND4D1BWP30P140LVT U190 ( .A1(n156), .A2(n155), .A3(n154), .A4(n153), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U191 ( .A1(n267), .A2(i_data_bus[86]), .B1(n242), .B2(
        i_data_bus[54]), .ZN(n163) );
  AOI22D1BWP30P140LVT U192 ( .A1(n3), .A2(i_data_bus[118]), .B1(n268), .B2(
        i_data_bus[150]), .ZN(n162) );
  INVD1BWP30P140LVT U193 ( .I(i_data_bus[214]), .ZN(n158) );
  INVD1BWP30P140LVT U194 ( .I(i_data_bus[182]), .ZN(n157) );
  OAI22D1BWP30P140LVT U195 ( .A1(n272), .A2(n158), .B1(n253), .B2(n157), .ZN(
        n159) );
  AOI21D1BWP30P140LVT U196 ( .A1(n262), .A2(i_data_bus[246]), .B(n159), .ZN(
        n161) );
  ND2D1BWP30P140LVT U197 ( .A1(n275), .A2(i_data_bus[22]), .ZN(n160) );
  ND4D1BWP30P140LVT U198 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U199 ( .A1(n267), .A2(i_data_bus[85]), .B1(n242), .B2(
        i_data_bus[53]), .ZN(n170) );
  AOI22D1BWP30P140LVT U200 ( .A1(n3), .A2(i_data_bus[117]), .B1(n268), .B2(
        i_data_bus[149]), .ZN(n169) );
  INVD1BWP30P140LVT U201 ( .I(i_data_bus[213]), .ZN(n165) );
  INVD1BWP30P140LVT U202 ( .I(i_data_bus[181]), .ZN(n164) );
  OAI22D1BWP30P140LVT U203 ( .A1(n272), .A2(n165), .B1(n253), .B2(n164), .ZN(
        n166) );
  AOI21D1BWP30P140LVT U204 ( .A1(n262), .A2(i_data_bus[245]), .B(n166), .ZN(
        n168) );
  ND2D1BWP30P140LVT U205 ( .A1(n275), .A2(i_data_bus[21]), .ZN(n167) );
  ND4D1BWP30P140LVT U206 ( .A1(n170), .A2(n169), .A3(n168), .A4(n167), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U207 ( .A1(n267), .A2(i_data_bus[84]), .B1(n242), .B2(
        i_data_bus[52]), .ZN(n177) );
  AOI22D1BWP30P140LVT U208 ( .A1(n3), .A2(i_data_bus[116]), .B1(n268), .B2(
        i_data_bus[148]), .ZN(n176) );
  INVD1BWP30P140LVT U209 ( .I(i_data_bus[212]), .ZN(n172) );
  INVD1BWP30P140LVT U210 ( .I(i_data_bus[180]), .ZN(n171) );
  OAI22D1BWP30P140LVT U211 ( .A1(n272), .A2(n172), .B1(n253), .B2(n171), .ZN(
        n173) );
  AOI21D1BWP30P140LVT U212 ( .A1(n262), .A2(i_data_bus[244]), .B(n173), .ZN(
        n175) );
  ND2D1BWP30P140LVT U213 ( .A1(n275), .A2(i_data_bus[20]), .ZN(n174) );
  ND4D1BWP30P140LVT U214 ( .A1(n177), .A2(n176), .A3(n175), .A4(n174), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U215 ( .A1(n267), .A2(i_data_bus[83]), .B1(n242), .B2(
        i_data_bus[51]), .ZN(n183) );
  AOI22D1BWP30P140LVT U216 ( .A1(n3), .A2(i_data_bus[115]), .B1(n268), .B2(
        i_data_bus[147]), .ZN(n182) );
  INVD1BWP30P140LVT U217 ( .I(i_data_bus[179]), .ZN(n178) );
  MOAI22D1BWP30P140LVT U218 ( .A1(n253), .A2(n178), .B1(n259), .B2(
        i_data_bus[211]), .ZN(n179) );
  AOI21D1BWP30P140LVT U219 ( .A1(n262), .A2(i_data_bus[243]), .B(n179), .ZN(
        n181) );
  ND2D1BWP30P140LVT U220 ( .A1(n275), .A2(i_data_bus[19]), .ZN(n180) );
  ND4D1BWP30P140LVT U221 ( .A1(n183), .A2(n182), .A3(n181), .A4(n180), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U222 ( .A1(n267), .A2(i_data_bus[82]), .B1(n242), .B2(
        i_data_bus[50]), .ZN(n189) );
  AOI22D1BWP30P140LVT U223 ( .A1(n3), .A2(i_data_bus[114]), .B1(n268), .B2(
        i_data_bus[146]), .ZN(n188) );
  INVD1BWP30P140LVT U224 ( .I(i_data_bus[178]), .ZN(n184) );
  MOAI22D1BWP30P140LVT U225 ( .A1(n253), .A2(n184), .B1(n259), .B2(
        i_data_bus[210]), .ZN(n185) );
  AOI21D1BWP30P140LVT U226 ( .A1(n262), .A2(i_data_bus[242]), .B(n185), .ZN(
        n187) );
  ND2D1BWP30P140LVT U227 ( .A1(n275), .A2(i_data_bus[18]), .ZN(n186) );
  ND4D1BWP30P140LVT U228 ( .A1(n189), .A2(n188), .A3(n187), .A4(n186), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U229 ( .A1(n267), .A2(i_data_bus[81]), .B1(n242), .B2(
        i_data_bus[49]), .ZN(n195) );
  AOI22D1BWP30P140LVT U230 ( .A1(n3), .A2(i_data_bus[113]), .B1(n268), .B2(
        i_data_bus[145]), .ZN(n194) );
  INVD1BWP30P140LVT U231 ( .I(i_data_bus[177]), .ZN(n190) );
  MOAI22D1BWP30P140LVT U232 ( .A1(n253), .A2(n190), .B1(n259), .B2(
        i_data_bus[209]), .ZN(n191) );
  AOI21D1BWP30P140LVT U233 ( .A1(n262), .A2(i_data_bus[241]), .B(n191), .ZN(
        n193) );
  ND2D1BWP30P140LVT U234 ( .A1(n275), .A2(i_data_bus[17]), .ZN(n192) );
  ND4D1BWP30P140LVT U235 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U236 ( .A1(n267), .A2(i_data_bus[80]), .B1(n242), .B2(
        i_data_bus[48]), .ZN(n201) );
  AOI22D1BWP30P140LVT U237 ( .A1(n3), .A2(i_data_bus[112]), .B1(n268), .B2(
        i_data_bus[144]), .ZN(n200) );
  INVD1BWP30P140LVT U238 ( .I(i_data_bus[176]), .ZN(n196) );
  MOAI22D1BWP30P140LVT U239 ( .A1(n253), .A2(n196), .B1(n259), .B2(
        i_data_bus[208]), .ZN(n197) );
  AOI21D1BWP30P140LVT U240 ( .A1(n262), .A2(i_data_bus[240]), .B(n197), .ZN(
        n199) );
  ND2D1BWP30P140LVT U241 ( .A1(n275), .A2(i_data_bus[16]), .ZN(n198) );
  ND4D1BWP30P140LVT U242 ( .A1(n201), .A2(n200), .A3(n199), .A4(n198), .ZN(
        N385) );
  AOI22D1BWP30P140LVT U243 ( .A1(n243), .A2(i_data_bus[70]), .B1(n242), .B2(
        i_data_bus[38]), .ZN(n208) );
  AOI22D1BWP30P140LVT U244 ( .A1(n3), .A2(i_data_bus[102]), .B1(n244), .B2(
        i_data_bus[134]), .ZN(n207) );
  INVD1BWP30P140LVT U245 ( .I(i_data_bus[198]), .ZN(n203) );
  INVD1BWP30P140LVT U246 ( .I(i_data_bus[166]), .ZN(n202) );
  OAI22D1BWP30P140LVT U247 ( .A1(n272), .A2(n203), .B1(n270), .B2(n202), .ZN(
        n204) );
  AOI21D1BWP30P140LVT U248 ( .A1(n274), .A2(i_data_bus[230]), .B(n204), .ZN(
        n206) );
  ND2D1BWP30P140LVT U249 ( .A1(n247), .A2(i_data_bus[6]), .ZN(n205) );
  ND4D1BWP30P140LVT U250 ( .A1(n208), .A2(n207), .A3(n206), .A4(n205), .ZN(
        N375) );
  AOI22D1BWP30P140LVT U251 ( .A1(n243), .A2(i_data_bus[69]), .B1(n242), .B2(
        i_data_bus[37]), .ZN(n215) );
  AOI22D1BWP30P140LVT U252 ( .A1(n3), .A2(i_data_bus[101]), .B1(n244), .B2(
        i_data_bus[133]), .ZN(n214) );
  INVD1BWP30P140LVT U253 ( .I(i_data_bus[197]), .ZN(n210) );
  INVD1BWP30P140LVT U254 ( .I(i_data_bus[165]), .ZN(n209) );
  OAI22D1BWP30P140LVT U255 ( .A1(n272), .A2(n210), .B1(n270), .B2(n209), .ZN(
        n211) );
  AOI21D1BWP30P140LVT U256 ( .A1(n274), .A2(i_data_bus[229]), .B(n211), .ZN(
        n213) );
  ND2D1BWP30P140LVT U257 ( .A1(n247), .A2(i_data_bus[5]), .ZN(n212) );
  ND4D1BWP30P140LVT U258 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .ZN(
        N374) );
  AOI22D1BWP30P140LVT U259 ( .A1(n243), .A2(i_data_bus[64]), .B1(n242), .B2(
        i_data_bus[32]), .ZN(n221) );
  AOI22D1BWP30P140LVT U260 ( .A1(n3), .A2(i_data_bus[96]), .B1(n244), .B2(
        i_data_bus[128]), .ZN(n220) );
  INR2D1BWP30P140LVT U261 ( .A1(i_data_bus[192]), .B1(n272), .ZN(n217) );
  INR2D1BWP30P140LVT U262 ( .A1(i_data_bus[160]), .B1(n270), .ZN(n216) );
  AOI211D1BWP30P140LVT U263 ( .A1(i_data_bus[224]), .A2(n274), .B(n217), .C(
        n216), .ZN(n219) );
  ND2D1BWP30P140LVT U264 ( .A1(n247), .A2(i_data_bus[0]), .ZN(n218) );
  ND4D1BWP30P140LVT U265 ( .A1(n221), .A2(n220), .A3(n219), .A4(n218), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U266 ( .A1(n243), .A2(i_data_bus[68]), .B1(n242), .B2(
        i_data_bus[36]), .ZN(n228) );
  AOI22D1BWP30P140LVT U267 ( .A1(n3), .A2(i_data_bus[100]), .B1(n244), .B2(
        i_data_bus[132]), .ZN(n227) );
  INVD1BWP30P140LVT U268 ( .I(i_data_bus[196]), .ZN(n223) );
  INVD1BWP30P140LVT U269 ( .I(i_data_bus[164]), .ZN(n222) );
  OAI22D1BWP30P140LVT U270 ( .A1(n272), .A2(n223), .B1(n270), .B2(n222), .ZN(
        n224) );
  ND2D1BWP30P140LVT U271 ( .A1(n247), .A2(i_data_bus[4]), .ZN(n225) );
  ND4D1BWP30P140LVT U272 ( .A1(n228), .A2(n227), .A3(n226), .A4(n225), .ZN(
        N373) );
  AOI22D1BWP30P140LVT U273 ( .A1(n243), .A2(i_data_bus[67]), .B1(n242), .B2(
        i_data_bus[35]), .ZN(n235) );
  AOI22D1BWP30P140LVT U274 ( .A1(n3), .A2(i_data_bus[99]), .B1(n244), .B2(
        i_data_bus[131]), .ZN(n234) );
  INVD1BWP30P140LVT U275 ( .I(i_data_bus[195]), .ZN(n230) );
  INVD1BWP30P140LVT U276 ( .I(i_data_bus[163]), .ZN(n229) );
  OAI22D1BWP30P140LVT U277 ( .A1(n272), .A2(n230), .B1(n270), .B2(n229), .ZN(
        n231) );
  ND2D1BWP30P140LVT U278 ( .A1(n247), .A2(i_data_bus[3]), .ZN(n232) );
  ND4D1BWP30P140LVT U279 ( .A1(n235), .A2(n234), .A3(n233), .A4(n232), .ZN(
        N372) );
  AOI22D1BWP30P140LVT U280 ( .A1(n243), .A2(i_data_bus[66]), .B1(n242), .B2(
        i_data_bus[34]), .ZN(n241) );
  AOI22D1BWP30P140LVT U281 ( .A1(n3), .A2(i_data_bus[98]), .B1(n244), .B2(
        i_data_bus[130]), .ZN(n240) );
  INVD1BWP30P140LVT U282 ( .I(i_data_bus[162]), .ZN(n236) );
  MOAI22D1BWP30P140LVT U283 ( .A1(n270), .A2(n236), .B1(n259), .B2(
        i_data_bus[194]), .ZN(n237) );
  AOI21D1BWP30P140LVT U284 ( .A1(n274), .A2(i_data_bus[226]), .B(n237), .ZN(
        n239) );
  ND2D1BWP30P140LVT U285 ( .A1(n247), .A2(i_data_bus[2]), .ZN(n238) );
  ND4D1BWP30P140LVT U286 ( .A1(n241), .A2(n240), .A3(n239), .A4(n238), .ZN(
        N371) );
  AOI22D1BWP30P140LVT U287 ( .A1(n243), .A2(i_data_bus[65]), .B1(n242), .B2(
        i_data_bus[33]), .ZN(n251) );
  AOI22D1BWP30P140LVT U288 ( .A1(n3), .A2(i_data_bus[97]), .B1(n244), .B2(
        i_data_bus[129]), .ZN(n250) );
  INVD1BWP30P140LVT U289 ( .I(i_data_bus[161]), .ZN(n245) );
  MOAI22D1BWP30P140LVT U290 ( .A1(n270), .A2(n245), .B1(n259), .B2(
        i_data_bus[193]), .ZN(n246) );
  AOI21D1BWP30P140LVT U291 ( .A1(n274), .A2(i_data_bus[225]), .B(n246), .ZN(
        n249) );
  ND2D1BWP30P140LVT U292 ( .A1(n247), .A2(i_data_bus[1]), .ZN(n248) );
  ND4D1BWP30P140LVT U293 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U294 ( .A1(n267), .A2(i_data_bus[79]), .B1(n242), .B2(
        i_data_bus[47]), .ZN(n258) );
  AOI22D1BWP30P140LVT U295 ( .A1(n3), .A2(i_data_bus[111]), .B1(n268), .B2(
        i_data_bus[143]), .ZN(n257) );
  INVD1BWP30P140LVT U296 ( .I(i_data_bus[175]), .ZN(n252) );
  MOAI22D1BWP30P140LVT U297 ( .A1(n253), .A2(n252), .B1(n259), .B2(
        i_data_bus[207]), .ZN(n254) );
  AOI21D1BWP30P140LVT U298 ( .A1(n262), .A2(i_data_bus[239]), .B(n254), .ZN(
        n256) );
  ND2D1BWP30P140LVT U299 ( .A1(n275), .A2(i_data_bus[15]), .ZN(n255) );
  ND4D1BWP30P140LVT U300 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U301 ( .A1(n267), .A2(i_data_bus[78]), .B1(n242), .B2(
        i_data_bus[46]), .ZN(n266) );
  AOI22D1BWP30P140LVT U302 ( .A1(n3), .A2(i_data_bus[110]), .B1(n268), .B2(
        i_data_bus[142]), .ZN(n265) );
  INVD1BWP30P140LVT U303 ( .I(i_data_bus[174]), .ZN(n260) );
  MOAI22D1BWP30P140LVT U304 ( .A1(n270), .A2(n260), .B1(n259), .B2(
        i_data_bus[206]), .ZN(n261) );
  AOI21D1BWP30P140LVT U305 ( .A1(n262), .A2(i_data_bus[238]), .B(n261), .ZN(
        n264) );
  ND2D1BWP30P140LVT U306 ( .A1(n275), .A2(i_data_bus[14]), .ZN(n263) );
  ND4D1BWP30P140LVT U307 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U308 ( .A1(n267), .A2(i_data_bus[77]), .B1(n242), .B2(
        i_data_bus[45]), .ZN(n279) );
  AOI22D1BWP30P140LVT U309 ( .A1(n3), .A2(i_data_bus[109]), .B1(n268), .B2(
        i_data_bus[141]), .ZN(n278) );
  INVD1BWP30P140LVT U310 ( .I(i_data_bus[205]), .ZN(n271) );
  INVD1BWP30P140LVT U311 ( .I(i_data_bus[173]), .ZN(n269) );
  OAI22D1BWP30P140LVT U312 ( .A1(n272), .A2(n271), .B1(n270), .B2(n269), .ZN(
        n273) );
  ND2D1BWP30P140LVT U313 ( .A1(n275), .A2(i_data_bus[13]), .ZN(n276) );
  ND4D1BWP30P140LVT U314 ( .A1(n279), .A2(n278), .A3(n277), .A4(n276), .ZN(
        N382) );
endmodule


module crossbar_8_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA8_1 ( clk, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [63:0] i_cmd;
  input clk, rst, i_en;

  wire   [63:0] o_inner_cmd_wire;
  wire   [255:0] bottom_half_0__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_0__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_1__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_1__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_2__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_2__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_3__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_3__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_4__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_4__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_5__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_5__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_6__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_6__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_7__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_7__inner_valid_i_mux_tree_wire;

  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_8 top_half_0__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[0]), .i_data_bus(
        i_data_bus[31:0]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[0], 
        bottom_half_6__inner_valid_i_mux_tree_wire[0], 
        bottom_half_5__inner_valid_i_mux_tree_wire[0], 
        bottom_half_4__inner_valid_i_mux_tree_wire[0], 
        bottom_half_3__inner_valid_i_mux_tree_wire[0], 
        bottom_half_2__inner_valid_i_mux_tree_wire[0], 
        bottom_half_1__inner_valid_i_mux_tree_wire[0], 
        bottom_half_0__inner_valid_i_mux_tree_wire[0]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_6__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_5__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_4__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_3__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_2__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_1__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_0__inner_data_i_mux_tree_wire[31:0]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 top_half_1__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[1]), .i_data_bus(
        i_data_bus[63:32]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[1], 
        bottom_half_6__inner_valid_i_mux_tree_wire[1], 
        bottom_half_5__inner_valid_i_mux_tree_wire[1], 
        bottom_half_4__inner_valid_i_mux_tree_wire[1], 
        bottom_half_3__inner_valid_i_mux_tree_wire[1], 
        bottom_half_2__inner_valid_i_mux_tree_wire[1], 
        bottom_half_1__inner_valid_i_mux_tree_wire[1], 
        bottom_half_0__inner_valid_i_mux_tree_wire[1]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_6__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_5__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_4__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_3__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_2__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_1__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_0__inner_data_i_mux_tree_wire[63:32]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 top_half_2__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[2]), .i_data_bus(
        i_data_bus[95:64]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[2], 
        bottom_half_6__inner_valid_i_mux_tree_wire[2], 
        bottom_half_5__inner_valid_i_mux_tree_wire[2], 
        bottom_half_4__inner_valid_i_mux_tree_wire[2], 
        bottom_half_3__inner_valid_i_mux_tree_wire[2], 
        bottom_half_2__inner_valid_i_mux_tree_wire[2], 
        bottom_half_1__inner_valid_i_mux_tree_wire[2], 
        bottom_half_0__inner_valid_i_mux_tree_wire[2]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_6__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_5__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_4__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_3__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_2__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_1__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_0__inner_data_i_mux_tree_wire[95:64]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 top_half_3__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[3]), .i_data_bus(
        i_data_bus[127:96]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[3], 
        bottom_half_6__inner_valid_i_mux_tree_wire[3], 
        bottom_half_5__inner_valid_i_mux_tree_wire[3], 
        bottom_half_4__inner_valid_i_mux_tree_wire[3], 
        bottom_half_3__inner_valid_i_mux_tree_wire[3], 
        bottom_half_2__inner_valid_i_mux_tree_wire[3], 
        bottom_half_1__inner_valid_i_mux_tree_wire[3], 
        bottom_half_0__inner_valid_i_mux_tree_wire[3]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_6__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_5__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_4__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_3__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_2__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_1__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_0__inner_data_i_mux_tree_wire[127:96]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 top_half_4__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[4]), .i_data_bus(
        i_data_bus[159:128]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[4], 
        bottom_half_6__inner_valid_i_mux_tree_wire[4], 
        bottom_half_5__inner_valid_i_mux_tree_wire[4], 
        bottom_half_4__inner_valid_i_mux_tree_wire[4], 
        bottom_half_3__inner_valid_i_mux_tree_wire[4], 
        bottom_half_2__inner_valid_i_mux_tree_wire[4], 
        bottom_half_1__inner_valid_i_mux_tree_wire[4], 
        bottom_half_0__inner_valid_i_mux_tree_wire[4]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_6__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_5__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_4__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_3__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_2__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_1__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_0__inner_data_i_mux_tree_wire[159:128]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 top_half_5__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[5]), .i_data_bus(
        i_data_bus[191:160]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[5], 
        bottom_half_6__inner_valid_i_mux_tree_wire[5], 
        bottom_half_5__inner_valid_i_mux_tree_wire[5], 
        bottom_half_4__inner_valid_i_mux_tree_wire[5], 
        bottom_half_3__inner_valid_i_mux_tree_wire[5], 
        bottom_half_2__inner_valid_i_mux_tree_wire[5], 
        bottom_half_1__inner_valid_i_mux_tree_wire[5], 
        bottom_half_0__inner_valid_i_mux_tree_wire[5]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_6__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_5__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_4__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_3__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_2__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_1__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_0__inner_data_i_mux_tree_wire[191:160]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 top_half_6__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[6]), .i_data_bus(
        i_data_bus[223:192]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[6], 
        bottom_half_6__inner_valid_i_mux_tree_wire[6], 
        bottom_half_5__inner_valid_i_mux_tree_wire[6], 
        bottom_half_4__inner_valid_i_mux_tree_wire[6], 
        bottom_half_3__inner_valid_i_mux_tree_wire[6], 
        bottom_half_2__inner_valid_i_mux_tree_wire[6], 
        bottom_half_1__inner_valid_i_mux_tree_wire[6], 
        bottom_half_0__inner_valid_i_mux_tree_wire[6]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_6__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_5__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_4__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_3__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_2__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_1__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_0__inner_data_i_mux_tree_wire[223:192]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 top_half_7__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[7]), .i_data_bus(
        i_data_bus[255:224]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[7], 
        bottom_half_6__inner_valid_i_mux_tree_wire[7], 
        bottom_half_5__inner_valid_i_mux_tree_wire[7], 
        bottom_half_4__inner_valid_i_mux_tree_wire[7], 
        bottom_half_3__inner_valid_i_mux_tree_wire[7], 
        bottom_half_2__inner_valid_i_mux_tree_wire[7], 
        bottom_half_1__inner_valid_i_mux_tree_wire[7], 
        bottom_half_0__inner_valid_i_mux_tree_wire[7]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_6__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_5__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_4__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_3__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_2__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_1__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_0__inner_data_i_mux_tree_wire[255:224]}), .i_en(i_en) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_8 i_cmd_id_0__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[0]), .o_cmd_1(
        o_inner_cmd_wire[8]), .o_cmd_2(o_inner_cmd_wire[16]), .o_cmd_3(
        o_inner_cmd_wire[24]), .o_cmd_4(o_inner_cmd_wire[32]), .o_cmd_5(
        o_inner_cmd_wire[40]), .o_cmd_6(o_inner_cmd_wire[48]), .o_cmd_7(
        o_inner_cmd_wire[56]), .i_en(i_en), .i_cmd(i_cmd[7:0]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 i_cmd_id_1__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[1]), .o_cmd_1(
        o_inner_cmd_wire[9]), .o_cmd_2(o_inner_cmd_wire[17]), .o_cmd_3(
        o_inner_cmd_wire[25]), .o_cmd_4(o_inner_cmd_wire[33]), .o_cmd_5(
        o_inner_cmd_wire[41]), .o_cmd_6(o_inner_cmd_wire[49]), .o_cmd_7(
        o_inner_cmd_wire[57]), .i_en(i_en), .i_cmd(i_cmd[15:8]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 i_cmd_id_2__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[2]), .o_cmd_1(
        o_inner_cmd_wire[10]), .o_cmd_2(o_inner_cmd_wire[18]), .o_cmd_3(
        o_inner_cmd_wire[26]), .o_cmd_4(o_inner_cmd_wire[34]), .o_cmd_5(
        o_inner_cmd_wire[42]), .o_cmd_6(o_inner_cmd_wire[50]), .o_cmd_7(
        o_inner_cmd_wire[58]), .i_en(i_en), .i_cmd(i_cmd[23:16]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 i_cmd_id_3__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[3]), .o_cmd_1(
        o_inner_cmd_wire[11]), .o_cmd_2(o_inner_cmd_wire[19]), .o_cmd_3(
        o_inner_cmd_wire[27]), .o_cmd_4(o_inner_cmd_wire[35]), .o_cmd_5(
        o_inner_cmd_wire[43]), .o_cmd_6(o_inner_cmd_wire[51]), .o_cmd_7(
        o_inner_cmd_wire[59]), .i_en(i_en), .i_cmd(i_cmd[31:24]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 i_cmd_id_4__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[4]), .o_cmd_1(
        o_inner_cmd_wire[12]), .o_cmd_2(o_inner_cmd_wire[20]), .o_cmd_3(
        o_inner_cmd_wire[28]), .o_cmd_4(o_inner_cmd_wire[36]), .o_cmd_5(
        o_inner_cmd_wire[44]), .o_cmd_6(o_inner_cmd_wire[52]), .o_cmd_7(
        o_inner_cmd_wire[60]), .i_en(i_en), .i_cmd(i_cmd[39:32]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 i_cmd_id_5__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[5]), .o_cmd_1(
        o_inner_cmd_wire[13]), .o_cmd_2(o_inner_cmd_wire[21]), .o_cmd_3(
        o_inner_cmd_wire[29]), .o_cmd_4(o_inner_cmd_wire[37]), .o_cmd_5(
        o_inner_cmd_wire[45]), .o_cmd_6(o_inner_cmd_wire[53]), .o_cmd_7(
        o_inner_cmd_wire[61]), .i_en(i_en), .i_cmd(i_cmd[47:40]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 i_cmd_id_6__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[6]), .o_cmd_1(
        o_inner_cmd_wire[14]), .o_cmd_2(o_inner_cmd_wire[22]), .o_cmd_3(
        o_inner_cmd_wire[30]), .o_cmd_4(o_inner_cmd_wire[38]), .o_cmd_5(
        o_inner_cmd_wire[46]), .o_cmd_6(o_inner_cmd_wire[54]), .o_cmd_7(
        o_inner_cmd_wire[62]), .i_en(i_en), .i_cmd(i_cmd[55:48]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 i_cmd_id_7__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(o_inner_cmd_wire[7]), .o_cmd_1(
        o_inner_cmd_wire[15]), .o_cmd_2(o_inner_cmd_wire[23]), .o_cmd_3(
        o_inner_cmd_wire[31]), .o_cmd_4(o_inner_cmd_wire[39]), .o_cmd_5(
        o_inner_cmd_wire[47]), .o_cmd_6(o_inner_cmd_wire[55]), .o_cmd_7(
        o_inner_cmd_wire[63]), .i_en(i_en), .i_cmd(i_cmd[63:56]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_8 bottom_half_0__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_0__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_0__inner_data_i_mux_tree_wire), .o_valid(o_valid[0]), 
        .o_data_bus(o_data_bus[31:0]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[7:0]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_7 bottom_half_1__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_1__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_1__inner_data_i_mux_tree_wire), .o_valid(o_valid[1]), 
        .o_data_bus(o_data_bus[63:32]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[15:8]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_6 bottom_half_2__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_2__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_2__inner_data_i_mux_tree_wire), .o_valid(o_valid[2]), 
        .o_data_bus(o_data_bus[95:64]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[23:16]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_5 bottom_half_3__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_3__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_3__inner_data_i_mux_tree_wire), .o_valid(o_valid[3]), 
        .o_data_bus(o_data_bus[127:96]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[31:24]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_4 bottom_half_4__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_4__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_4__inner_data_i_mux_tree_wire), .o_valid(o_valid[4]), 
        .o_data_bus(o_data_bus[159:128]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[39:32]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_3 bottom_half_5__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_5__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_5__inner_data_i_mux_tree_wire), .o_valid(o_valid[5]), 
        .o_data_bus(o_data_bus[191:160]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[47:40]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_2 bottom_half_6__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_6__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_6__inner_data_i_mux_tree_wire), .o_valid(o_valid[6]), 
        .o_data_bus(o_data_bus[223:192]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[55:48]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_1 bottom_half_7__mux_tree ( 
        .clk(clk), .rst(rst), .i_valid(
        bottom_half_7__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_7__inner_data_i_mux_tree_wire), .o_valid(o_valid[7]), 
        .o_data_bus(o_data_bus[255:224]), .i_en(i_en), .i_cmd(
        o_inner_cmd_wire[63:56]) );
endmodule


module crossbar_one_hot_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [15:0] i_valid;
  input [511:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [127:0] i_cmd;
  input clk, rst, i_en;
  wire   N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129,
         N130, N131, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N268,
         N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279,
         N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290,
         N291, N292, N293, N294, N295, N296, N297, N298, N299, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N392, N401, N410, N419,
         N428, N437, N446, N455, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51;
  wire   [7:0] first_stage_output_def_0__o_valid_wire;
  wire   [255:0] first_stage_output_def_0__o_data_bus_wire;
  wire   [7:0] first_stage_output_def_1__o_valid_wire;
  wire   [255:0] first_stage_output_def_1__o_data_bus_wire;

  crossbar_8_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA8_0 xbar_8_8_0__xba8_8 ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[7:0]), .i_data_bus(
        i_data_bus[255:0]), .o_valid(first_stage_output_def_0__o_valid_wire), 
        .o_data_bus(first_stage_output_def_0__o_data_bus_wire), .i_en(i_en), 
        .i_cmd(i_cmd[63:0]) );
  crossbar_8_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA8_1 xbar_8_8_1__xba8_8 ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[15:8]), .i_data_bus(
        i_data_bus[511:256]), .o_valid(first_stage_output_def_1__o_valid_wire), 
        .o_data_bus(first_stage_output_def_1__o_data_bus_wire), .i_en(i_en), 
        .i_cmd(i_cmd[127:64]) );
  EDFQD4BWP30P140LVT o_valid_reg_reg_7_ ( .D(N455), .E(n51), .CP(clk), .Q(
        o_valid[7]) );
  EDFQD4BWP30P140LVT o_valid_reg_reg_6_ ( .D(N446), .E(n51), .CP(clk), .Q(
        o_valid[6]) );
  EDFQD4BWP30P140LVT o_valid_reg_reg_5_ ( .D(N437), .E(n50), .CP(clk), .Q(
        o_valid[5]) );
  EDFQD4BWP30P140LVT o_valid_reg_reg_4_ ( .D(N428), .E(n51), .CP(clk), .Q(
        o_valid[4]) );
  EDFQD4BWP30P140LVT o_valid_reg_reg_3_ ( .D(N419), .E(n51), .CP(clk), .Q(
        o_valid[3]) );
  EDFQD4BWP30P140LVT o_valid_reg_reg_2_ ( .D(N410), .E(n51), .CP(clk), .Q(
        o_valid[2]) );
  EDFQD4BWP30P140LVT o_valid_reg_reg_1_ ( .D(N401), .E(n50), .CP(clk), .Q(
        o_valid[1]) );
  EDFQD4BWP30P140LVT o_valid_reg_reg_0_ ( .D(N392), .E(n51), .CP(clk), .Q(
        o_valid[0]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N383), .E(n50), .CP(clk), 
        .Q(o_data_bus[255]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N382), .E(n51), .CP(clk), 
        .Q(o_data_bus[254]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N381), .E(n50), .CP(clk), 
        .Q(o_data_bus[253]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N380), .E(n51), .CP(clk), 
        .Q(o_data_bus[252]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N379), .E(n50), .CP(clk), 
        .Q(o_data_bus[251]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N378), .E(n50), .CP(clk), 
        .Q(o_data_bus[250]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N377), .E(n50), .CP(clk), 
        .Q(o_data_bus[249]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N376), .E(n50), .CP(clk), 
        .Q(o_data_bus[248]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N375), .E(n50), .CP(clk), 
        .Q(o_data_bus[247]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N374), .E(n50), .CP(clk), 
        .Q(o_data_bus[246]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N373), .E(n50), .CP(clk), 
        .Q(o_data_bus[245]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N372), .E(n50), .CP(clk), 
        .Q(o_data_bus[244]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N371), .E(n50), .CP(clk), 
        .Q(o_data_bus[243]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N370), .E(n50), .CP(clk), 
        .Q(o_data_bus[242]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N369), .E(n50), .CP(clk), 
        .Q(o_data_bus[241]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N368), .E(n50), .CP(clk), 
        .Q(o_data_bus[240]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N367), .E(n50), .CP(clk), 
        .Q(o_data_bus[239]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N366), .E(n50), .CP(clk), 
        .Q(o_data_bus[238]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N365), .E(n50), .CP(clk), 
        .Q(o_data_bus[237]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N364), .E(n50), .CP(clk), 
        .Q(o_data_bus[236]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N363), .E(n50), .CP(clk), 
        .Q(o_data_bus[235]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N362), .E(n50), .CP(clk), 
        .Q(o_data_bus[234]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N361), .E(n50), .CP(clk), 
        .Q(o_data_bus[233]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N360), .E(n50), .CP(clk), 
        .Q(o_data_bus[232]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N359), .E(n50), .CP(clk), 
        .Q(o_data_bus[231]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N358), .E(n50), .CP(clk), 
        .Q(o_data_bus[230]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N357), .E(n50), .CP(clk), 
        .Q(o_data_bus[229]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N356), .E(n50), .CP(clk), 
        .Q(o_data_bus[228]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N355), .E(n50), .CP(clk), 
        .Q(o_data_bus[227]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N354), .E(n50), .CP(clk), 
        .Q(o_data_bus[226]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N353), .E(n50), .CP(clk), 
        .Q(o_data_bus[225]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N352), .E(n51), .CP(clk), 
        .Q(o_data_bus[224]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N341), .E(n50), .CP(clk), 
        .Q(o_data_bus[223]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N340), .E(n51), .CP(clk), 
        .Q(o_data_bus[222]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N339), .E(n50), .CP(clk), 
        .Q(o_data_bus[221]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N338), .E(n50), .CP(clk), 
        .Q(o_data_bus[220]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N337), .E(n50), .CP(clk), 
        .Q(o_data_bus[219]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N336), .E(n51), .CP(clk), 
        .Q(o_data_bus[218]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N335), .E(n50), .CP(clk), 
        .Q(o_data_bus[217]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N334), .E(n50), .CP(clk), 
        .Q(o_data_bus[216]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N333), .E(n50), .CP(clk), 
        .Q(o_data_bus[215]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N332), .E(n51), .CP(clk), 
        .Q(o_data_bus[214]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N331), .E(n50), .CP(clk), 
        .Q(o_data_bus[213]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N330), .E(n50), .CP(clk), 
        .Q(o_data_bus[212]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N329), .E(n50), .CP(clk), 
        .Q(o_data_bus[211]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N328), .E(n50), .CP(clk), 
        .Q(o_data_bus[210]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N327), .E(n51), .CP(clk), 
        .Q(o_data_bus[209]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N326), .E(n50), .CP(clk), 
        .Q(o_data_bus[208]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N325), .E(n50), .CP(clk), 
        .Q(o_data_bus[207]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N324), .E(n51), .CP(clk), 
        .Q(o_data_bus[206]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N323), .E(n50), .CP(clk), 
        .Q(o_data_bus[205]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N322), .E(n50), .CP(clk), 
        .Q(o_data_bus[204]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N321), .E(n50), .CP(clk), 
        .Q(o_data_bus[203]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N320), .E(n50), .CP(clk), 
        .Q(o_data_bus[202]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N319), .E(n50), .CP(clk), 
        .Q(o_data_bus[201]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N318), .E(n50), .CP(clk), 
        .Q(o_data_bus[200]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N317), .E(n50), .CP(clk), 
        .Q(o_data_bus[199]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N316), .E(n50), .CP(clk), 
        .Q(o_data_bus[198]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N315), .E(n51), .CP(clk), 
        .Q(o_data_bus[197]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N314), .E(n50), .CP(clk), 
        .Q(o_data_bus[196]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N313), .E(n50), .CP(clk), 
        .Q(o_data_bus[195]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N312), .E(n50), .CP(clk), 
        .Q(o_data_bus[194]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N311), .E(n50), .CP(clk), 
        .Q(o_data_bus[193]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N310), .E(n51), .CP(clk), 
        .Q(o_data_bus[192]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N299), .E(n50), .CP(clk), 
        .Q(o_data_bus[191]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N298), .E(n50), .CP(clk), 
        .Q(o_data_bus[190]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N297), .E(n50), .CP(clk), 
        .Q(o_data_bus[189]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N296), .E(n50), .CP(clk), 
        .Q(o_data_bus[188]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N295), .E(n50), .CP(clk), 
        .Q(o_data_bus[187]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N294), .E(n50), .CP(clk), 
        .Q(o_data_bus[186]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N293), .E(n50), .CP(clk), 
        .Q(o_data_bus[185]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N292), .E(n50), .CP(clk), 
        .Q(o_data_bus[184]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N291), .E(n50), .CP(clk), 
        .Q(o_data_bus[183]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N290), .E(n50), .CP(clk), 
        .Q(o_data_bus[182]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N289), .E(n50), .CP(clk), 
        .Q(o_data_bus[181]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N288), .E(n50), .CP(clk), 
        .Q(o_data_bus[180]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N287), .E(n50), .CP(clk), 
        .Q(o_data_bus[179]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N286), .E(n50), .CP(clk), 
        .Q(o_data_bus[178]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N285), .E(n50), .CP(clk), 
        .Q(o_data_bus[177]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N284), .E(n50), .CP(clk), 
        .Q(o_data_bus[176]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N283), .E(n50), .CP(clk), 
        .Q(o_data_bus[175]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N282), .E(n50), .CP(clk), 
        .Q(o_data_bus[174]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N281), .E(n50), .CP(clk), 
        .Q(o_data_bus[173]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N280), .E(n50), .CP(clk), 
        .Q(o_data_bus[172]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N279), .E(n50), .CP(clk), 
        .Q(o_data_bus[171]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N278), .E(n50), .CP(clk), 
        .Q(o_data_bus[170]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N277), .E(n50), .CP(clk), 
        .Q(o_data_bus[169]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N276), .E(n50), .CP(clk), 
        .Q(o_data_bus[168]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N275), .E(n50), .CP(clk), 
        .Q(o_data_bus[167]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N274), .E(n50), .CP(clk), 
        .Q(o_data_bus[166]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N273), .E(n50), .CP(clk), 
        .Q(o_data_bus[165]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N272), .E(n50), .CP(clk), 
        .Q(o_data_bus[164]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N271), .E(n50), .CP(clk), 
        .Q(o_data_bus[163]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N270), .E(n50), .CP(clk), 
        .Q(o_data_bus[162]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N269), .E(n50), .CP(clk), 
        .Q(o_data_bus[161]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N268), .E(n50), .CP(clk), 
        .Q(o_data_bus[160]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N257), .E(n50), .CP(clk), 
        .Q(o_data_bus[159]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N256), .E(n50), .CP(clk), 
        .Q(o_data_bus[158]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N255), .E(n50), .CP(clk), 
        .Q(o_data_bus[157]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N254), .E(n50), .CP(clk), 
        .Q(o_data_bus[156]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N253), .E(n50), .CP(clk), 
        .Q(o_data_bus[155]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N252), .E(n50), .CP(clk), 
        .Q(o_data_bus[154]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N251), .E(n50), .CP(clk), 
        .Q(o_data_bus[153]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N250), .E(n50), .CP(clk), 
        .Q(o_data_bus[152]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N249), .E(n50), .CP(clk), 
        .Q(o_data_bus[151]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N248), .E(n50), .CP(clk), 
        .Q(o_data_bus[150]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N247), .E(n50), .CP(clk), 
        .Q(o_data_bus[149]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N246), .E(n50), .CP(clk), 
        .Q(o_data_bus[148]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N245), .E(n50), .CP(clk), 
        .Q(o_data_bus[147]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N244), .E(n51), .CP(clk), 
        .Q(o_data_bus[146]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N243), .E(n51), .CP(clk), 
        .Q(o_data_bus[145]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N242), .E(n51), .CP(clk), 
        .Q(o_data_bus[144]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N241), .E(n50), .CP(clk), 
        .Q(o_data_bus[143]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N240), .E(n51), .CP(clk), 
        .Q(o_data_bus[142]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N239), .E(n50), .CP(clk), 
        .Q(o_data_bus[141]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N238), .E(n51), .CP(clk), 
        .Q(o_data_bus[140]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N237), .E(n51), .CP(clk), 
        .Q(o_data_bus[139]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N236), .E(n51), .CP(clk), 
        .Q(o_data_bus[138]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N235), .E(n51), .CP(clk), 
        .Q(o_data_bus[137]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N234), .E(n51), .CP(clk), 
        .Q(o_data_bus[136]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N233), .E(n50), .CP(clk), 
        .Q(o_data_bus[135]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N232), .E(n51), .CP(clk), 
        .Q(o_data_bus[134]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N231), .E(n51), .CP(clk), 
        .Q(o_data_bus[133]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N230), .E(n51), .CP(clk), 
        .Q(o_data_bus[132]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N229), .E(n50), .CP(clk), 
        .Q(o_data_bus[131]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N228), .E(n51), .CP(clk), 
        .Q(o_data_bus[130]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N227), .E(n51), .CP(clk), 
        .Q(o_data_bus[129]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N226), .E(n50), .CP(clk), 
        .Q(o_data_bus[128]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N215), .E(n51), .CP(clk), 
        .Q(o_data_bus[127]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N214), .E(n51), .CP(clk), 
        .Q(o_data_bus[126]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N213), .E(n51), .CP(clk), 
        .Q(o_data_bus[125]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N212), .E(n51), .CP(clk), 
        .Q(o_data_bus[124]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N211), .E(n50), .CP(clk), 
        .Q(o_data_bus[123]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N210), .E(n51), .CP(clk), 
        .Q(o_data_bus[122]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N209), .E(n51), .CP(clk), 
        .Q(o_data_bus[121]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N208), .E(n51), .CP(clk), 
        .Q(o_data_bus[120]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N207), .E(n51), .CP(clk), 
        .Q(o_data_bus[119]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N206), .E(n51), .CP(clk), 
        .Q(o_data_bus[118]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N205), .E(n51), .CP(clk), 
        .Q(o_data_bus[117]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N204), .E(n50), .CP(clk), 
        .Q(o_data_bus[116]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N203), .E(n51), .CP(clk), 
        .Q(o_data_bus[115]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N202), .E(n51), .CP(clk), 
        .Q(o_data_bus[114]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N201), .E(n51), .CP(clk), 
        .Q(o_data_bus[113]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N200), .E(n51), .CP(clk), 
        .Q(o_data_bus[112]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N199), .E(n51), .CP(clk), 
        .Q(o_data_bus[111]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N198), .E(n51), .CP(clk), 
        .Q(o_data_bus[110]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N197), .E(n51), .CP(clk), 
        .Q(o_data_bus[109]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N196), .E(n50), .CP(clk), 
        .Q(o_data_bus[108]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N195), .E(n50), .CP(clk), 
        .Q(o_data_bus[107]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N194), .E(n50), .CP(clk), 
        .Q(o_data_bus[106]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N193), .E(n50), .CP(clk), 
        .Q(o_data_bus[105]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N192), .E(n50), .CP(clk), 
        .Q(o_data_bus[104]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N191), .E(n50), .CP(clk), 
        .Q(o_data_bus[103]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N190), .E(n50), .CP(clk), 
        .Q(o_data_bus[102]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N189), .E(n50), .CP(clk), 
        .Q(o_data_bus[101]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N188), .E(n50), .CP(clk), 
        .Q(o_data_bus[100]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N187), .E(n50), .CP(clk), .Q(
        o_data_bus[99]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N186), .E(n50), .CP(clk), .Q(
        o_data_bus[98]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N185), .E(n50), .CP(clk), .Q(
        o_data_bus[97]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N184), .E(n50), .CP(clk), .Q(
        o_data_bus[96]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N173), .E(n50), .CP(clk), .Q(
        o_data_bus[95]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N172), .E(n50), .CP(clk), .Q(
        o_data_bus[94]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N171), .E(n50), .CP(clk), .Q(
        o_data_bus[93]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N170), .E(n50), .CP(clk), .Q(
        o_data_bus[92]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N169), .E(n50), .CP(clk), .Q(
        o_data_bus[91]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N168), .E(n50), .CP(clk), .Q(
        o_data_bus[90]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N167), .E(n50), .CP(clk), .Q(
        o_data_bus[89]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N166), .E(n50), .CP(clk), .Q(
        o_data_bus[88]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N165), .E(n50), .CP(clk), .Q(
        o_data_bus[87]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N164), .E(n50), .CP(clk), .Q(
        o_data_bus[86]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N163), .E(n50), .CP(clk), .Q(
        o_data_bus[85]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N162), .E(n50), .CP(clk), .Q(
        o_data_bus[84]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N161), .E(n50), .CP(clk), .Q(
        o_data_bus[83]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N160), .E(n50), .CP(clk), .Q(
        o_data_bus[82]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N159), .E(n50), .CP(clk), .Q(
        o_data_bus[81]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N158), .E(n50), .CP(clk), .Q(
        o_data_bus[80]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N157), .E(n50), .CP(clk), .Q(
        o_data_bus[79]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N156), .E(n50), .CP(clk), .Q(
        o_data_bus[78]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N155), .E(n50), .CP(clk), .Q(
        o_data_bus[77]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N154), .E(n50), .CP(clk), .Q(
        o_data_bus[76]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N153), .E(n50), .CP(clk), .Q(
        o_data_bus[75]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N152), .E(n50), .CP(clk), .Q(
        o_data_bus[74]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N151), .E(n50), .CP(clk), .Q(
        o_data_bus[73]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N150), .E(n50), .CP(clk), .Q(
        o_data_bus[72]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N149), .E(n50), .CP(clk), .Q(
        o_data_bus[71]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N148), .E(n50), .CP(clk), .Q(
        o_data_bus[70]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N147), .E(n50), .CP(clk), .Q(
        o_data_bus[69]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N146), .E(n50), .CP(clk), .Q(
        o_data_bus[68]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N145), .E(n50), .CP(clk), .Q(
        o_data_bus[67]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N144), .E(n50), .CP(clk), .Q(
        o_data_bus[66]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N143), .E(n50), .CP(clk), .Q(
        o_data_bus[65]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N142), .E(n50), .CP(clk), .Q(
        o_data_bus[64]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N131), .E(n50), .CP(clk), .Q(
        o_data_bus[63]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N130), .E(n50), .CP(clk), .Q(
        o_data_bus[62]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N129), .E(n50), .CP(clk), .Q(
        o_data_bus[61]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N128), .E(n50), .CP(clk), .Q(
        o_data_bus[60]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N127), .E(n50), .CP(clk), .Q(
        o_data_bus[59]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N126), .E(n50), .CP(clk), .Q(
        o_data_bus[58]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N125), .E(n50), .CP(clk), .Q(
        o_data_bus[57]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N124), .E(n50), .CP(clk), .Q(
        o_data_bus[56]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N123), .E(n50), .CP(clk), .Q(
        o_data_bus[55]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N122), .E(n50), .CP(clk), .Q(
        o_data_bus[54]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N121), .E(n50), .CP(clk), .Q(
        o_data_bus[53]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N120), .E(n50), .CP(clk), .Q(
        o_data_bus[52]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N119), .E(n50), .CP(clk), .Q(
        o_data_bus[51]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N118), .E(n50), .CP(clk), .Q(
        o_data_bus[50]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N117), .E(n50), .CP(clk), .Q(
        o_data_bus[49]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N116), .E(n50), .CP(clk), .Q(
        o_data_bus[48]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N115), .E(n50), .CP(clk), .Q(
        o_data_bus[47]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N114), .E(n50), .CP(clk), .Q(
        o_data_bus[46]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N113), .E(n50), .CP(clk), .Q(
        o_data_bus[45]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N112), .E(n50), .CP(clk), .Q(
        o_data_bus[44]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N111), .E(n50), .CP(clk), .Q(
        o_data_bus[43]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N110), .E(n50), .CP(clk), .Q(
        o_data_bus[42]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N109), .E(n50), .CP(clk), .Q(
        o_data_bus[41]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N108), .E(n50), .CP(clk), .Q(
        o_data_bus[40]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N107), .E(n50), .CP(clk), .Q(
        o_data_bus[39]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N106), .E(n50), .CP(clk), .Q(
        o_data_bus[38]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N105), .E(n50), .CP(clk), .Q(
        o_data_bus[37]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N104), .E(n50), .CP(clk), .Q(
        o_data_bus[36]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N103), .E(n50), .CP(clk), .Q(
        o_data_bus[35]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N102), .E(n50), .CP(clk), .Q(
        o_data_bus[34]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N101), .E(n50), .CP(clk), .Q(
        o_data_bus[33]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N100), .E(n50), .CP(clk), .Q(
        o_data_bus[32]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N89), .E(n50), .CP(clk), .Q(
        o_data_bus[31]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N88), .E(n50), .CP(clk), .Q(
        o_data_bus[30]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N87), .E(n51), .CP(clk), .Q(
        o_data_bus[29]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N86), .E(n51), .CP(clk), .Q(
        o_data_bus[28]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N85), .E(n50), .CP(clk), .Q(
        o_data_bus[27]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N84), .E(n51), .CP(clk), .Q(
        o_data_bus[26]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N83), .E(n51), .CP(clk), .Q(
        o_data_bus[25]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N82), .E(n50), .CP(clk), .Q(
        o_data_bus[24]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N81), .E(n51), .CP(clk), .Q(
        o_data_bus[23]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N80), .E(n51), .CP(clk), .Q(
        o_data_bus[22]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N79), .E(n51), .CP(clk), .Q(
        o_data_bus[21]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N78), .E(n51), .CP(clk), .Q(
        o_data_bus[20]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N77), .E(n50), .CP(clk), .Q(
        o_data_bus[19]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N76), .E(n51), .CP(clk), .Q(
        o_data_bus[18]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N75), .E(n51), .CP(clk), .Q(
        o_data_bus[17]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N74), .E(n50), .CP(clk), .Q(
        o_data_bus[16]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N73), .E(n51), .CP(clk), .Q(
        o_data_bus[15]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N72), .E(n50), .CP(clk), .Q(
        o_data_bus[14]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N71), .E(n51), .CP(clk), .Q(
        o_data_bus[13]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N70), .E(n51), .CP(clk), .Q(
        o_data_bus[12]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N69), .E(n50), .CP(clk), .Q(
        o_data_bus[11]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N68), .E(n51), .CP(clk), .Q(
        o_data_bus[10]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N67), .E(n51), .CP(clk), .Q(
        o_data_bus[9]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N66), .E(n50), .CP(clk), .Q(
        o_data_bus[8]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N65), .E(n51), .CP(clk), .Q(
        o_data_bus[7]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N64), .E(n50), .CP(clk), .Q(
        o_data_bus[6]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N63), .E(n51), .CP(clk), .Q(
        o_data_bus[5]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N62), .E(n51), .CP(clk), .Q(
        o_data_bus[4]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N61), .E(n51), .CP(clk), .Q(
        o_data_bus[3]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N60), .E(n51), .CP(clk), .Q(
        o_data_bus[2]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N59), .E(n51), .CP(clk), .Q(
        o_data_bus[1]) );
  EDFQD4BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N58), .E(n51), .CP(clk), .Q(
        o_data_bus[0]) );
  ND2OPTIBD1BWP30P140LVT U283 ( .A1(n43), .A2(n42), .ZN(N428) );
  ND2OPTIBD1BWP30P140LVT U284 ( .A1(n45), .A2(n44), .ZN(N437) );
  ND2OPTIBD1BWP30P140LVT U285 ( .A1(n41), .A2(n40), .ZN(N419) );
  ND2OPTIBD1BWP30P140LVT U286 ( .A1(n39), .A2(n38), .ZN(N410) );
  ND2OPTIBD1BWP30P140LVT U287 ( .A1(n47), .A2(n46), .ZN(N446) );
  ND2OPTIBD1BWP30P140LVT U288 ( .A1(n37), .A2(n36), .ZN(N401) );
  ND2OPTIBD1BWP30P140LVT U289 ( .A1(n35), .A2(n34), .ZN(N392) );
  ND2OPTIBD1BWP30P140LVT U290 ( .A1(n49), .A2(n48), .ZN(N455) );
  BUFFD2BWP30P140LVT U291 ( .I(n51), .Z(n50) );
  INVD1BWP30P140LVT U292 ( .I(i_en), .ZN(n17) );
  NR2D1BWP30P140LVT U293 ( .A1(rst), .A2(n17), .ZN(n51) );
  IND2D1BWP30P140LVT U294 ( .A1(first_stage_output_def_0__o_valid_wire[0]), 
        .B1(first_stage_output_def_1__o_valid_wire[0]), .ZN(n35) );
  INVD2BWP30P140LVT U295 ( .I(n35), .ZN(n19) );
  IND2D1BWP30P140LVT U296 ( .A1(first_stage_output_def_1__o_valid_wire[0]), 
        .B1(first_stage_output_def_0__o_valid_wire[0]), .ZN(n34) );
  INVD2BWP30P140LVT U297 ( .I(n34), .ZN(n18) );
  AO22D1BWP30P140LVT U298 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[0]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[0]), .Z(N58) );
  AO22D1BWP30P140LVT U299 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[1]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[1]), .Z(N59) );
  AO22D1BWP30P140LVT U300 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[2]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[2]), .Z(N60) );
  AO22D1BWP30P140LVT U301 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[3]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[3]), .Z(N61) );
  AO22D1BWP30P140LVT U302 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[4]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[4]), .Z(N62) );
  AO22D1BWP30P140LVT U303 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[5]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[5]), .Z(N63) );
  AO22D1BWP30P140LVT U304 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[6]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[6]), .Z(N64) );
  AO22D1BWP30P140LVT U305 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[7]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[7]), .Z(N65) );
  AO22D1BWP30P140LVT U306 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[8]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[8]), .Z(N66) );
  AO22D1BWP30P140LVT U307 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[9]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[9]), .Z(N67) );
  AO22D1BWP30P140LVT U308 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[10]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[10]), .Z(N68) );
  AO22D1BWP30P140LVT U309 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[11]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[11]), .Z(N69) );
  AO22D1BWP30P140LVT U310 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[12]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[12]), .Z(N70) );
  AO22D1BWP30P140LVT U311 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[13]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[13]), .Z(N71) );
  AO22D1BWP30P140LVT U312 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[14]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[14]), .Z(N72) );
  AO22D1BWP30P140LVT U313 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[15]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[15]), .Z(N73) );
  AO22D1BWP30P140LVT U314 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[16]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[16]), .Z(N74) );
  AO22D1BWP30P140LVT U315 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[17]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[17]), .Z(N75) );
  AO22D1BWP30P140LVT U316 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[18]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[18]), .Z(N76) );
  AO22D1BWP30P140LVT U317 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[19]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[19]), .Z(N77) );
  AO22D1BWP30P140LVT U318 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[20]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[20]), .Z(N78) );
  AO22D1BWP30P140LVT U319 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[21]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[21]), .Z(N79) );
  AO22D1BWP30P140LVT U320 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[22]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[22]), .Z(N80) );
  AO22D1BWP30P140LVT U321 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[23]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[23]), .Z(N81) );
  AO22D1BWP30P140LVT U322 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[24]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[24]), .Z(N82) );
  AO22D1BWP30P140LVT U323 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[25]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[25]), .Z(N83) );
  AO22D1BWP30P140LVT U324 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[26]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[26]), .Z(N84) );
  AO22D1BWP30P140LVT U325 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[27]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[27]), .Z(N85) );
  AO22D1BWP30P140LVT U326 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[28]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[28]), .Z(N86) );
  AO22D1BWP30P140LVT U327 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[29]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[29]), .Z(N87) );
  AO22D1BWP30P140LVT U328 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[30]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[30]), .Z(N88) );
  AO22D1BWP30P140LVT U329 ( .A1(n19), .A2(
        first_stage_output_def_1__o_data_bus_wire[31]), .B1(n18), .B2(
        first_stage_output_def_0__o_data_bus_wire[31]), .Z(N89) );
  IND2D1BWP30P140LVT U330 ( .A1(first_stage_output_def_0__o_valid_wire[1]), 
        .B1(first_stage_output_def_1__o_valid_wire[1]), .ZN(n37) );
  INVD2BWP30P140LVT U331 ( .I(n37), .ZN(n21) );
  IND2D1BWP30P140LVT U332 ( .A1(first_stage_output_def_1__o_valid_wire[1]), 
        .B1(first_stage_output_def_0__o_valid_wire[1]), .ZN(n36) );
  INVD2BWP30P140LVT U333 ( .I(n36), .ZN(n20) );
  AO22D1BWP30P140LVT U334 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[32]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[32]), .Z(N100) );
  AO22D1BWP30P140LVT U335 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[33]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[33]), .Z(N101) );
  AO22D1BWP30P140LVT U336 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[34]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[34]), .Z(N102) );
  AO22D1BWP30P140LVT U337 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[35]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[35]), .Z(N103) );
  AO22D1BWP30P140LVT U338 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[36]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[36]), .Z(N104) );
  AO22D1BWP30P140LVT U339 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[37]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[37]), .Z(N105) );
  AO22D1BWP30P140LVT U340 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[38]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[38]), .Z(N106) );
  AO22D1BWP30P140LVT U341 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[39]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[39]), .Z(N107) );
  AO22D1BWP30P140LVT U342 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[40]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[40]), .Z(N108) );
  AO22D1BWP30P140LVT U343 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[41]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[41]), .Z(N109) );
  AO22D1BWP30P140LVT U344 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[42]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[42]), .Z(N110) );
  AO22D1BWP30P140LVT U345 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[43]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[43]), .Z(N111) );
  AO22D1BWP30P140LVT U346 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[44]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[44]), .Z(N112) );
  AO22D1BWP30P140LVT U347 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[45]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[45]), .Z(N113) );
  AO22D1BWP30P140LVT U348 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[46]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[46]), .Z(N114) );
  AO22D1BWP30P140LVT U349 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[47]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[47]), .Z(N115) );
  AO22D1BWP30P140LVT U350 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[48]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[48]), .Z(N116) );
  AO22D1BWP30P140LVT U351 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[49]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[49]), .Z(N117) );
  AO22D1BWP30P140LVT U352 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[50]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[50]), .Z(N118) );
  AO22D1BWP30P140LVT U353 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[51]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[51]), .Z(N119) );
  AO22D1BWP30P140LVT U354 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[52]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[52]), .Z(N120) );
  AO22D1BWP30P140LVT U355 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[53]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[53]), .Z(N121) );
  AO22D1BWP30P140LVT U356 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[54]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[54]), .Z(N122) );
  AO22D1BWP30P140LVT U357 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[55]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[55]), .Z(N123) );
  AO22D1BWP30P140LVT U358 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[56]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[56]), .Z(N124) );
  AO22D1BWP30P140LVT U359 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[57]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[57]), .Z(N125) );
  AO22D1BWP30P140LVT U360 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[58]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[58]), .Z(N126) );
  AO22D1BWP30P140LVT U361 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[59]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[59]), .Z(N127) );
  AO22D1BWP30P140LVT U362 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[60]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[60]), .Z(N128) );
  AO22D1BWP30P140LVT U363 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[61]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[61]), .Z(N129) );
  AO22D1BWP30P140LVT U364 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[62]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[62]), .Z(N130) );
  AO22D1BWP30P140LVT U365 ( .A1(n21), .A2(
        first_stage_output_def_1__o_data_bus_wire[63]), .B1(n20), .B2(
        first_stage_output_def_0__o_data_bus_wire[63]), .Z(N131) );
  IND2D1BWP30P140LVT U366 ( .A1(first_stage_output_def_0__o_valid_wire[2]), 
        .B1(first_stage_output_def_1__o_valid_wire[2]), .ZN(n39) );
  INVD2BWP30P140LVT U367 ( .I(n39), .ZN(n23) );
  IND2D1BWP30P140LVT U368 ( .A1(first_stage_output_def_1__o_valid_wire[2]), 
        .B1(first_stage_output_def_0__o_valid_wire[2]), .ZN(n38) );
  INVD2BWP30P140LVT U369 ( .I(n38), .ZN(n22) );
  AO22D1BWP30P140LVT U370 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[64]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[64]), .Z(N142) );
  AO22D1BWP30P140LVT U371 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[65]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[65]), .Z(N143) );
  AO22D1BWP30P140LVT U372 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[66]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[66]), .Z(N144) );
  AO22D1BWP30P140LVT U373 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[67]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[67]), .Z(N145) );
  AO22D1BWP30P140LVT U374 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[68]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[68]), .Z(N146) );
  AO22D1BWP30P140LVT U375 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[69]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[69]), .Z(N147) );
  AO22D1BWP30P140LVT U376 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[70]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[70]), .Z(N148) );
  AO22D1BWP30P140LVT U377 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[71]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[71]), .Z(N149) );
  AO22D1BWP30P140LVT U378 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[72]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[72]), .Z(N150) );
  AO22D1BWP30P140LVT U379 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[73]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[73]), .Z(N151) );
  AO22D1BWP30P140LVT U380 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[74]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[74]), .Z(N152) );
  AO22D1BWP30P140LVT U381 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[75]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[75]), .Z(N153) );
  AO22D1BWP30P140LVT U382 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[76]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[76]), .Z(N154) );
  AO22D1BWP30P140LVT U383 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[77]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[77]), .Z(N155) );
  AO22D1BWP30P140LVT U384 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[78]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[78]), .Z(N156) );
  AO22D1BWP30P140LVT U385 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[79]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[79]), .Z(N157) );
  AO22D1BWP30P140LVT U386 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[80]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[80]), .Z(N158) );
  AO22D1BWP30P140LVT U387 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[81]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[81]), .Z(N159) );
  AO22D1BWP30P140LVT U388 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[82]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[82]), .Z(N160) );
  AO22D1BWP30P140LVT U389 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[83]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[83]), .Z(N161) );
  AO22D1BWP30P140LVT U390 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[84]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[84]), .Z(N162) );
  AO22D1BWP30P140LVT U391 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[85]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[85]), .Z(N163) );
  AO22D1BWP30P140LVT U392 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[86]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[86]), .Z(N164) );
  AO22D1BWP30P140LVT U393 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[87]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[87]), .Z(N165) );
  AO22D1BWP30P140LVT U394 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[88]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[88]), .Z(N166) );
  AO22D1BWP30P140LVT U395 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[89]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[89]), .Z(N167) );
  AO22D1BWP30P140LVT U396 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[90]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[90]), .Z(N168) );
  AO22D1BWP30P140LVT U397 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[91]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[91]), .Z(N169) );
  AO22D1BWP30P140LVT U398 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[92]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[92]), .Z(N170) );
  AO22D1BWP30P140LVT U399 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[93]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[93]), .Z(N171) );
  AO22D1BWP30P140LVT U400 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[94]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[94]), .Z(N172) );
  AO22D1BWP30P140LVT U401 ( .A1(n23), .A2(
        first_stage_output_def_1__o_data_bus_wire[95]), .B1(n22), .B2(
        first_stage_output_def_0__o_data_bus_wire[95]), .Z(N173) );
  IND2D1BWP30P140LVT U402 ( .A1(first_stage_output_def_0__o_valid_wire[3]), 
        .B1(first_stage_output_def_1__o_valid_wire[3]), .ZN(n41) );
  INVD2BWP30P140LVT U403 ( .I(n41), .ZN(n25) );
  IND2D1BWP30P140LVT U404 ( .A1(first_stage_output_def_1__o_valid_wire[3]), 
        .B1(first_stage_output_def_0__o_valid_wire[3]), .ZN(n40) );
  INVD2BWP30P140LVT U405 ( .I(n40), .ZN(n24) );
  AO22D1BWP30P140LVT U406 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[96]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[96]), .Z(N184) );
  AO22D1BWP30P140LVT U407 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[97]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[97]), .Z(N185) );
  AO22D1BWP30P140LVT U408 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[98]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[98]), .Z(N186) );
  AO22D1BWP30P140LVT U409 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[99]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[99]), .Z(N187) );
  AO22D1BWP30P140LVT U410 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[100]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[100]), .Z(N188) );
  AO22D1BWP30P140LVT U411 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[101]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[101]), .Z(N189) );
  AO22D1BWP30P140LVT U412 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[102]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[102]), .Z(N190) );
  AO22D1BWP30P140LVT U413 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[103]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[103]), .Z(N191) );
  AO22D1BWP30P140LVT U414 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[104]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[104]), .Z(N192) );
  AO22D1BWP30P140LVT U415 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[105]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[105]), .Z(N193) );
  AO22D1BWP30P140LVT U416 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[106]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[106]), .Z(N194) );
  AO22D1BWP30P140LVT U417 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[107]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[107]), .Z(N195) );
  AO22D1BWP30P140LVT U418 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[108]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[108]), .Z(N196) );
  AO22D1BWP30P140LVT U419 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[109]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[109]), .Z(N197) );
  AO22D1BWP30P140LVT U420 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[110]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[110]), .Z(N198) );
  AO22D1BWP30P140LVT U421 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[111]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[111]), .Z(N199) );
  AO22D1BWP30P140LVT U422 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[112]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[112]), .Z(N200) );
  AO22D1BWP30P140LVT U423 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[113]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[113]), .Z(N201) );
  AO22D1BWP30P140LVT U424 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[114]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[114]), .Z(N202) );
  AO22D1BWP30P140LVT U425 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[115]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[115]), .Z(N203) );
  AO22D1BWP30P140LVT U426 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[116]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[116]), .Z(N204) );
  AO22D1BWP30P140LVT U427 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[117]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[117]), .Z(N205) );
  AO22D1BWP30P140LVT U428 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[118]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[118]), .Z(N206) );
  AO22D1BWP30P140LVT U429 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[119]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[119]), .Z(N207) );
  AO22D1BWP30P140LVT U430 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[120]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[120]), .Z(N208) );
  AO22D1BWP30P140LVT U431 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[121]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[121]), .Z(N209) );
  AO22D1BWP30P140LVT U432 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[122]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[122]), .Z(N210) );
  AO22D1BWP30P140LVT U433 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[123]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[123]), .Z(N211) );
  AO22D1BWP30P140LVT U434 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[124]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[124]), .Z(N212) );
  AO22D1BWP30P140LVT U435 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[125]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[125]), .Z(N213) );
  AO22D1BWP30P140LVT U436 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[126]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[126]), .Z(N214) );
  AO22D1BWP30P140LVT U437 ( .A1(n25), .A2(
        first_stage_output_def_1__o_data_bus_wire[127]), .B1(n24), .B2(
        first_stage_output_def_0__o_data_bus_wire[127]), .Z(N215) );
  IND2D1BWP30P140LVT U438 ( .A1(first_stage_output_def_0__o_valid_wire[4]), 
        .B1(first_stage_output_def_1__o_valid_wire[4]), .ZN(n43) );
  INVD2BWP30P140LVT U439 ( .I(n43), .ZN(n27) );
  IND2D1BWP30P140LVT U440 ( .A1(first_stage_output_def_1__o_valid_wire[4]), 
        .B1(first_stage_output_def_0__o_valid_wire[4]), .ZN(n42) );
  INVD2BWP30P140LVT U441 ( .I(n42), .ZN(n26) );
  AO22D1BWP30P140LVT U442 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[128]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[128]), .Z(N226) );
  AO22D1BWP30P140LVT U443 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[129]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[129]), .Z(N227) );
  AO22D1BWP30P140LVT U444 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[130]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[130]), .Z(N228) );
  AO22D1BWP30P140LVT U445 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[131]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[131]), .Z(N229) );
  AO22D1BWP30P140LVT U446 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[132]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[132]), .Z(N230) );
  AO22D1BWP30P140LVT U447 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[133]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[133]), .Z(N231) );
  AO22D1BWP30P140LVT U448 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[134]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[134]), .Z(N232) );
  AO22D1BWP30P140LVT U449 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[135]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[135]), .Z(N233) );
  AO22D1BWP30P140LVT U450 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[136]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[136]), .Z(N234) );
  AO22D1BWP30P140LVT U451 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[137]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[137]), .Z(N235) );
  AO22D1BWP30P140LVT U452 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[138]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[138]), .Z(N236) );
  AO22D1BWP30P140LVT U453 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[139]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[139]), .Z(N237) );
  AO22D1BWP30P140LVT U454 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[140]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[140]), .Z(N238) );
  AO22D1BWP30P140LVT U455 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[141]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[141]), .Z(N239) );
  AO22D1BWP30P140LVT U456 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[142]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[142]), .Z(N240) );
  AO22D1BWP30P140LVT U457 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[143]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[143]), .Z(N241) );
  AO22D1BWP30P140LVT U458 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[144]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[144]), .Z(N242) );
  AO22D1BWP30P140LVT U459 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[145]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[145]), .Z(N243) );
  AO22D1BWP30P140LVT U460 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[146]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[146]), .Z(N244) );
  AO22D1BWP30P140LVT U461 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[147]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[147]), .Z(N245) );
  AO22D1BWP30P140LVT U462 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[148]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[148]), .Z(N246) );
  AO22D1BWP30P140LVT U463 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[149]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[149]), .Z(N247) );
  AO22D1BWP30P140LVT U464 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[150]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[150]), .Z(N248) );
  AO22D1BWP30P140LVT U465 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[151]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[151]), .Z(N249) );
  AO22D1BWP30P140LVT U466 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[152]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[152]), .Z(N250) );
  AO22D1BWP30P140LVT U467 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[153]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[153]), .Z(N251) );
  AO22D1BWP30P140LVT U468 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[154]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[154]), .Z(N252) );
  AO22D1BWP30P140LVT U469 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[155]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[155]), .Z(N253) );
  AO22D1BWP30P140LVT U470 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[156]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[156]), .Z(N254) );
  AO22D1BWP30P140LVT U471 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[157]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[157]), .Z(N255) );
  AO22D1BWP30P140LVT U472 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[158]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[158]), .Z(N256) );
  AO22D1BWP30P140LVT U473 ( .A1(n27), .A2(
        first_stage_output_def_1__o_data_bus_wire[159]), .B1(n26), .B2(
        first_stage_output_def_0__o_data_bus_wire[159]), .Z(N257) );
  IND2D1BWP30P140LVT U474 ( .A1(first_stage_output_def_0__o_valid_wire[5]), 
        .B1(first_stage_output_def_1__o_valid_wire[5]), .ZN(n45) );
  INVD2BWP30P140LVT U475 ( .I(n45), .ZN(n29) );
  IND2D1BWP30P140LVT U476 ( .A1(first_stage_output_def_1__o_valid_wire[5]), 
        .B1(first_stage_output_def_0__o_valid_wire[5]), .ZN(n44) );
  INVD2BWP30P140LVT U477 ( .I(n44), .ZN(n28) );
  AO22D1BWP30P140LVT U478 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[160]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[160]), .Z(N268) );
  AO22D1BWP30P140LVT U479 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[161]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[161]), .Z(N269) );
  AO22D1BWP30P140LVT U480 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[162]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[162]), .Z(N270) );
  AO22D1BWP30P140LVT U481 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[163]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[163]), .Z(N271) );
  AO22D1BWP30P140LVT U482 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[164]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[164]), .Z(N272) );
  AO22D1BWP30P140LVT U483 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[165]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[165]), .Z(N273) );
  AO22D1BWP30P140LVT U484 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[166]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[166]), .Z(N274) );
  AO22D1BWP30P140LVT U485 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[167]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[167]), .Z(N275) );
  AO22D1BWP30P140LVT U486 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[168]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[168]), .Z(N276) );
  AO22D1BWP30P140LVT U487 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[169]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[169]), .Z(N277) );
  AO22D1BWP30P140LVT U488 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[170]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[170]), .Z(N278) );
  AO22D1BWP30P140LVT U489 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[171]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[171]), .Z(N279) );
  AO22D1BWP30P140LVT U490 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[172]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[172]), .Z(N280) );
  AO22D1BWP30P140LVT U491 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[173]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[173]), .Z(N281) );
  AO22D1BWP30P140LVT U492 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[174]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[174]), .Z(N282) );
  AO22D1BWP30P140LVT U493 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[175]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[175]), .Z(N283) );
  AO22D1BWP30P140LVT U494 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[176]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[176]), .Z(N284) );
  AO22D1BWP30P140LVT U495 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[177]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[177]), .Z(N285) );
  AO22D1BWP30P140LVT U496 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[178]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[178]), .Z(N286) );
  AO22D1BWP30P140LVT U497 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[179]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[179]), .Z(N287) );
  AO22D1BWP30P140LVT U498 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[180]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[180]), .Z(N288) );
  AO22D1BWP30P140LVT U499 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[181]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[181]), .Z(N289) );
  AO22D1BWP30P140LVT U500 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[182]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[182]), .Z(N290) );
  AO22D1BWP30P140LVT U501 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[183]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[183]), .Z(N291) );
  AO22D1BWP30P140LVT U502 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[184]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[184]), .Z(N292) );
  AO22D1BWP30P140LVT U503 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[185]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[185]), .Z(N293) );
  AO22D1BWP30P140LVT U504 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[186]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[186]), .Z(N294) );
  AO22D1BWP30P140LVT U505 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[187]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[187]), .Z(N295) );
  AO22D1BWP30P140LVT U506 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[188]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[188]), .Z(N296) );
  AO22D1BWP30P140LVT U507 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[189]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[189]), .Z(N297) );
  AO22D1BWP30P140LVT U508 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[190]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[190]), .Z(N298) );
  AO22D1BWP30P140LVT U509 ( .A1(n29), .A2(
        first_stage_output_def_1__o_data_bus_wire[191]), .B1(n28), .B2(
        first_stage_output_def_0__o_data_bus_wire[191]), .Z(N299) );
  IND2D1BWP30P140LVT U510 ( .A1(first_stage_output_def_0__o_valid_wire[6]), 
        .B1(first_stage_output_def_1__o_valid_wire[6]), .ZN(n47) );
  INVD2BWP30P140LVT U511 ( .I(n47), .ZN(n31) );
  IND2D1BWP30P140LVT U512 ( .A1(first_stage_output_def_1__o_valid_wire[6]), 
        .B1(first_stage_output_def_0__o_valid_wire[6]), .ZN(n46) );
  INVD2BWP30P140LVT U513 ( .I(n46), .ZN(n30) );
  AO22D1BWP30P140LVT U514 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[192]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[192]), .Z(N310) );
  AO22D1BWP30P140LVT U515 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[193]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[193]), .Z(N311) );
  AO22D1BWP30P140LVT U516 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[194]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[194]), .Z(N312) );
  AO22D1BWP30P140LVT U517 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[195]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[195]), .Z(N313) );
  AO22D1BWP30P140LVT U518 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[196]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[196]), .Z(N314) );
  AO22D1BWP30P140LVT U519 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[197]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[197]), .Z(N315) );
  AO22D1BWP30P140LVT U520 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[198]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[198]), .Z(N316) );
  AO22D1BWP30P140LVT U521 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[199]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[199]), .Z(N317) );
  AO22D1BWP30P140LVT U522 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[200]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[200]), .Z(N318) );
  AO22D1BWP30P140LVT U523 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[201]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[201]), .Z(N319) );
  AO22D1BWP30P140LVT U524 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[202]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[202]), .Z(N320) );
  AO22D1BWP30P140LVT U525 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[203]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[203]), .Z(N321) );
  AO22D1BWP30P140LVT U526 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[204]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[204]), .Z(N322) );
  AO22D1BWP30P140LVT U527 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[205]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[205]), .Z(N323) );
  AO22D1BWP30P140LVT U528 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[206]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[206]), .Z(N324) );
  AO22D1BWP30P140LVT U529 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[207]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[207]), .Z(N325) );
  AO22D1BWP30P140LVT U530 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[208]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[208]), .Z(N326) );
  AO22D1BWP30P140LVT U531 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[209]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[209]), .Z(N327) );
  AO22D1BWP30P140LVT U532 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[210]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[210]), .Z(N328) );
  AO22D1BWP30P140LVT U533 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[211]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[211]), .Z(N329) );
  AO22D1BWP30P140LVT U534 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[212]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[212]), .Z(N330) );
  AO22D1BWP30P140LVT U535 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[213]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[213]), .Z(N331) );
  AO22D1BWP30P140LVT U536 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[214]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[214]), .Z(N332) );
  AO22D1BWP30P140LVT U537 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[215]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[215]), .Z(N333) );
  AO22D1BWP30P140LVT U538 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[216]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[216]), .Z(N334) );
  AO22D1BWP30P140LVT U539 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[217]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[217]), .Z(N335) );
  AO22D1BWP30P140LVT U540 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[218]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[218]), .Z(N336) );
  AO22D1BWP30P140LVT U541 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[219]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[219]), .Z(N337) );
  AO22D1BWP30P140LVT U542 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[220]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[220]), .Z(N338) );
  AO22D1BWP30P140LVT U543 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[221]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[221]), .Z(N339) );
  AO22D1BWP30P140LVT U544 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[222]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[222]), .Z(N340) );
  AO22D1BWP30P140LVT U545 ( .A1(n31), .A2(
        first_stage_output_def_1__o_data_bus_wire[223]), .B1(n30), .B2(
        first_stage_output_def_0__o_data_bus_wire[223]), .Z(N341) );
  IND2D1BWP30P140LVT U546 ( .A1(first_stage_output_def_0__o_valid_wire[7]), 
        .B1(first_stage_output_def_1__o_valid_wire[7]), .ZN(n49) );
  INVD2BWP30P140LVT U547 ( .I(n49), .ZN(n33) );
  IND2D1BWP30P140LVT U548 ( .A1(first_stage_output_def_1__o_valid_wire[7]), 
        .B1(first_stage_output_def_0__o_valid_wire[7]), .ZN(n48) );
  INVD2BWP30P140LVT U549 ( .I(n48), .ZN(n32) );
  AO22D1BWP30P140LVT U550 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[224]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[224]), .Z(N352) );
  AO22D1BWP30P140LVT U551 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[225]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[225]), .Z(N353) );
  AO22D1BWP30P140LVT U552 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[226]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[226]), .Z(N354) );
  AO22D1BWP30P140LVT U553 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[227]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[227]), .Z(N355) );
  AO22D1BWP30P140LVT U554 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[228]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[228]), .Z(N356) );
  AO22D1BWP30P140LVT U555 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[229]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[229]), .Z(N357) );
  AO22D1BWP30P140LVT U556 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[230]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[230]), .Z(N358) );
  AO22D1BWP30P140LVT U557 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[231]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[231]), .Z(N359) );
  AO22D1BWP30P140LVT U558 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[232]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[232]), .Z(N360) );
  AO22D1BWP30P140LVT U559 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[233]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[233]), .Z(N361) );
  AO22D1BWP30P140LVT U560 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[234]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[234]), .Z(N362) );
  AO22D1BWP30P140LVT U561 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[235]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[235]), .Z(N363) );
  AO22D1BWP30P140LVT U562 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[236]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[236]), .Z(N364) );
  AO22D1BWP30P140LVT U563 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[237]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[237]), .Z(N365) );
  AO22D1BWP30P140LVT U564 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[238]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[238]), .Z(N366) );
  AO22D1BWP30P140LVT U565 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[239]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[239]), .Z(N367) );
  AO22D1BWP30P140LVT U566 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[240]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[240]), .Z(N368) );
  AO22D1BWP30P140LVT U567 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[241]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[241]), .Z(N369) );
  AO22D1BWP30P140LVT U568 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[242]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[242]), .Z(N370) );
  AO22D1BWP30P140LVT U569 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[243]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[243]), .Z(N371) );
  AO22D1BWP30P140LVT U570 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[244]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[244]), .Z(N372) );
  AO22D1BWP30P140LVT U571 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[245]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[245]), .Z(N373) );
  AO22D1BWP30P140LVT U572 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[246]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[246]), .Z(N374) );
  AO22D1BWP30P140LVT U573 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[247]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[247]), .Z(N375) );
  AO22D1BWP30P140LVT U574 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[248]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[248]), .Z(N376) );
  AO22D1BWP30P140LVT U575 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[249]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[249]), .Z(N377) );
  AO22D1BWP30P140LVT U576 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[250]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[250]), .Z(N378) );
  AO22D1BWP30P140LVT U577 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[251]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[251]), .Z(N379) );
  AO22D1BWP30P140LVT U578 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[252]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[252]), .Z(N380) );
  AO22D1BWP30P140LVT U579 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[253]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[253]), .Z(N381) );
  AO22D1BWP30P140LVT U580 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[254]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[254]), .Z(N382) );
  AO22D1BWP30P140LVT U581 ( .A1(n33), .A2(
        first_stage_output_def_1__o_data_bus_wire[255]), .B1(n32), .B2(
        first_stage_output_def_0__o_data_bus_wire[255]), .Z(N383) );
endmodule

