

    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1, n2;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  CKBD1BWP30P140LVT U3 ( .I(n1), .Z(n2) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n2), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[119]), 
        .Z(N487) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[120]), 
        .Z(N488) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[122]), 
        .Z(N490) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[123]), 
        .Z(N491) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[125]), 
        .Z(N493) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[126]), 
        .Z(N494) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n2), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n2), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n2), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n2), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[29]), .Z(N32) );
  INR2D1BWP30P140LVT U137 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U268 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1, n2;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  CKBD1BWP30P140LVT U3 ( .I(n1), .Z(n2) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[119]), 
        .Z(N487) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[120]), 
        .Z(N488) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[122]), 
        .Z(N490) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[123]), 
        .Z(N491) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[125]), 
        .Z(N493) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[126]), 
        .Z(N494) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n2), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n2), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n2), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n2), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n2), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[29]), .Z(N32) );
  INR2D1BWP30P140LVT U137 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U268 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1, n2;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  CKBD1BWP30P140LVT U3 ( .I(n1), .Z(n2) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[119]), 
        .Z(N487) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[120]), 
        .Z(N488) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[122]), 
        .Z(N490) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[123]), 
        .Z(N491) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[125]), 
        .Z(N493) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[126]), 
        .Z(N494) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n2), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n2), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n2), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n2), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n2), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[29]), .Z(N32) );
  INR2D1BWP30P140LVT U137 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U268 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1, n2;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  CKBD1BWP30P140LVT U3 ( .I(n1), .Z(n2) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[119]), 
        .Z(N487) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[120]), 
        .Z(N488) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[122]), 
        .Z(N490) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[123]), 
        .Z(N491) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[125]), 
        .Z(N493) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[126]), 
        .Z(N494) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n2), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n2), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n2), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n2), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n2), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[29]), .Z(N32) );
  INR2D1BWP30P140LVT U137 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U268 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1, n2;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  CKBD1BWP30P140LVT U3 ( .I(n1), .Z(n2) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[119]), 
        .Z(N487) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[120]), 
        .Z(N488) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[122]), 
        .Z(N490) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[123]), 
        .Z(N491) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[125]), 
        .Z(N493) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[126]), 
        .Z(N494) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n2), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n2), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n2), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n2), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n2), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[29]), .Z(N32) );
  INR2D1BWP30P140LVT U137 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U268 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1, n2;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  CKBD1BWP30P140LVT U3 ( .I(n1), .Z(n2) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[119]), 
        .Z(N487) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[120]), 
        .Z(N488) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[122]), 
        .Z(N490) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[123]), 
        .Z(N491) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[125]), 
        .Z(N493) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[126]), 
        .Z(N494) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n2), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n2), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n2), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n2), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n2), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[29]), .Z(N32) );
  INR2D1BWP30P140LVT U137 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U268 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1, n2;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  CKBD1BWP30P140LVT U3 ( .I(n1), .Z(n2) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[119]), 
        .Z(N487) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[120]), 
        .Z(N488) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[122]), 
        .Z(N490) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[123]), 
        .Z(N491) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[125]), 
        .Z(N493) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[126]), 
        .Z(N494) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n2), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n2), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n2), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n2), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n2), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[29]), .Z(N32) );
  INR2D1BWP30P140LVT U137 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U268 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        clk, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input clk, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1, n2;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;

  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(clk), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(clk), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(clk), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(clk), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(clk), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(clk), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(clk), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(clk), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(clk), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(clk), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(clk), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(clk), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(clk), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(clk), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(clk), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(clk), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(clk), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(clk), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(clk), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(clk), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(clk), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(clk), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(clk), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(clk), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(clk), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(clk), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(clk), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(clk), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(clk), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(clk), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(clk), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(clk), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(clk), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(clk), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(clk), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(clk), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(clk), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(clk), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(clk), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(clk), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(clk), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(clk), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(clk), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(clk), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(clk), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(clk), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(clk), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(clk), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(clk), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(clk), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(clk), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(clk), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(clk), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(clk), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(clk), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(clk), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(clk), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        clk), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(clk), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(clk), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(clk), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(clk), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(clk), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(clk), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(clk), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(clk), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(clk), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(clk), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        clk), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        clk), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(clk), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(clk), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(clk), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(clk), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(clk), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(clk), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(clk), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(clk), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(clk), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(clk), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(clk), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(clk), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(clk), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(clk), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(clk), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(clk), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(clk), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(clk), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(clk), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(clk), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(clk), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(clk), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(clk), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(clk), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(clk), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(clk), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(clk), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(clk), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(clk), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(clk), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(clk), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(clk), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(clk), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(clk), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(clk), .Q(o_valid[6]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(clk), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(clk), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(clk), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(clk), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(clk), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(clk), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(clk), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(clk), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(clk), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(clk), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(clk), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(clk), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(clk), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(clk), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(clk), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(clk), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(clk), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(clk), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(clk), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(clk), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(clk), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(clk), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(clk), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(clk), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(clk), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(clk), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(clk), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(clk), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(clk), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(clk), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(clk), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(clk), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(clk), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(clk), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(clk), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(clk), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(clk), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(clk), .Q(
        o_data_bus[224]) );
  CKBD1BWP30P140LVT U3 ( .I(n1), .Z(n2) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n2), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[101]), 
        .Z(N469) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[102]), 
        .Z(N470) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[105]), 
        .Z(N473) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[107]), 
        .Z(N475) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[109]), 
        .Z(N477) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[110]), 
        .Z(N478) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[111]), 
        .Z(N479) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[112]), 
        .Z(N480) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[115]), 
        .Z(N483) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[119]), 
        .Z(N487) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[120]), 
        .Z(N488) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[122]), 
        .Z(N490) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[123]), 
        .Z(N491) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[125]), 
        .Z(N493) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[126]), 
        .Z(N494) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[64]), 
        .Z(N398) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[65]), 
        .Z(N399) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[68]), 
        .Z(N402) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[69]), 
        .Z(N403) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[70]), 
        .Z(N404) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[71]), 
        .Z(N405) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[72]), 
        .Z(N406) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[74]), 
        .Z(N408) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[75]), 
        .Z(N409) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[76]), 
        .Z(N410) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[78]), 
        .Z(N412) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[81]), 
        .Z(N415) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[83]), 
        .Z(N417) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[88]), 
        .Z(N422) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[93]), 
        .Z(N427) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[32]), 
        .Z(N332) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[34]), 
        .Z(N334) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[35]), 
        .Z(N335) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[39]), 
        .Z(N339) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[40]), 
        .Z(N340) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[42]), 
        .Z(N342) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[44]), 
        .Z(N344) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[45]), 
        .Z(N345) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[48]), 
        .Z(N348) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[49]), 
        .Z(N349) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[54]), 
        .Z(N354) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[55]), 
        .Z(N355) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[58]), 
        .Z(N358) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[59]), 
        .Z(N359) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[61]), 
        .Z(N361) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[7]), 
        .Z(N273) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[8]), 
        .Z(N274) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[9]), 
        .Z(N275) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[12]), 
        .Z(N278) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[13]), 
        .Z(N279) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[14]), 
        .Z(N280) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[15]), 
        .Z(N281) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[16]), 
        .Z(N282) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[17]), 
        .Z(N283) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[18]), 
        .Z(N284) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[19]), 
        .Z(N285) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[20]), 
        .Z(N286) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[21]), 
        .Z(N287) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[24]), 
        .Z(N290) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[26]), 
        .Z(N292) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[27]), 
        .Z(N293) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[29]), 
        .Z(N295) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n2), .A2(wire_tree_level_2__i_data_latch[30]), 
        .Z(N296) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n2), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n2), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n2), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n2), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n2), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n2), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n2), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n2), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U135 ( .A1(n2), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n2), .A2(i_data_bus[29]), .Z(N32) );
  INR2D1BWP30P140LVT U137 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[31]), 
        .Z(N297) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[28]), 
        .Z(N294) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[25]), 
        .Z(N291) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[23]), 
        .Z(N289) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[22]), 
        .Z(N288) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[11]), 
        .Z(N277) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[10]), 
        .Z(N276) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[5]), 
        .Z(N271) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[4]), 
        .Z(N270) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[3]), 
        .Z(N269) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[1]), 
        .Z(N267) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[0]), 
        .Z(N266) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[63]), 
        .Z(N363) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[62]), 
        .Z(N362) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[60]), 
        .Z(N360) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[57]), 
        .Z(N357) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[56]), 
        .Z(N356) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[53]), 
        .Z(N353) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[52]), 
        .Z(N352) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[51]), 
        .Z(N351) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[50]), 
        .Z(N350) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[47]), 
        .Z(N347) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[46]), 
        .Z(N346) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[43]), 
        .Z(N343) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[41]), 
        .Z(N341) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[38]), 
        .Z(N338) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[37]), 
        .Z(N337) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[36]), 
        .Z(N336) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[33]), 
        .Z(N333) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[95]), 
        .Z(N429) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[94]), 
        .Z(N428) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[92]), 
        .Z(N426) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[91]), 
        .Z(N425) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[90]), 
        .Z(N424) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[89]), 
        .Z(N423) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[87]), 
        .Z(N421) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[86]), 
        .Z(N420) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[85]), 
        .Z(N419) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[84]), 
        .Z(N418) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[82]), 
        .Z(N416) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[80]), 
        .Z(N414) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[79]), 
        .Z(N413) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[77]), 
        .Z(N411) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[73]), 
        .Z(N407) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[67]), 
        .Z(N401) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[66]), 
        .Z(N400) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(wire_tree_level_2__i_data_latch[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  CKAN2D1BWP30P140LVT U268 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        clk, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input clk, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(clk), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(clk), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        clk), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        clk), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        clk), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        clk), .Q(o_cmd_3) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        clk), .Q(o_cmd_4) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        clk), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        clk), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        clk), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule


module binary_tree_8_64_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, o_cmd, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [63:0] o_valid;
  output [2047:0] o_data_bus;
  output [63:0] o_cmd;
  input [63:0] i_cmd;
  input clk, rst, i_en;
  wire   n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352;

  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 top_half_0__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[0]), .i_data_bus(
        i_data_bus[31:0]), .o_valid({n2184, n2192, n2200, n2208, n2216, n2224, 
        n2232, n2240}), .o_data_bus({n2465, n2466, n2467, n2468, n2469, n2470, 
        n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
        n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2721, n2722, n2723, n2724, 
        n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, 
        n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, 
        n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2977, n2978, 
        n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
        n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
        n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
        n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
        n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
        n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
        n3263, n3264, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
        n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
        n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
        n3517, n3518, n3519, n3520, n3745, n3746, n3747, n3748, n3749, n3750, 
        n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, 
        n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, 
        n3771, n3772, n3773, n3774, n3775, n3776, n4001, n4002, n4003, n4004, 
        n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, 
        n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, 
        n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4257, n4258, 
        n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, 
        n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, 
        n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288}), 
        .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 top_half_1__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[1]), .i_data_bus(
        i_data_bus[63:32]), .o_valid({n2183, n2191, n2199, n2207, n2215, n2223, 
        n2231, n2239}), .o_data_bus({n2433, n2434, n2435, n2436, n2437, n2438, 
        n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, 
        n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, 
        n2459, n2460, n2461, n2462, n2463, n2464, n2689, n2690, n2691, n2692, 
        n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
        n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, 
        n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2945, n2946, 
        n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
        n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
        n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
        n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, 
        n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, 
        n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
        n3231, n3232, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, 
        n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, 
        n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, 
        n3485, n3486, n3487, n3488, n3713, n3714, n3715, n3716, n3717, n3718, 
        n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, 
        n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, 
        n3739, n3740, n3741, n3742, n3743, n3744, n3969, n3970, n3971, n3972, 
        n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
        n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
        n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4225, n4226, 
        n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, 
        n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, 
        n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256}), 
        .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 top_half_2__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[2]), .i_data_bus(
        i_data_bus[95:64]), .o_valid({n2182, n2190, n2198, n2206, n2214, n2222, 
        n2230, n2238}), .o_data_bus({n2401, n2402, n2403, n2404, n2405, n2406, 
        n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
        n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
        n2427, n2428, n2429, n2430, n2431, n2432, n2657, n2658, n2659, n2660, 
        n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, 
        n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, 
        n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2913, n2914, 
        n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, 
        n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, 
        n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, 
        n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, 
        n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
        n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
        n3199, n3200, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
        n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
        n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
        n3453, n3454, n3455, n3456, n3681, n3682, n3683, n3684, n3685, n3686, 
        n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, 
        n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, 
        n3707, n3708, n3709, n3710, n3711, n3712, n3937, n3938, n3939, n3940, 
        n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, 
        n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, 
        n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n4193, n4194, 
        n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, 
        n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, 
        n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224}), 
        .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 top_half_3__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[3]), .i_data_bus(
        i_data_bus[127:96]), .o_valid({n2181, n2189, n2197, n2205, n2213, 
        n2221, n2229, n2237}), .o_data_bus({n2369, n2370, n2371, n2372, n2373, 
        n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, 
        n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
        n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2625, n2626, n2627, 
        n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
        n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, 
        n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2881, 
        n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
        n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
        n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, 
        n2912, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, 
        n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, 
        n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, 
        n3166, n3167, n3168, n3393, n3394, n3395, n3396, n3397, n3398, n3399, 
        n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, 
        n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, 
        n3420, n3421, n3422, n3423, n3424, n3649, n3650, n3651, n3652, n3653, 
        n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, 
        n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
        n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3905, n3906, n3907, 
        n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, 
        n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, 
        n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n4161, 
        n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, 
        n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, 
        n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, 
        n4192}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 top_half_4__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[4]), .i_data_bus(
        i_data_bus[159:128]), .o_valid({n2180, n2188, n2196, n2204, n2212, 
        n2220, n2228, n2236}), .o_data_bus({n2337, n2338, n2339, n2340, n2341, 
        n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, 
        n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, 
        n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2593, n2594, n2595, 
        n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, 
        n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, 
        n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2849, 
        n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
        n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, 
        n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, 
        n2880, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
        n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
        n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
        n3134, n3135, n3136, n3361, n3362, n3363, n3364, n3365, n3366, n3367, 
        n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, 
        n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, 
        n3388, n3389, n3390, n3391, n3392, n3617, n3618, n3619, n3620, n3621, 
        n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, 
        n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, 
        n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3873, n3874, n3875, 
        n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, 
        n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, 
        n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n4129, 
        n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, 
        n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, 
        n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, 
        n4160}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 top_half_5__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[5]), .i_data_bus(
        i_data_bus[191:160]), .o_valid({n2179, n2187, n2195, n2203, n2211, 
        n2219, n2227, n2235}), .o_data_bus({n2305, n2306, n2307, n2308, n2309, 
        n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
        n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, 
        n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2561, n2562, n2563, 
        n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, 
        n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, 
        n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2817, 
        n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, 
        n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, 
        n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, 
        n2848, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
        n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
        n3102, n3103, n3104, n3329, n3330, n3331, n3332, n3333, n3334, n3335, 
        n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, 
        n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, 
        n3356, n3357, n3358, n3359, n3360, n3585, n3586, n3587, n3588, n3589, 
        n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, 
        n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, 
        n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3841, n3842, n3843, 
        n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, 
        n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, 
        n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n4097, 
        n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, 
        n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
        n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
        n4128}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 top_half_6__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[6]), .i_data_bus(
        i_data_bus[223:192]), .o_valid({n2178, n2186, n2194, n2202, n2210, 
        n2218, n2226, n2234}), .o_data_bus({n2273, n2274, n2275, n2276, n2277, 
        n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
        n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
        n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2529, n2530, n2531, 
        n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, 
        n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, 
        n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2785, 
        n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, 
        n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, 
        n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
        n2816, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, 
        n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, 
        n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, 
        n3070, n3071, n3072, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
        n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
        n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, 
        n3324, n3325, n3326, n3327, n3328, n3553, n3554, n3555, n3556, n3557, 
        n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, 
        n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, 
        n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3809, n3810, n3811, 
        n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, 
        n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, 
        n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n4065, 
        n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, 
        n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, 
        n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, 
        n4096}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 top_half_7__wire_pipeline ( 
        .clk(clk), .rst(rst), .i_valid(i_valid[7]), .i_data_bus(
        i_data_bus[255:224]), .o_valid({n2177, n2185, n2193, n2201, n2209, 
        n2217, n2225, n2233}), .o_data_bus({n2241, n2242, n2243, n2244, n2245, 
        n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, 
        n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, 
        n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2497, n2498, n2499, 
        n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, 
        n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
        n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2753, 
        n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, 
        n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, 
        n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
        n2784, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
        n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, 
        n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, 
        n3038, n3039, n3040, n3265, n3266, n3267, n3268, n3269, n3270, n3271, 
        n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
        n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, 
        n3292, n3293, n3294, n3295, n3296, n3521, n3522, n3523, n3524, n3525, 
        n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, 
        n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, 
        n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3777, n3778, n3779, 
        n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, 
        n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, 
        n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n4033, 
        n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, 
        n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, 
        n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, 
        n4064}), .i_en(i_en) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 i_cmd_id_0__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(n4352), .o_cmd_1(n4344), .o_cmd_2(n4336), .o_cmd_3(n4328), .o_cmd_4(n4320), .o_cmd_5(n4312), .o_cmd_6(n4304), 
        .o_cmd_7(n4296), .i_en(i_en), .i_cmd(i_cmd[7:0]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 i_cmd_id_1__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(n4351), .o_cmd_1(n4343), .o_cmd_2(n4335), .o_cmd_3(n4327), .o_cmd_4(n4319), .o_cmd_5(n4311), .o_cmd_6(n4303), 
        .o_cmd_7(n4295), .i_en(i_en), .i_cmd(i_cmd[15:8]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 i_cmd_id_2__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(n4350), .o_cmd_1(n4342), .o_cmd_2(n4334), .o_cmd_3(n4326), .o_cmd_4(n4318), .o_cmd_5(n4310), .o_cmd_6(n4302), 
        .o_cmd_7(n4294), .i_en(i_en), .i_cmd(i_cmd[23:16]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 i_cmd_id_3__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(n4349), .o_cmd_1(n4341), .o_cmd_2(n4333), .o_cmd_3(n4325), .o_cmd_4(n4317), .o_cmd_5(n4309), .o_cmd_6(n4301), 
        .o_cmd_7(n4293), .i_en(i_en), .i_cmd(i_cmd[31:24]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 i_cmd_id_4__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(n4348), .o_cmd_1(n4340), .o_cmd_2(n4332), .o_cmd_3(n4324), .o_cmd_4(n4316), .o_cmd_5(n4308), .o_cmd_6(n4300), 
        .o_cmd_7(n4292), .i_en(i_en), .i_cmd(i_cmd[39:32]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 i_cmd_id_5__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(n4347), .o_cmd_1(n4339), .o_cmd_2(n4331), .o_cmd_3(n4323), .o_cmd_4(n4315), .o_cmd_5(n4307), .o_cmd_6(n4299), 
        .o_cmd_7(n4291), .i_en(i_en), .i_cmd(i_cmd[47:40]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 i_cmd_id_6__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(n4346), .o_cmd_1(n4338), .o_cmd_2(n4330), .o_cmd_3(n4322), .o_cmd_4(n4314), .o_cmd_5(n4306), .o_cmd_6(n4298), 
        .o_cmd_7(n4290), .i_en(i_en), .i_cmd(i_cmd[55:48]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 i_cmd_id_7__cmd_pipeline ( 
        .clk(clk), .rst(rst), .o_cmd_0(n4345), .o_cmd_1(n4337), .o_cmd_2(n4329), .o_cmd_3(n4321), .o_cmd_4(n4313), .o_cmd_5(n4305), .o_cmd_6(n4297), 
        .o_cmd_7(n4289), .i_en(i_en), .i_cmd(i_cmd[63:56]) );
  BUFFD6BWP30P140LVT U1 ( .I(n2923), .Z(o_data_bus[1365]) );
  BUFFD6BWP30P140LVT U2 ( .I(n2991), .Z(o_data_bus[1297]) );
  BUFFD6BWP30P140LVT U3 ( .I(n2920), .Z(o_data_bus[1368]) );
  BUFFD6BWP30P140LVT U4 ( .I(n2921), .Z(o_data_bus[1367]) );
  BUFFD6BWP30P140LVT U5 ( .I(n2918), .Z(o_data_bus[1370]) );
  BUFFD6BWP30P140LVT U6 ( .I(n2919), .Z(o_data_bus[1369]) );
  BUFFD6BWP30P140LVT U7 ( .I(n2916), .Z(o_data_bus[1372]) );
  BUFFD6BWP30P140LVT U8 ( .I(n2915), .Z(o_data_bus[1373]) );
  BUFFD6BWP30P140LVT U9 ( .I(n2914), .Z(o_data_bus[1374]) );
  BUFFD6BWP30P140LVT U10 ( .I(n2913), .Z(o_data_bus[1375]) );
  BUFFD6BWP30P140LVT U11 ( .I(n2912), .Z(o_data_bus[1376]) );
  BUFFD6BWP30P140LVT U12 ( .I(n2911), .Z(o_data_bus[1377]) );
  BUFFD6BWP30P140LVT U13 ( .I(n2910), .Z(o_data_bus[1378]) );
  BUFFD6BWP30P140LVT U14 ( .I(n2909), .Z(o_data_bus[1379]) );
  BUFFD6BWP30P140LVT U15 ( .I(n2908), .Z(o_data_bus[1380]) );
  BUFFD6BWP30P140LVT U16 ( .I(n2907), .Z(o_data_bus[1381]) );
  BUFFD6BWP30P140LVT U17 ( .I(n2906), .Z(o_data_bus[1382]) );
  BUFFD6BWP30P140LVT U18 ( .I(n2905), .Z(o_data_bus[1383]) );
  BUFFD6BWP30P140LVT U19 ( .I(n2917), .Z(o_data_bus[1371]) );
  BUFFD6BWP30P140LVT U20 ( .I(n2904), .Z(o_data_bus[1384]) );
  BUFFD6BWP30P140LVT U21 ( .I(n2903), .Z(o_data_bus[1385]) );
  BUFFD6BWP30P140LVT U22 ( .I(n2902), .Z(o_data_bus[1386]) );
  BUFFD6BWP30P140LVT U23 ( .I(n2901), .Z(o_data_bus[1387]) );
  BUFFD6BWP30P140LVT U24 ( .I(n2900), .Z(o_data_bus[1388]) );
  BUFFD6BWP30P140LVT U25 ( .I(n2899), .Z(o_data_bus[1389]) );
  BUFFD6BWP30P140LVT U26 ( .I(n2898), .Z(o_data_bus[1390]) );
  BUFFD6BWP30P140LVT U27 ( .I(n2897), .Z(o_data_bus[1391]) );
  BUFFD6BWP30P140LVT U28 ( .I(n2896), .Z(o_data_bus[1392]) );
  BUFFD6BWP30P140LVT U29 ( .I(n2895), .Z(o_data_bus[1393]) );
  BUFFD6BWP30P140LVT U30 ( .I(n2922), .Z(o_data_bus[1366]) );
  BUFFD6BWP30P140LVT U31 ( .I(n2894), .Z(o_data_bus[1394]) );
  BUFFD6BWP30P140LVT U32 ( .I(n2893), .Z(o_data_bus[1395]) );
  BUFFD6BWP30P140LVT U33 ( .I(n2892), .Z(o_data_bus[1396]) );
  BUFFD6BWP30P140LVT U34 ( .I(n2924), .Z(o_data_bus[1364]) );
  BUFFD6BWP30P140LVT U35 ( .I(n2891), .Z(o_data_bus[1397]) );
  BUFFD6BWP30P140LVT U36 ( .I(n2890), .Z(o_data_bus[1398]) );
  BUFFD6BWP30P140LVT U37 ( .I(n2888), .Z(o_data_bus[1400]) );
  BUFFD6BWP30P140LVT U38 ( .I(n2887), .Z(o_data_bus[1401]) );
  BUFFD6BWP30P140LVT U39 ( .I(n2886), .Z(o_data_bus[1402]) );
  BUFFD6BWP30P140LVT U40 ( .I(n2885), .Z(o_data_bus[1403]) );
  BUFFD6BWP30P140LVT U41 ( .I(n2884), .Z(o_data_bus[1404]) );
  BUFFD6BWP30P140LVT U42 ( .I(n2883), .Z(o_data_bus[1405]) );
  BUFFD6BWP30P140LVT U43 ( .I(n2882), .Z(o_data_bus[1406]) );
  BUFFD6BWP30P140LVT U44 ( .I(n2881), .Z(o_data_bus[1407]) );
  BUFFD6BWP30P140LVT U45 ( .I(n2880), .Z(o_data_bus[1408]) );
  BUFFD6BWP30P140LVT U46 ( .I(n2879), .Z(o_data_bus[1409]) );
  BUFFD6BWP30P140LVT U47 ( .I(n2878), .Z(o_data_bus[1410]) );
  BUFFD6BWP30P140LVT U48 ( .I(n2877), .Z(o_data_bus[1411]) );
  BUFFD6BWP30P140LVT U49 ( .I(n2876), .Z(o_data_bus[1412]) );
  BUFFD6BWP30P140LVT U50 ( .I(n2875), .Z(o_data_bus[1413]) );
  BUFFD6BWP30P140LVT U51 ( .I(n2874), .Z(o_data_bus[1414]) );
  BUFFD6BWP30P140LVT U52 ( .I(n2873), .Z(o_data_bus[1415]) );
  BUFFD6BWP30P140LVT U53 ( .I(n2872), .Z(o_data_bus[1416]) );
  BUFFD6BWP30P140LVT U54 ( .I(n2871), .Z(o_data_bus[1417]) );
  BUFFD6BWP30P140LVT U55 ( .I(n2870), .Z(o_data_bus[1418]) );
  BUFFD6BWP30P140LVT U56 ( .I(n2869), .Z(o_data_bus[1419]) );
  BUFFD6BWP30P140LVT U57 ( .I(n2868), .Z(o_data_bus[1420]) );
  BUFFD6BWP30P140LVT U58 ( .I(n2867), .Z(o_data_bus[1421]) );
  BUFFD6BWP30P140LVT U59 ( .I(n2866), .Z(o_data_bus[1422]) );
  BUFFD6BWP30P140LVT U60 ( .I(n2865), .Z(o_data_bus[1423]) );
  BUFFD6BWP30P140LVT U61 ( .I(n2864), .Z(o_data_bus[1424]) );
  BUFFD6BWP30P140LVT U62 ( .I(n2863), .Z(o_data_bus[1425]) );
  BUFFD6BWP30P140LVT U63 ( .I(n2862), .Z(o_data_bus[1426]) );
  BUFFD6BWP30P140LVT U64 ( .I(n2861), .Z(o_data_bus[1427]) );
  BUFFD6BWP30P140LVT U65 ( .I(n2860), .Z(o_data_bus[1428]) );
  BUFFD6BWP30P140LVT U66 ( .I(n2859), .Z(o_data_bus[1429]) );
  BUFFD6BWP30P140LVT U67 ( .I(n2858), .Z(o_data_bus[1430]) );
  BUFFD6BWP30P140LVT U68 ( .I(n2925), .Z(o_data_bus[1363]) );
  BUFFD6BWP30P140LVT U69 ( .I(n2926), .Z(o_data_bus[1362]) );
  BUFFD6BWP30P140LVT U70 ( .I(n2927), .Z(o_data_bus[1361]) );
  BUFFD6BWP30P140LVT U71 ( .I(n2928), .Z(o_data_bus[1360]) );
  BUFFD6BWP30P140LVT U72 ( .I(n2929), .Z(o_data_bus[1359]) );
  BUFFD6BWP30P140LVT U73 ( .I(n2930), .Z(o_data_bus[1358]) );
  BUFFD6BWP30P140LVT U74 ( .I(n2931), .Z(o_data_bus[1357]) );
  BUFFD6BWP30P140LVT U75 ( .I(n2932), .Z(o_data_bus[1356]) );
  BUFFD6BWP30P140LVT U76 ( .I(n2933), .Z(o_data_bus[1355]) );
  BUFFD6BWP30P140LVT U77 ( .I(n2934), .Z(o_data_bus[1354]) );
  BUFFD6BWP30P140LVT U78 ( .I(n2935), .Z(o_data_bus[1353]) );
  BUFFD6BWP30P140LVT U79 ( .I(n2936), .Z(o_data_bus[1352]) );
  BUFFD6BWP30P140LVT U80 ( .I(n2937), .Z(o_data_bus[1351]) );
  BUFFD6BWP30P140LVT U81 ( .I(n2938), .Z(o_data_bus[1350]) );
  BUFFD6BWP30P140LVT U82 ( .I(n2939), .Z(o_data_bus[1349]) );
  BUFFD6BWP30P140LVT U83 ( .I(n2940), .Z(o_data_bus[1348]) );
  BUFFD6BWP30P140LVT U84 ( .I(n2941), .Z(o_data_bus[1347]) );
  BUFFD6BWP30P140LVT U85 ( .I(n2942), .Z(o_data_bus[1346]) );
  BUFFD6BWP30P140LVT U86 ( .I(n2943), .Z(o_data_bus[1345]) );
  BUFFD6BWP30P140LVT U87 ( .I(n2944), .Z(o_data_bus[1344]) );
  BUFFD6BWP30P140LVT U88 ( .I(n2945), .Z(o_data_bus[1343]) );
  BUFFD6BWP30P140LVT U89 ( .I(n2946), .Z(o_data_bus[1342]) );
  BUFFD6BWP30P140LVT U90 ( .I(n2947), .Z(o_data_bus[1341]) );
  BUFFD6BWP30P140LVT U91 ( .I(n2948), .Z(o_data_bus[1340]) );
  BUFFD6BWP30P140LVT U92 ( .I(n2949), .Z(o_data_bus[1339]) );
  BUFFD6BWP30P140LVT U93 ( .I(n2950), .Z(o_data_bus[1338]) );
  BUFFD6BWP30P140LVT U94 ( .I(n2951), .Z(o_data_bus[1337]) );
  BUFFD6BWP30P140LVT U95 ( .I(n2952), .Z(o_data_bus[1336]) );
  BUFFD6BWP30P140LVT U96 ( .I(n2953), .Z(o_data_bus[1335]) );
  BUFFD6BWP30P140LVT U97 ( .I(n2954), .Z(o_data_bus[1334]) );
  BUFFD6BWP30P140LVT U98 ( .I(n2955), .Z(o_data_bus[1333]) );
  BUFFD6BWP30P140LVT U99 ( .I(n2956), .Z(o_data_bus[1332]) );
  BUFFD6BWP30P140LVT U100 ( .I(n2957), .Z(o_data_bus[1331]) );
  BUFFD6BWP30P140LVT U101 ( .I(n2958), .Z(o_data_bus[1330]) );
  BUFFD6BWP30P140LVT U102 ( .I(n2959), .Z(o_data_bus[1329]) );
  BUFFD6BWP30P140LVT U103 ( .I(n2960), .Z(o_data_bus[1328]) );
  BUFFD6BWP30P140LVT U104 ( .I(n2961), .Z(o_data_bus[1327]) );
  BUFFD6BWP30P140LVT U105 ( .I(n2962), .Z(o_data_bus[1326]) );
  BUFFD6BWP30P140LVT U106 ( .I(n2963), .Z(o_data_bus[1325]) );
  BUFFD6BWP30P140LVT U107 ( .I(n2964), .Z(o_data_bus[1324]) );
  BUFFD6BWP30P140LVT U108 ( .I(n2965), .Z(o_data_bus[1323]) );
  BUFFD6BWP30P140LVT U109 ( .I(n2966), .Z(o_data_bus[1322]) );
  BUFFD6BWP30P140LVT U110 ( .I(n2967), .Z(o_data_bus[1321]) );
  BUFFD6BWP30P140LVT U111 ( .I(n2968), .Z(o_data_bus[1320]) );
  BUFFD6BWP30P140LVT U112 ( .I(n2969), .Z(o_data_bus[1319]) );
  BUFFD6BWP30P140LVT U113 ( .I(n2970), .Z(o_data_bus[1318]) );
  BUFFD6BWP30P140LVT U114 ( .I(n2971), .Z(o_data_bus[1317]) );
  BUFFD6BWP30P140LVT U115 ( .I(n2972), .Z(o_data_bus[1316]) );
  BUFFD6BWP30P140LVT U116 ( .I(n2973), .Z(o_data_bus[1315]) );
  BUFFD6BWP30P140LVT U117 ( .I(n2974), .Z(o_data_bus[1314]) );
  BUFFD6BWP30P140LVT U118 ( .I(n2975), .Z(o_data_bus[1313]) );
  BUFFD6BWP30P140LVT U119 ( .I(n2976), .Z(o_data_bus[1312]) );
  BUFFD6BWP30P140LVT U120 ( .I(n2977), .Z(o_data_bus[1311]) );
  BUFFD6BWP30P140LVT U121 ( .I(n2978), .Z(o_data_bus[1310]) );
  BUFFD6BWP30P140LVT U122 ( .I(n2979), .Z(o_data_bus[1309]) );
  BUFFD6BWP30P140LVT U123 ( .I(n2980), .Z(o_data_bus[1308]) );
  BUFFD6BWP30P140LVT U124 ( .I(n2981), .Z(o_data_bus[1307]) );
  BUFFD6BWP30P140LVT U125 ( .I(n2982), .Z(o_data_bus[1306]) );
  BUFFD6BWP30P140LVT U126 ( .I(n2983), .Z(o_data_bus[1305]) );
  BUFFD6BWP30P140LVT U127 ( .I(n2984), .Z(o_data_bus[1304]) );
  BUFFD6BWP30P140LVT U128 ( .I(n2985), .Z(o_data_bus[1303]) );
  BUFFD6BWP30P140LVT U129 ( .I(n2986), .Z(o_data_bus[1302]) );
  BUFFD6BWP30P140LVT U130 ( .I(n2987), .Z(o_data_bus[1301]) );
  BUFFD6BWP30P140LVT U131 ( .I(n2988), .Z(o_data_bus[1300]) );
  BUFFD6BWP30P140LVT U132 ( .I(n2989), .Z(o_data_bus[1299]) );
  BUFFD6BWP30P140LVT U133 ( .I(n2990), .Z(o_data_bus[1298]) );
  BUFFD6BWP30P140LVT U134 ( .I(n2721), .Z(o_data_bus[1567]) );
  BUFFD6BWP30P140LVT U135 ( .I(n2857), .Z(o_data_bus[1431]) );
  BUFFD6BWP30P140LVT U136 ( .I(n2723), .Z(o_data_bus[1565]) );
  BUFFD6BWP30P140LVT U137 ( .I(n2724), .Z(o_data_bus[1564]) );
  BUFFD6BWP30P140LVT U138 ( .I(n2725), .Z(o_data_bus[1563]) );
  BUFFD6BWP30P140LVT U139 ( .I(n2726), .Z(o_data_bus[1562]) );
  BUFFD6BWP30P140LVT U140 ( .I(n2727), .Z(o_data_bus[1561]) );
  BUFFD6BWP30P140LVT U141 ( .I(n2728), .Z(o_data_bus[1560]) );
  BUFFD6BWP30P140LVT U142 ( .I(n2729), .Z(o_data_bus[1559]) );
  BUFFD6BWP30P140LVT U143 ( .I(n2730), .Z(o_data_bus[1558]) );
  BUFFD6BWP30P140LVT U144 ( .I(n2731), .Z(o_data_bus[1557]) );
  BUFFD6BWP30P140LVT U145 ( .I(n2732), .Z(o_data_bus[1556]) );
  BUFFD6BWP30P140LVT U146 ( .I(n2733), .Z(o_data_bus[1555]) );
  BUFFD6BWP30P140LVT U147 ( .I(n2734), .Z(o_data_bus[1554]) );
  BUFFD6BWP30P140LVT U148 ( .I(n2735), .Z(o_data_bus[1553]) );
  BUFFD6BWP30P140LVT U149 ( .I(n2736), .Z(o_data_bus[1552]) );
  BUFFD6BWP30P140LVT U150 ( .I(n2737), .Z(o_data_bus[1551]) );
  BUFFD6BWP30P140LVT U151 ( .I(n2738), .Z(o_data_bus[1550]) );
  BUFFD6BWP30P140LVT U152 ( .I(n2739), .Z(o_data_bus[1549]) );
  BUFFD6BWP30P140LVT U153 ( .I(n2740), .Z(o_data_bus[1548]) );
  BUFFD6BWP30P140LVT U154 ( .I(n2741), .Z(o_data_bus[1547]) );
  BUFFD6BWP30P140LVT U155 ( .I(n2742), .Z(o_data_bus[1546]) );
  BUFFD6BWP30P140LVT U156 ( .I(n2743), .Z(o_data_bus[1545]) );
  BUFFD6BWP30P140LVT U157 ( .I(n2744), .Z(o_data_bus[1544]) );
  BUFFD6BWP30P140LVT U158 ( .I(n2745), .Z(o_data_bus[1543]) );
  BUFFD6BWP30P140LVT U159 ( .I(n2746), .Z(o_data_bus[1542]) );
  BUFFD6BWP30P140LVT U160 ( .I(n2747), .Z(o_data_bus[1541]) );
  BUFFD6BWP30P140LVT U161 ( .I(n2748), .Z(o_data_bus[1540]) );
  BUFFD6BWP30P140LVT U162 ( .I(n2749), .Z(o_data_bus[1539]) );
  BUFFD6BWP30P140LVT U163 ( .I(n2750), .Z(o_data_bus[1538]) );
  BUFFD6BWP30P140LVT U164 ( .I(n2751), .Z(o_data_bus[1537]) );
  BUFFD6BWP30P140LVT U165 ( .I(n2752), .Z(o_data_bus[1536]) );
  BUFFD6BWP30P140LVT U166 ( .I(n2753), .Z(o_data_bus[1535]) );
  BUFFD6BWP30P140LVT U167 ( .I(n2754), .Z(o_data_bus[1534]) );
  BUFFD6BWP30P140LVT U168 ( .I(n2755), .Z(o_data_bus[1533]) );
  BUFFD6BWP30P140LVT U169 ( .I(n2756), .Z(o_data_bus[1532]) );
  BUFFD6BWP30P140LVT U170 ( .I(n2757), .Z(o_data_bus[1531]) );
  BUFFD6BWP30P140LVT U171 ( .I(n2758), .Z(o_data_bus[1530]) );
  BUFFD6BWP30P140LVT U172 ( .I(n2759), .Z(o_data_bus[1529]) );
  BUFFD6BWP30P140LVT U173 ( .I(n2760), .Z(o_data_bus[1528]) );
  BUFFD6BWP30P140LVT U174 ( .I(n2761), .Z(o_data_bus[1527]) );
  BUFFD6BWP30P140LVT U175 ( .I(n2762), .Z(o_data_bus[1526]) );
  BUFFD6BWP30P140LVT U176 ( .I(n2763), .Z(o_data_bus[1525]) );
  BUFFD6BWP30P140LVT U177 ( .I(n2764), .Z(o_data_bus[1524]) );
  BUFFD6BWP30P140LVT U178 ( .I(n2765), .Z(o_data_bus[1523]) );
  BUFFD6BWP30P140LVT U179 ( .I(n2766), .Z(o_data_bus[1522]) );
  BUFFD6BWP30P140LVT U180 ( .I(n2767), .Z(o_data_bus[1521]) );
  BUFFD6BWP30P140LVT U181 ( .I(n2768), .Z(o_data_bus[1520]) );
  BUFFD6BWP30P140LVT U182 ( .I(n2769), .Z(o_data_bus[1519]) );
  BUFFD6BWP30P140LVT U183 ( .I(n2770), .Z(o_data_bus[1518]) );
  BUFFD6BWP30P140LVT U184 ( .I(n2771), .Z(o_data_bus[1517]) );
  BUFFD6BWP30P140LVT U185 ( .I(n2772), .Z(o_data_bus[1516]) );
  BUFFD6BWP30P140LVT U186 ( .I(n2773), .Z(o_data_bus[1515]) );
  BUFFD6BWP30P140LVT U187 ( .I(n2774), .Z(o_data_bus[1514]) );
  BUFFD6BWP30P140LVT U188 ( .I(n2775), .Z(o_data_bus[1513]) );
  BUFFD6BWP30P140LVT U189 ( .I(n2776), .Z(o_data_bus[1512]) );
  BUFFD6BWP30P140LVT U190 ( .I(n2777), .Z(o_data_bus[1511]) );
  BUFFD6BWP30P140LVT U191 ( .I(n2778), .Z(o_data_bus[1510]) );
  BUFFD6BWP30P140LVT U192 ( .I(n2779), .Z(o_data_bus[1509]) );
  BUFFD6BWP30P140LVT U193 ( .I(n2780), .Z(o_data_bus[1508]) );
  BUFFD6BWP30P140LVT U194 ( .I(n2781), .Z(o_data_bus[1507]) );
  BUFFD6BWP30P140LVT U195 ( .I(n2782), .Z(o_data_bus[1506]) );
  BUFFD6BWP30P140LVT U196 ( .I(n2783), .Z(o_data_bus[1505]) );
  BUFFD6BWP30P140LVT U197 ( .I(n2784), .Z(o_data_bus[1504]) );
  BUFFD6BWP30P140LVT U198 ( .I(n2785), .Z(o_data_bus[1503]) );
  BUFFD6BWP30P140LVT U199 ( .I(n2786), .Z(o_data_bus[1502]) );
  BUFFD6BWP30P140LVT U200 ( .I(n2787), .Z(o_data_bus[1501]) );
  BUFFD6BWP30P140LVT U201 ( .I(n2788), .Z(o_data_bus[1500]) );
  BUFFD6BWP30P140LVT U202 ( .I(n2789), .Z(o_data_bus[1499]) );
  BUFFD6BWP30P140LVT U203 ( .I(n2790), .Z(o_data_bus[1498]) );
  BUFFD6BWP30P140LVT U204 ( .I(n2722), .Z(o_data_bus[1566]) );
  BUFFD6BWP30P140LVT U205 ( .I(n2791), .Z(o_data_bus[1497]) );
  BUFFD6BWP30P140LVT U206 ( .I(n2792), .Z(o_data_bus[1496]) );
  BUFFD6BWP30P140LVT U207 ( .I(n2793), .Z(o_data_bus[1495]) );
  BUFFD6BWP30P140LVT U208 ( .I(n2794), .Z(o_data_bus[1494]) );
  BUFFD6BWP30P140LVT U209 ( .I(n2795), .Z(o_data_bus[1493]) );
  BUFFD6BWP30P140LVT U210 ( .I(n2796), .Z(o_data_bus[1492]) );
  BUFFD6BWP30P140LVT U211 ( .I(n2797), .Z(o_data_bus[1491]) );
  BUFFD6BWP30P140LVT U212 ( .I(n2798), .Z(o_data_bus[1490]) );
  BUFFD6BWP30P140LVT U213 ( .I(n2799), .Z(o_data_bus[1489]) );
  BUFFD6BWP30P140LVT U214 ( .I(n2800), .Z(o_data_bus[1488]) );
  BUFFD6BWP30P140LVT U215 ( .I(n2801), .Z(o_data_bus[1487]) );
  BUFFD6BWP30P140LVT U216 ( .I(n2802), .Z(o_data_bus[1486]) );
  BUFFD6BWP30P140LVT U217 ( .I(n2803), .Z(o_data_bus[1485]) );
  BUFFD6BWP30P140LVT U218 ( .I(n2804), .Z(o_data_bus[1484]) );
  BUFFD6BWP30P140LVT U219 ( .I(n2805), .Z(o_data_bus[1483]) );
  BUFFD6BWP30P140LVT U220 ( .I(n2806), .Z(o_data_bus[1482]) );
  BUFFD6BWP30P140LVT U221 ( .I(n2807), .Z(o_data_bus[1481]) );
  BUFFD6BWP30P140LVT U222 ( .I(n2808), .Z(o_data_bus[1480]) );
  BUFFD6BWP30P140LVT U223 ( .I(n2809), .Z(o_data_bus[1479]) );
  BUFFD6BWP30P140LVT U224 ( .I(n2810), .Z(o_data_bus[1478]) );
  BUFFD6BWP30P140LVT U225 ( .I(n2811), .Z(o_data_bus[1477]) );
  BUFFD6BWP30P140LVT U226 ( .I(n2812), .Z(o_data_bus[1476]) );
  BUFFD6BWP30P140LVT U227 ( .I(n2813), .Z(o_data_bus[1475]) );
  BUFFD6BWP30P140LVT U228 ( .I(n2814), .Z(o_data_bus[1474]) );
  BUFFD6BWP30P140LVT U229 ( .I(n2815), .Z(o_data_bus[1473]) );
  BUFFD6BWP30P140LVT U230 ( .I(n2816), .Z(o_data_bus[1472]) );
  BUFFD6BWP30P140LVT U231 ( .I(n2817), .Z(o_data_bus[1471]) );
  BUFFD6BWP30P140LVT U232 ( .I(n2818), .Z(o_data_bus[1470]) );
  BUFFD6BWP30P140LVT U233 ( .I(n2819), .Z(o_data_bus[1469]) );
  BUFFD6BWP30P140LVT U234 ( .I(n2820), .Z(o_data_bus[1468]) );
  BUFFD6BWP30P140LVT U235 ( .I(n2821), .Z(o_data_bus[1467]) );
  BUFFD6BWP30P140LVT U236 ( .I(n2822), .Z(o_data_bus[1466]) );
  BUFFD6BWP30P140LVT U237 ( .I(n2823), .Z(o_data_bus[1465]) );
  BUFFD6BWP30P140LVT U238 ( .I(n2824), .Z(o_data_bus[1464]) );
  BUFFD6BWP30P140LVT U239 ( .I(n2825), .Z(o_data_bus[1463]) );
  BUFFD6BWP30P140LVT U240 ( .I(n2826), .Z(o_data_bus[1462]) );
  BUFFD6BWP30P140LVT U241 ( .I(n2827), .Z(o_data_bus[1461]) );
  BUFFD6BWP30P140LVT U242 ( .I(n2828), .Z(o_data_bus[1460]) );
  BUFFD6BWP30P140LVT U243 ( .I(n2829), .Z(o_data_bus[1459]) );
  BUFFD6BWP30P140LVT U244 ( .I(n2830), .Z(o_data_bus[1458]) );
  BUFFD6BWP30P140LVT U245 ( .I(n2831), .Z(o_data_bus[1457]) );
  BUFFD6BWP30P140LVT U246 ( .I(n2832), .Z(o_data_bus[1456]) );
  BUFFD6BWP30P140LVT U247 ( .I(n2833), .Z(o_data_bus[1455]) );
  BUFFD6BWP30P140LVT U248 ( .I(n2834), .Z(o_data_bus[1454]) );
  BUFFD6BWP30P140LVT U249 ( .I(n2835), .Z(o_data_bus[1453]) );
  BUFFD6BWP30P140LVT U250 ( .I(n2836), .Z(o_data_bus[1452]) );
  BUFFD6BWP30P140LVT U251 ( .I(n2837), .Z(o_data_bus[1451]) );
  BUFFD6BWP30P140LVT U252 ( .I(n2838), .Z(o_data_bus[1450]) );
  BUFFD6BWP30P140LVT U253 ( .I(n2839), .Z(o_data_bus[1449]) );
  BUFFD6BWP30P140LVT U254 ( .I(n2840), .Z(o_data_bus[1448]) );
  BUFFD6BWP30P140LVT U255 ( .I(n2841), .Z(o_data_bus[1447]) );
  BUFFD6BWP30P140LVT U256 ( .I(n2842), .Z(o_data_bus[1446]) );
  BUFFD6BWP30P140LVT U257 ( .I(n2843), .Z(o_data_bus[1445]) );
  BUFFD6BWP30P140LVT U258 ( .I(n2844), .Z(o_data_bus[1444]) );
  BUFFD6BWP30P140LVT U259 ( .I(n2845), .Z(o_data_bus[1443]) );
  BUFFD6BWP30P140LVT U260 ( .I(n2846), .Z(o_data_bus[1442]) );
  BUFFD6BWP30P140LVT U261 ( .I(n2847), .Z(o_data_bus[1441]) );
  BUFFD6BWP30P140LVT U262 ( .I(n2848), .Z(o_data_bus[1440]) );
  BUFFD6BWP30P140LVT U263 ( .I(n2849), .Z(o_data_bus[1439]) );
  BUFFD6BWP30P140LVT U264 ( .I(n2850), .Z(o_data_bus[1438]) );
  BUFFD6BWP30P140LVT U265 ( .I(n2851), .Z(o_data_bus[1437]) );
  BUFFD6BWP30P140LVT U266 ( .I(n2852), .Z(o_data_bus[1436]) );
  BUFFD6BWP30P140LVT U267 ( .I(n2853), .Z(o_data_bus[1435]) );
  BUFFD6BWP30P140LVT U268 ( .I(n2854), .Z(o_data_bus[1434]) );
  BUFFD6BWP30P140LVT U269 ( .I(n2855), .Z(o_data_bus[1433]) );
  BUFFD6BWP30P140LVT U270 ( .I(n2856), .Z(o_data_bus[1432]) );
  BUFFD6BWP30P140LVT U271 ( .I(n2992), .Z(o_data_bus[1296]) );
  BUFFD6BWP30P140LVT U272 ( .I(n2889), .Z(o_data_bus[1399]) );
  BUFFD6BWP30P140LVT U273 ( .I(n3130), .Z(o_data_bus[1158]) );
  BUFFD6BWP30P140LVT U274 ( .I(n3131), .Z(o_data_bus[1157]) );
  BUFFD6BWP30P140LVT U275 ( .I(n3132), .Z(o_data_bus[1156]) );
  BUFFD6BWP30P140LVT U276 ( .I(n3133), .Z(o_data_bus[1155]) );
  BUFFD6BWP30P140LVT U277 ( .I(n3134), .Z(o_data_bus[1154]) );
  BUFFD6BWP30P140LVT U278 ( .I(n3135), .Z(o_data_bus[1153]) );
  BUFFD6BWP30P140LVT U279 ( .I(n3136), .Z(o_data_bus[1152]) );
  BUFFD6BWP30P140LVT U280 ( .I(n3137), .Z(o_data_bus[1151]) );
  BUFFD6BWP30P140LVT U281 ( .I(n3138), .Z(o_data_bus[1150]) );
  BUFFD6BWP30P140LVT U282 ( .I(n3139), .Z(o_data_bus[1149]) );
  BUFFD6BWP30P140LVT U283 ( .I(n3140), .Z(o_data_bus[1148]) );
  BUFFD6BWP30P140LVT U284 ( .I(n3141), .Z(o_data_bus[1147]) );
  BUFFD6BWP30P140LVT U285 ( .I(n3142), .Z(o_data_bus[1146]) );
  BUFFD6BWP30P140LVT U286 ( .I(n3143), .Z(o_data_bus[1145]) );
  BUFFD6BWP30P140LVT U287 ( .I(n3144), .Z(o_data_bus[1144]) );
  BUFFD6BWP30P140LVT U288 ( .I(n3145), .Z(o_data_bus[1143]) );
  BUFFD6BWP30P140LVT U289 ( .I(n3146), .Z(o_data_bus[1142]) );
  BUFFD6BWP30P140LVT U290 ( .I(n3147), .Z(o_data_bus[1141]) );
  BUFFD6BWP30P140LVT U291 ( .I(n3148), .Z(o_data_bus[1140]) );
  BUFFD6BWP30P140LVT U292 ( .I(n3149), .Z(o_data_bus[1139]) );
  BUFFD6BWP30P140LVT U293 ( .I(n3150), .Z(o_data_bus[1138]) );
  BUFFD6BWP30P140LVT U294 ( .I(n3151), .Z(o_data_bus[1137]) );
  BUFFD6BWP30P140LVT U295 ( .I(n3152), .Z(o_data_bus[1136]) );
  BUFFD6BWP30P140LVT U296 ( .I(n3153), .Z(o_data_bus[1135]) );
  BUFFD6BWP30P140LVT U297 ( .I(n3154), .Z(o_data_bus[1134]) );
  BUFFD6BWP30P140LVT U298 ( .I(n3155), .Z(o_data_bus[1133]) );
  BUFFD6BWP30P140LVT U299 ( .I(n3156), .Z(o_data_bus[1132]) );
  BUFFD6BWP30P140LVT U300 ( .I(n3157), .Z(o_data_bus[1131]) );
  BUFFD6BWP30P140LVT U301 ( .I(n3158), .Z(o_data_bus[1130]) );
  BUFFD6BWP30P140LVT U302 ( .I(n3159), .Z(o_data_bus[1129]) );
  BUFFD6BWP30P140LVT U303 ( .I(n3160), .Z(o_data_bus[1128]) );
  BUFFD6BWP30P140LVT U304 ( .I(n3161), .Z(o_data_bus[1127]) );
  BUFFD6BWP30P140LVT U305 ( .I(n3162), .Z(o_data_bus[1126]) );
  BUFFD6BWP30P140LVT U306 ( .I(n3163), .Z(o_data_bus[1125]) );
  BUFFD6BWP30P140LVT U307 ( .I(n3164), .Z(o_data_bus[1124]) );
  BUFFD6BWP30P140LVT U308 ( .I(n3165), .Z(o_data_bus[1123]) );
  BUFFD6BWP30P140LVT U309 ( .I(n3166), .Z(o_data_bus[1122]) );
  BUFFD6BWP30P140LVT U310 ( .I(n3167), .Z(o_data_bus[1121]) );
  BUFFD6BWP30P140LVT U311 ( .I(n3168), .Z(o_data_bus[1120]) );
  BUFFD6BWP30P140LVT U312 ( .I(n3169), .Z(o_data_bus[1119]) );
  BUFFD6BWP30P140LVT U313 ( .I(n3170), .Z(o_data_bus[1118]) );
  BUFFD6BWP30P140LVT U314 ( .I(n3171), .Z(o_data_bus[1117]) );
  BUFFD6BWP30P140LVT U315 ( .I(n3172), .Z(o_data_bus[1116]) );
  BUFFD6BWP30P140LVT U316 ( .I(n3173), .Z(o_data_bus[1115]) );
  BUFFD6BWP30P140LVT U317 ( .I(n3174), .Z(o_data_bus[1114]) );
  BUFFD6BWP30P140LVT U318 ( .I(n3175), .Z(o_data_bus[1113]) );
  BUFFD6BWP30P140LVT U319 ( .I(n3176), .Z(o_data_bus[1112]) );
  BUFFD6BWP30P140LVT U320 ( .I(n3177), .Z(o_data_bus[1111]) );
  BUFFD6BWP30P140LVT U321 ( .I(n3178), .Z(o_data_bus[1110]) );
  BUFFD6BWP30P140LVT U322 ( .I(n3179), .Z(o_data_bus[1109]) );
  BUFFD6BWP30P140LVT U323 ( .I(n3180), .Z(o_data_bus[1108]) );
  BUFFD6BWP30P140LVT U324 ( .I(n3181), .Z(o_data_bus[1107]) );
  BUFFD6BWP30P140LVT U325 ( .I(n3182), .Z(o_data_bus[1106]) );
  BUFFD6BWP30P140LVT U326 ( .I(n3183), .Z(o_data_bus[1105]) );
  BUFFD6BWP30P140LVT U327 ( .I(n3184), .Z(o_data_bus[1104]) );
  BUFFD6BWP30P140LVT U328 ( .I(n3185), .Z(o_data_bus[1103]) );
  BUFFD6BWP30P140LVT U329 ( .I(n3186), .Z(o_data_bus[1102]) );
  BUFFD6BWP30P140LVT U330 ( .I(n3187), .Z(o_data_bus[1101]) );
  BUFFD6BWP30P140LVT U331 ( .I(n3188), .Z(o_data_bus[1100]) );
  BUFFD6BWP30P140LVT U332 ( .I(n3189), .Z(o_data_bus[1099]) );
  BUFFD6BWP30P140LVT U333 ( .I(n3190), .Z(o_data_bus[1098]) );
  BUFFD6BWP30P140LVT U334 ( .I(n3191), .Z(o_data_bus[1097]) );
  BUFFD6BWP30P140LVT U335 ( .I(n3192), .Z(o_data_bus[1096]) );
  BUFFD6BWP30P140LVT U336 ( .I(n3193), .Z(o_data_bus[1095]) );
  BUFFD6BWP30P140LVT U337 ( .I(n3194), .Z(o_data_bus[1094]) );
  BUFFD6BWP30P140LVT U338 ( .I(n3195), .Z(o_data_bus[1093]) );
  BUFFD6BWP30P140LVT U339 ( .I(n3196), .Z(o_data_bus[1092]) );
  BUFFD6BWP30P140LVT U340 ( .I(n3129), .Z(o_data_bus[1159]) );
  BUFFD6BWP30P140LVT U341 ( .I(n3197), .Z(o_data_bus[1091]) );
  BUFFD6BWP30P140LVT U342 ( .I(n3198), .Z(o_data_bus[1090]) );
  BUFFD6BWP30P140LVT U343 ( .I(n3199), .Z(o_data_bus[1089]) );
  BUFFD6BWP30P140LVT U344 ( .I(n3200), .Z(o_data_bus[1088]) );
  BUFFD6BWP30P140LVT U345 ( .I(n3201), .Z(o_data_bus[1087]) );
  BUFFD6BWP30P140LVT U346 ( .I(n3202), .Z(o_data_bus[1086]) );
  BUFFD6BWP30P140LVT U347 ( .I(n3203), .Z(o_data_bus[1085]) );
  BUFFD6BWP30P140LVT U348 ( .I(n3204), .Z(o_data_bus[1084]) );
  BUFFD6BWP30P140LVT U349 ( .I(n3205), .Z(o_data_bus[1083]) );
  BUFFD6BWP30P140LVT U350 ( .I(n3206), .Z(o_data_bus[1082]) );
  BUFFD6BWP30P140LVT U351 ( .I(n3207), .Z(o_data_bus[1081]) );
  BUFFD6BWP30P140LVT U352 ( .I(n3208), .Z(o_data_bus[1080]) );
  BUFFD6BWP30P140LVT U353 ( .I(n3209), .Z(o_data_bus[1079]) );
  BUFFD6BWP30P140LVT U354 ( .I(n3210), .Z(o_data_bus[1078]) );
  BUFFD6BWP30P140LVT U355 ( .I(n3211), .Z(o_data_bus[1077]) );
  BUFFD6BWP30P140LVT U356 ( .I(n3212), .Z(o_data_bus[1076]) );
  BUFFD6BWP30P140LVT U357 ( .I(n3213), .Z(o_data_bus[1075]) );
  BUFFD6BWP30P140LVT U358 ( .I(n3214), .Z(o_data_bus[1074]) );
  BUFFD6BWP30P140LVT U359 ( .I(n3215), .Z(o_data_bus[1073]) );
  BUFFD6BWP30P140LVT U360 ( .I(n3216), .Z(o_data_bus[1072]) );
  BUFFD6BWP30P140LVT U361 ( .I(n3217), .Z(o_data_bus[1071]) );
  BUFFD6BWP30P140LVT U362 ( .I(n3218), .Z(o_data_bus[1070]) );
  BUFFD6BWP30P140LVT U363 ( .I(n3219), .Z(o_data_bus[1069]) );
  BUFFD6BWP30P140LVT U364 ( .I(n3220), .Z(o_data_bus[1068]) );
  BUFFD6BWP30P140LVT U365 ( .I(n3221), .Z(o_data_bus[1067]) );
  BUFFD6BWP30P140LVT U366 ( .I(n3222), .Z(o_data_bus[1066]) );
  BUFFD6BWP30P140LVT U367 ( .I(n3223), .Z(o_data_bus[1065]) );
  BUFFD6BWP30P140LVT U368 ( .I(n3224), .Z(o_data_bus[1064]) );
  BUFFD6BWP30P140LVT U369 ( .I(n3225), .Z(o_data_bus[1063]) );
  BUFFD6BWP30P140LVT U370 ( .I(n3226), .Z(o_data_bus[1062]) );
  BUFFD6BWP30P140LVT U371 ( .I(n3227), .Z(o_data_bus[1061]) );
  BUFFD6BWP30P140LVT U372 ( .I(n3228), .Z(o_data_bus[1060]) );
  BUFFD6BWP30P140LVT U373 ( .I(n3229), .Z(o_data_bus[1059]) );
  BUFFD6BWP30P140LVT U374 ( .I(n3230), .Z(o_data_bus[1058]) );
  BUFFD6BWP30P140LVT U375 ( .I(n3231), .Z(o_data_bus[1057]) );
  BUFFD6BWP30P140LVT U376 ( .I(n3232), .Z(o_data_bus[1056]) );
  BUFFD6BWP30P140LVT U377 ( .I(n3233), .Z(o_data_bus[1055]) );
  BUFFD6BWP30P140LVT U378 ( .I(n3234), .Z(o_data_bus[1054]) );
  BUFFD6BWP30P140LVT U379 ( .I(n3235), .Z(o_data_bus[1053]) );
  BUFFD6BWP30P140LVT U380 ( .I(n3236), .Z(o_data_bus[1052]) );
  BUFFD6BWP30P140LVT U381 ( .I(n3237), .Z(o_data_bus[1051]) );
  BUFFD6BWP30P140LVT U382 ( .I(n3238), .Z(o_data_bus[1050]) );
  BUFFD6BWP30P140LVT U383 ( .I(n3239), .Z(o_data_bus[1049]) );
  BUFFD6BWP30P140LVT U384 ( .I(n3240), .Z(o_data_bus[1048]) );
  BUFFD6BWP30P140LVT U385 ( .I(n3241), .Z(o_data_bus[1047]) );
  BUFFD6BWP30P140LVT U386 ( .I(n3242), .Z(o_data_bus[1046]) );
  BUFFD6BWP30P140LVT U387 ( .I(n3243), .Z(o_data_bus[1045]) );
  BUFFD6BWP30P140LVT U388 ( .I(n3244), .Z(o_data_bus[1044]) );
  BUFFD6BWP30P140LVT U389 ( .I(n3245), .Z(o_data_bus[1043]) );
  BUFFD6BWP30P140LVT U390 ( .I(n3246), .Z(o_data_bus[1042]) );
  BUFFD6BWP30P140LVT U391 ( .I(n3247), .Z(o_data_bus[1041]) );
  BUFFD6BWP30P140LVT U392 ( .I(n3248), .Z(o_data_bus[1040]) );
  BUFFD6BWP30P140LVT U393 ( .I(n3249), .Z(o_data_bus[1039]) );
  BUFFD6BWP30P140LVT U394 ( .I(n3250), .Z(o_data_bus[1038]) );
  BUFFD6BWP30P140LVT U395 ( .I(n3251), .Z(o_data_bus[1037]) );
  BUFFD6BWP30P140LVT U396 ( .I(n3252), .Z(o_data_bus[1036]) );
  BUFFD6BWP30P140LVT U397 ( .I(n3253), .Z(o_data_bus[1035]) );
  BUFFD6BWP30P140LVT U398 ( .I(n3254), .Z(o_data_bus[1034]) );
  BUFFD6BWP30P140LVT U399 ( .I(n3255), .Z(o_data_bus[1033]) );
  BUFFD6BWP30P140LVT U400 ( .I(n3256), .Z(o_data_bus[1032]) );
  BUFFD6BWP30P140LVT U401 ( .I(n3257), .Z(o_data_bus[1031]) );
  BUFFD6BWP30P140LVT U402 ( .I(n3258), .Z(o_data_bus[1030]) );
  BUFFD6BWP30P140LVT U403 ( .I(n3259), .Z(o_data_bus[1029]) );
  BUFFD6BWP30P140LVT U404 ( .I(n3260), .Z(o_data_bus[1028]) );
  BUFFD6BWP30P140LVT U405 ( .I(n3261), .Z(o_data_bus[1027]) );
  BUFFD6BWP30P140LVT U406 ( .I(n3262), .Z(o_data_bus[1026]) );
  BUFFD6BWP30P140LVT U407 ( .I(n3263), .Z(o_data_bus[1025]) );
  BUFFD6BWP30P140LVT U408 ( .I(n2994), .Z(o_data_bus[1294]) );
  BUFFD6BWP30P140LVT U409 ( .I(n2995), .Z(o_data_bus[1293]) );
  BUFFD6BWP30P140LVT U410 ( .I(n2996), .Z(o_data_bus[1292]) );
  BUFFD6BWP30P140LVT U411 ( .I(n2997), .Z(o_data_bus[1291]) );
  BUFFD6BWP30P140LVT U412 ( .I(n2998), .Z(o_data_bus[1290]) );
  BUFFD6BWP30P140LVT U413 ( .I(n2999), .Z(o_data_bus[1289]) );
  BUFFD6BWP30P140LVT U414 ( .I(n3000), .Z(o_data_bus[1288]) );
  BUFFD6BWP30P140LVT U415 ( .I(n3001), .Z(o_data_bus[1287]) );
  BUFFD6BWP30P140LVT U416 ( .I(n3002), .Z(o_data_bus[1286]) );
  BUFFD6BWP30P140LVT U417 ( .I(n3003), .Z(o_data_bus[1285]) );
  BUFFD6BWP30P140LVT U418 ( .I(n3004), .Z(o_data_bus[1284]) );
  BUFFD6BWP30P140LVT U419 ( .I(n3005), .Z(o_data_bus[1283]) );
  BUFFD6BWP30P140LVT U420 ( .I(n3006), .Z(o_data_bus[1282]) );
  BUFFD6BWP30P140LVT U421 ( .I(n3007), .Z(o_data_bus[1281]) );
  BUFFD6BWP30P140LVT U422 ( .I(n3008), .Z(o_data_bus[1280]) );
  BUFFD6BWP30P140LVT U423 ( .I(n3009), .Z(o_data_bus[1279]) );
  BUFFD6BWP30P140LVT U424 ( .I(n3010), .Z(o_data_bus[1278]) );
  BUFFD6BWP30P140LVT U425 ( .I(n3011), .Z(o_data_bus[1277]) );
  BUFFD6BWP30P140LVT U426 ( .I(n3012), .Z(o_data_bus[1276]) );
  BUFFD6BWP30P140LVT U427 ( .I(n3013), .Z(o_data_bus[1275]) );
  BUFFD6BWP30P140LVT U428 ( .I(n3014), .Z(o_data_bus[1274]) );
  BUFFD6BWP30P140LVT U429 ( .I(n3015), .Z(o_data_bus[1273]) );
  BUFFD6BWP30P140LVT U430 ( .I(n3016), .Z(o_data_bus[1272]) );
  BUFFD6BWP30P140LVT U431 ( .I(n3017), .Z(o_data_bus[1271]) );
  BUFFD6BWP30P140LVT U432 ( .I(n3018), .Z(o_data_bus[1270]) );
  BUFFD6BWP30P140LVT U433 ( .I(n3019), .Z(o_data_bus[1269]) );
  BUFFD6BWP30P140LVT U434 ( .I(n3020), .Z(o_data_bus[1268]) );
  BUFFD6BWP30P140LVT U435 ( .I(n3021), .Z(o_data_bus[1267]) );
  BUFFD6BWP30P140LVT U436 ( .I(n3022), .Z(o_data_bus[1266]) );
  BUFFD6BWP30P140LVT U437 ( .I(n3023), .Z(o_data_bus[1265]) );
  BUFFD6BWP30P140LVT U438 ( .I(n3024), .Z(o_data_bus[1264]) );
  BUFFD6BWP30P140LVT U439 ( .I(n3025), .Z(o_data_bus[1263]) );
  BUFFD6BWP30P140LVT U440 ( .I(n3026), .Z(o_data_bus[1262]) );
  BUFFD6BWP30P140LVT U441 ( .I(n3027), .Z(o_data_bus[1261]) );
  BUFFD6BWP30P140LVT U442 ( .I(n3028), .Z(o_data_bus[1260]) );
  BUFFD6BWP30P140LVT U443 ( .I(n3029), .Z(o_data_bus[1259]) );
  BUFFD6BWP30P140LVT U444 ( .I(n3030), .Z(o_data_bus[1258]) );
  BUFFD6BWP30P140LVT U445 ( .I(n3031), .Z(o_data_bus[1257]) );
  BUFFD6BWP30P140LVT U446 ( .I(n3032), .Z(o_data_bus[1256]) );
  BUFFD6BWP30P140LVT U447 ( .I(n3033), .Z(o_data_bus[1255]) );
  BUFFD6BWP30P140LVT U448 ( .I(n3034), .Z(o_data_bus[1254]) );
  BUFFD6BWP30P140LVT U449 ( .I(n3035), .Z(o_data_bus[1253]) );
  BUFFD6BWP30P140LVT U450 ( .I(n3036), .Z(o_data_bus[1252]) );
  BUFFD6BWP30P140LVT U451 ( .I(n3037), .Z(o_data_bus[1251]) );
  BUFFD6BWP30P140LVT U452 ( .I(n3038), .Z(o_data_bus[1250]) );
  BUFFD6BWP30P140LVT U453 ( .I(n3039), .Z(o_data_bus[1249]) );
  BUFFD6BWP30P140LVT U454 ( .I(n3040), .Z(o_data_bus[1248]) );
  BUFFD6BWP30P140LVT U455 ( .I(n3041), .Z(o_data_bus[1247]) );
  BUFFD6BWP30P140LVT U456 ( .I(n3042), .Z(o_data_bus[1246]) );
  BUFFD6BWP30P140LVT U457 ( .I(n3043), .Z(o_data_bus[1245]) );
  BUFFD6BWP30P140LVT U458 ( .I(n3044), .Z(o_data_bus[1244]) );
  BUFFD6BWP30P140LVT U459 ( .I(n3045), .Z(o_data_bus[1243]) );
  BUFFD6BWP30P140LVT U460 ( .I(n3046), .Z(o_data_bus[1242]) );
  BUFFD6BWP30P140LVT U461 ( .I(n3047), .Z(o_data_bus[1241]) );
  BUFFD6BWP30P140LVT U462 ( .I(n3048), .Z(o_data_bus[1240]) );
  BUFFD6BWP30P140LVT U463 ( .I(n3049), .Z(o_data_bus[1239]) );
  BUFFD6BWP30P140LVT U464 ( .I(n3050), .Z(o_data_bus[1238]) );
  BUFFD6BWP30P140LVT U465 ( .I(n3051), .Z(o_data_bus[1237]) );
  BUFFD6BWP30P140LVT U466 ( .I(n3052), .Z(o_data_bus[1236]) );
  BUFFD6BWP30P140LVT U467 ( .I(n3053), .Z(o_data_bus[1235]) );
  BUFFD6BWP30P140LVT U468 ( .I(n3054), .Z(o_data_bus[1234]) );
  BUFFD6BWP30P140LVT U469 ( .I(n3055), .Z(o_data_bus[1233]) );
  BUFFD6BWP30P140LVT U470 ( .I(n3056), .Z(o_data_bus[1232]) );
  BUFFD6BWP30P140LVT U471 ( .I(n3057), .Z(o_data_bus[1231]) );
  BUFFD6BWP30P140LVT U472 ( .I(n3058), .Z(o_data_bus[1230]) );
  BUFFD6BWP30P140LVT U473 ( .I(n3059), .Z(o_data_bus[1229]) );
  BUFFD6BWP30P140LVT U474 ( .I(n3060), .Z(o_data_bus[1228]) );
  BUFFD6BWP30P140LVT U475 ( .I(n2993), .Z(o_data_bus[1295]) );
  BUFFD6BWP30P140LVT U476 ( .I(n3061), .Z(o_data_bus[1227]) );
  BUFFD6BWP30P140LVT U477 ( .I(n3062), .Z(o_data_bus[1226]) );
  BUFFD6BWP30P140LVT U478 ( .I(n3063), .Z(o_data_bus[1225]) );
  BUFFD6BWP30P140LVT U479 ( .I(n3064), .Z(o_data_bus[1224]) );
  BUFFD6BWP30P140LVT U480 ( .I(n3065), .Z(o_data_bus[1223]) );
  BUFFD6BWP30P140LVT U481 ( .I(n3066), .Z(o_data_bus[1222]) );
  BUFFD6BWP30P140LVT U482 ( .I(n3067), .Z(o_data_bus[1221]) );
  BUFFD6BWP30P140LVT U483 ( .I(n3068), .Z(o_data_bus[1220]) );
  BUFFD6BWP30P140LVT U484 ( .I(n3069), .Z(o_data_bus[1219]) );
  BUFFD6BWP30P140LVT U485 ( .I(n3070), .Z(o_data_bus[1218]) );
  BUFFD6BWP30P140LVT U486 ( .I(n3071), .Z(o_data_bus[1217]) );
  BUFFD6BWP30P140LVT U487 ( .I(n3072), .Z(o_data_bus[1216]) );
  BUFFD6BWP30P140LVT U488 ( .I(n3073), .Z(o_data_bus[1215]) );
  BUFFD6BWP30P140LVT U489 ( .I(n3074), .Z(o_data_bus[1214]) );
  BUFFD6BWP30P140LVT U490 ( .I(n3075), .Z(o_data_bus[1213]) );
  BUFFD6BWP30P140LVT U491 ( .I(n3076), .Z(o_data_bus[1212]) );
  BUFFD6BWP30P140LVT U492 ( .I(n3077), .Z(o_data_bus[1211]) );
  BUFFD6BWP30P140LVT U493 ( .I(n3078), .Z(o_data_bus[1210]) );
  BUFFD6BWP30P140LVT U494 ( .I(n3079), .Z(o_data_bus[1209]) );
  BUFFD6BWP30P140LVT U495 ( .I(n3080), .Z(o_data_bus[1208]) );
  BUFFD6BWP30P140LVT U496 ( .I(n3082), .Z(o_data_bus[1206]) );
  BUFFD6BWP30P140LVT U497 ( .I(n3083), .Z(o_data_bus[1205]) );
  BUFFD6BWP30P140LVT U498 ( .I(n3084), .Z(o_data_bus[1204]) );
  BUFFD6BWP30P140LVT U499 ( .I(n3085), .Z(o_data_bus[1203]) );
  BUFFD6BWP30P140LVT U500 ( .I(n3086), .Z(o_data_bus[1202]) );
  BUFFD6BWP30P140LVT U501 ( .I(n3087), .Z(o_data_bus[1201]) );
  BUFFD6BWP30P140LVT U502 ( .I(n3088), .Z(o_data_bus[1200]) );
  BUFFD6BWP30P140LVT U503 ( .I(n3089), .Z(o_data_bus[1199]) );
  BUFFD6BWP30P140LVT U504 ( .I(n3090), .Z(o_data_bus[1198]) );
  BUFFD6BWP30P140LVT U505 ( .I(n3091), .Z(o_data_bus[1197]) );
  BUFFD6BWP30P140LVT U506 ( .I(n3092), .Z(o_data_bus[1196]) );
  BUFFD6BWP30P140LVT U507 ( .I(n3093), .Z(o_data_bus[1195]) );
  BUFFD6BWP30P140LVT U508 ( .I(n3094), .Z(o_data_bus[1194]) );
  BUFFD6BWP30P140LVT U509 ( .I(n3095), .Z(o_data_bus[1193]) );
  BUFFD6BWP30P140LVT U510 ( .I(n3096), .Z(o_data_bus[1192]) );
  BUFFD6BWP30P140LVT U511 ( .I(n3097), .Z(o_data_bus[1191]) );
  BUFFD6BWP30P140LVT U512 ( .I(n3098), .Z(o_data_bus[1190]) );
  BUFFD6BWP30P140LVT U513 ( .I(n3099), .Z(o_data_bus[1189]) );
  BUFFD6BWP30P140LVT U514 ( .I(n3100), .Z(o_data_bus[1188]) );
  BUFFD6BWP30P140LVT U515 ( .I(n3101), .Z(o_data_bus[1187]) );
  BUFFD6BWP30P140LVT U516 ( .I(n3102), .Z(o_data_bus[1186]) );
  BUFFD6BWP30P140LVT U517 ( .I(n3103), .Z(o_data_bus[1185]) );
  BUFFD6BWP30P140LVT U518 ( .I(n3104), .Z(o_data_bus[1184]) );
  BUFFD6BWP30P140LVT U519 ( .I(n3105), .Z(o_data_bus[1183]) );
  BUFFD6BWP30P140LVT U520 ( .I(n3106), .Z(o_data_bus[1182]) );
  BUFFD6BWP30P140LVT U521 ( .I(n3107), .Z(o_data_bus[1181]) );
  BUFFD6BWP30P140LVT U522 ( .I(n3108), .Z(o_data_bus[1180]) );
  BUFFD6BWP30P140LVT U523 ( .I(n3109), .Z(o_data_bus[1179]) );
  BUFFD6BWP30P140LVT U524 ( .I(n3110), .Z(o_data_bus[1178]) );
  BUFFD6BWP30P140LVT U525 ( .I(n3111), .Z(o_data_bus[1177]) );
  BUFFD6BWP30P140LVT U526 ( .I(n3112), .Z(o_data_bus[1176]) );
  BUFFD6BWP30P140LVT U527 ( .I(n3113), .Z(o_data_bus[1175]) );
  BUFFD6BWP30P140LVT U528 ( .I(n3114), .Z(o_data_bus[1174]) );
  BUFFD6BWP30P140LVT U529 ( .I(n3115), .Z(o_data_bus[1173]) );
  BUFFD6BWP30P140LVT U530 ( .I(n3116), .Z(o_data_bus[1172]) );
  BUFFD6BWP30P140LVT U531 ( .I(n3117), .Z(o_data_bus[1171]) );
  BUFFD6BWP30P140LVT U532 ( .I(n3118), .Z(o_data_bus[1170]) );
  BUFFD6BWP30P140LVT U533 ( .I(n3119), .Z(o_data_bus[1169]) );
  BUFFD6BWP30P140LVT U534 ( .I(n3120), .Z(o_data_bus[1168]) );
  BUFFD6BWP30P140LVT U535 ( .I(n3121), .Z(o_data_bus[1167]) );
  BUFFD6BWP30P140LVT U536 ( .I(n3122), .Z(o_data_bus[1166]) );
  BUFFD6BWP30P140LVT U537 ( .I(n3123), .Z(o_data_bus[1165]) );
  BUFFD6BWP30P140LVT U538 ( .I(n3124), .Z(o_data_bus[1164]) );
  BUFFD6BWP30P140LVT U539 ( .I(n3125), .Z(o_data_bus[1163]) );
  BUFFD6BWP30P140LVT U540 ( .I(n3126), .Z(o_data_bus[1162]) );
  BUFFD6BWP30P140LVT U541 ( .I(n3127), .Z(o_data_bus[1161]) );
  BUFFD6BWP30P140LVT U542 ( .I(n3128), .Z(o_data_bus[1160]) );
  BUFFD6BWP30P140LVT U543 ( .I(n3264), .Z(o_data_bus[1024]) );
  BUFFD6BWP30P140LVT U544 ( .I(n2677), .Z(o_data_bus[1611]) );
  BUFFD6BWP30P140LVT U545 ( .I(n2678), .Z(o_data_bus[1610]) );
  BUFFD6BWP30P140LVT U546 ( .I(n2679), .Z(o_data_bus[1609]) );
  BUFFD6BWP30P140LVT U547 ( .I(n2680), .Z(o_data_bus[1608]) );
  BUFFD6BWP30P140LVT U548 ( .I(n2681), .Z(o_data_bus[1607]) );
  BUFFD6BWP30P140LVT U549 ( .I(n2682), .Z(o_data_bus[1606]) );
  BUFFD6BWP30P140LVT U550 ( .I(n2683), .Z(o_data_bus[1605]) );
  BUFFD6BWP30P140LVT U551 ( .I(n2684), .Z(o_data_bus[1604]) );
  BUFFD6BWP30P140LVT U552 ( .I(n2685), .Z(o_data_bus[1603]) );
  BUFFD6BWP30P140LVT U553 ( .I(n2686), .Z(o_data_bus[1602]) );
  BUFFD6BWP30P140LVT U554 ( .I(n2687), .Z(o_data_bus[1601]) );
  BUFFD6BWP30P140LVT U555 ( .I(n2688), .Z(o_data_bus[1600]) );
  BUFFD6BWP30P140LVT U556 ( .I(n2689), .Z(o_data_bus[1599]) );
  BUFFD6BWP30P140LVT U557 ( .I(n2690), .Z(o_data_bus[1598]) );
  BUFFD6BWP30P140LVT U558 ( .I(n2691), .Z(o_data_bus[1597]) );
  BUFFD6BWP30P140LVT U559 ( .I(n2692), .Z(o_data_bus[1596]) );
  BUFFD6BWP30P140LVT U560 ( .I(n2693), .Z(o_data_bus[1595]) );
  BUFFD6BWP30P140LVT U561 ( .I(n2694), .Z(o_data_bus[1594]) );
  BUFFD6BWP30P140LVT U562 ( .I(n2695), .Z(o_data_bus[1593]) );
  BUFFD6BWP30P140LVT U563 ( .I(n2696), .Z(o_data_bus[1592]) );
  BUFFD6BWP30P140LVT U564 ( .I(n2697), .Z(o_data_bus[1591]) );
  BUFFD6BWP30P140LVT U565 ( .I(n2698), .Z(o_data_bus[1590]) );
  BUFFD6BWP30P140LVT U566 ( .I(n2699), .Z(o_data_bus[1589]) );
  BUFFD6BWP30P140LVT U567 ( .I(n2700), .Z(o_data_bus[1588]) );
  BUFFD6BWP30P140LVT U568 ( .I(n2701), .Z(o_data_bus[1587]) );
  BUFFD6BWP30P140LVT U569 ( .I(n2702), .Z(o_data_bus[1586]) );
  BUFFD6BWP30P140LVT U570 ( .I(n2703), .Z(o_data_bus[1585]) );
  BUFFD6BWP30P140LVT U571 ( .I(n2704), .Z(o_data_bus[1584]) );
  BUFFD6BWP30P140LVT U572 ( .I(n2705), .Z(o_data_bus[1583]) );
  BUFFD6BWP30P140LVT U573 ( .I(n2706), .Z(o_data_bus[1582]) );
  BUFFD6BWP30P140LVT U574 ( .I(n2707), .Z(o_data_bus[1581]) );
  BUFFD6BWP30P140LVT U575 ( .I(n2708), .Z(o_data_bus[1580]) );
  BUFFD6BWP30P140LVT U576 ( .I(n2709), .Z(o_data_bus[1579]) );
  BUFFD6BWP30P140LVT U577 ( .I(n2710), .Z(o_data_bus[1578]) );
  BUFFD6BWP30P140LVT U578 ( .I(n2711), .Z(o_data_bus[1577]) );
  BUFFD6BWP30P140LVT U579 ( .I(n2712), .Z(o_data_bus[1576]) );
  BUFFD6BWP30P140LVT U580 ( .I(n2713), .Z(o_data_bus[1575]) );
  BUFFD6BWP30P140LVT U581 ( .I(n2714), .Z(o_data_bus[1574]) );
  BUFFD6BWP30P140LVT U582 ( .I(n2715), .Z(o_data_bus[1573]) );
  BUFFD6BWP30P140LVT U583 ( .I(n2716), .Z(o_data_bus[1572]) );
  BUFFD6BWP30P140LVT U584 ( .I(n2717), .Z(o_data_bus[1571]) );
  BUFFD6BWP30P140LVT U585 ( .I(n2718), .Z(o_data_bus[1570]) );
  BUFFD6BWP30P140LVT U586 ( .I(n2719), .Z(o_data_bus[1569]) );
  BUFFD6BWP30P140LVT U587 ( .I(n2720), .Z(o_data_bus[1568]) );
  BUFFD6BWP30P140LVT U588 ( .I(n3265), .Z(o_data_bus[1023]) );
  BUFFD6BWP30P140LVT U589 ( .I(n3946), .Z(o_data_bus[342]) );
  BUFFD6BWP30P140LVT U590 ( .I(n3947), .Z(o_data_bus[341]) );
  BUFFD6BWP30P140LVT U591 ( .I(n3948), .Z(o_data_bus[340]) );
  BUFFD6BWP30P140LVT U592 ( .I(n3949), .Z(o_data_bus[339]) );
  BUFFD6BWP30P140LVT U593 ( .I(n3950), .Z(o_data_bus[338]) );
  BUFFD6BWP30P140LVT U594 ( .I(n3951), .Z(o_data_bus[337]) );
  BUFFD6BWP30P140LVT U595 ( .I(n3952), .Z(o_data_bus[336]) );
  BUFFD6BWP30P140LVT U596 ( .I(n3953), .Z(o_data_bus[335]) );
  BUFFD6BWP30P140LVT U597 ( .I(n3954), .Z(o_data_bus[334]) );
  BUFFD6BWP30P140LVT U598 ( .I(n3955), .Z(o_data_bus[333]) );
  BUFFD6BWP30P140LVT U599 ( .I(n3956), .Z(o_data_bus[332]) );
  BUFFD6BWP30P140LVT U600 ( .I(n3957), .Z(o_data_bus[331]) );
  BUFFD6BWP30P140LVT U601 ( .I(n3958), .Z(o_data_bus[330]) );
  BUFFD6BWP30P140LVT U602 ( .I(n3959), .Z(o_data_bus[329]) );
  BUFFD6BWP30P140LVT U603 ( .I(n3960), .Z(o_data_bus[328]) );
  BUFFD6BWP30P140LVT U604 ( .I(n3961), .Z(o_data_bus[327]) );
  BUFFD6BWP30P140LVT U605 ( .I(n3962), .Z(o_data_bus[326]) );
  BUFFD6BWP30P140LVT U606 ( .I(n3963), .Z(o_data_bus[325]) );
  BUFFD6BWP30P140LVT U607 ( .I(n3964), .Z(o_data_bus[324]) );
  BUFFD6BWP30P140LVT U608 ( .I(n3965), .Z(o_data_bus[323]) );
  BUFFD6BWP30P140LVT U609 ( .I(n3966), .Z(o_data_bus[322]) );
  BUFFD6BWP30P140LVT U610 ( .I(n3967), .Z(o_data_bus[321]) );
  BUFFD6BWP30P140LVT U611 ( .I(n3968), .Z(o_data_bus[320]) );
  BUFFD6BWP30P140LVT U612 ( .I(n3969), .Z(o_data_bus[319]) );
  BUFFD6BWP30P140LVT U613 ( .I(n3970), .Z(o_data_bus[318]) );
  BUFFD6BWP30P140LVT U614 ( .I(n3971), .Z(o_data_bus[317]) );
  BUFFD6BWP30P140LVT U615 ( .I(n3972), .Z(o_data_bus[316]) );
  BUFFD6BWP30P140LVT U616 ( .I(n3973), .Z(o_data_bus[315]) );
  BUFFD6BWP30P140LVT U617 ( .I(n3974), .Z(o_data_bus[314]) );
  BUFFD6BWP30P140LVT U618 ( .I(n3975), .Z(o_data_bus[313]) );
  BUFFD6BWP30P140LVT U619 ( .I(n3976), .Z(o_data_bus[312]) );
  BUFFD6BWP30P140LVT U620 ( .I(n3977), .Z(o_data_bus[311]) );
  BUFFD6BWP30P140LVT U621 ( .I(n3978), .Z(o_data_bus[310]) );
  BUFFD6BWP30P140LVT U622 ( .I(n3979), .Z(o_data_bus[309]) );
  BUFFD6BWP30P140LVT U623 ( .I(n3980), .Z(o_data_bus[308]) );
  BUFFD6BWP30P140LVT U624 ( .I(n3981), .Z(o_data_bus[307]) );
  BUFFD6BWP30P140LVT U625 ( .I(n3982), .Z(o_data_bus[306]) );
  BUFFD6BWP30P140LVT U626 ( .I(n3983), .Z(o_data_bus[305]) );
  BUFFD6BWP30P140LVT U627 ( .I(n3984), .Z(o_data_bus[304]) );
  BUFFD6BWP30P140LVT U628 ( .I(n3985), .Z(o_data_bus[303]) );
  BUFFD6BWP30P140LVT U629 ( .I(n3986), .Z(o_data_bus[302]) );
  BUFFD6BWP30P140LVT U630 ( .I(n3987), .Z(o_data_bus[301]) );
  BUFFD6BWP30P140LVT U631 ( .I(n3988), .Z(o_data_bus[300]) );
  BUFFD6BWP30P140LVT U632 ( .I(n3989), .Z(o_data_bus[299]) );
  BUFFD6BWP30P140LVT U633 ( .I(n3990), .Z(o_data_bus[298]) );
  BUFFD6BWP30P140LVT U634 ( .I(n3991), .Z(o_data_bus[297]) );
  BUFFD6BWP30P140LVT U635 ( .I(n3992), .Z(o_data_bus[296]) );
  BUFFD6BWP30P140LVT U636 ( .I(n3993), .Z(o_data_bus[295]) );
  BUFFD6BWP30P140LVT U637 ( .I(n3994), .Z(o_data_bus[294]) );
  BUFFD6BWP30P140LVT U638 ( .I(n3995), .Z(o_data_bus[293]) );
  BUFFD6BWP30P140LVT U639 ( .I(n3996), .Z(o_data_bus[292]) );
  BUFFD6BWP30P140LVT U640 ( .I(n3997), .Z(o_data_bus[291]) );
  BUFFD6BWP30P140LVT U641 ( .I(n3998), .Z(o_data_bus[290]) );
  BUFFD6BWP30P140LVT U642 ( .I(n3999), .Z(o_data_bus[289]) );
  BUFFD6BWP30P140LVT U643 ( .I(n4000), .Z(o_data_bus[288]) );
  BUFFD6BWP30P140LVT U644 ( .I(n4001), .Z(o_data_bus[287]) );
  BUFFD6BWP30P140LVT U645 ( .I(n4002), .Z(o_data_bus[286]) );
  BUFFD6BWP30P140LVT U646 ( .I(n4003), .Z(o_data_bus[285]) );
  BUFFD6BWP30P140LVT U647 ( .I(n4004), .Z(o_data_bus[284]) );
  BUFFD6BWP30P140LVT U648 ( .I(n4005), .Z(o_data_bus[283]) );
  BUFFD6BWP30P140LVT U649 ( .I(n4006), .Z(o_data_bus[282]) );
  BUFFD6BWP30P140LVT U650 ( .I(n4007), .Z(o_data_bus[281]) );
  BUFFD6BWP30P140LVT U651 ( .I(n4008), .Z(o_data_bus[280]) );
  BUFFD6BWP30P140LVT U652 ( .I(n4009), .Z(o_data_bus[279]) );
  BUFFD6BWP30P140LVT U653 ( .I(n4010), .Z(o_data_bus[278]) );
  BUFFD6BWP30P140LVT U654 ( .I(n4011), .Z(o_data_bus[277]) );
  BUFFD6BWP30P140LVT U655 ( .I(n4012), .Z(o_data_bus[276]) );
  BUFFD6BWP30P140LVT U656 ( .I(n3945), .Z(o_data_bus[343]) );
  BUFFD6BWP30P140LVT U657 ( .I(n4013), .Z(o_data_bus[275]) );
  BUFFD6BWP30P140LVT U658 ( .I(n4014), .Z(o_data_bus[274]) );
  BUFFD6BWP30P140LVT U659 ( .I(n4015), .Z(o_data_bus[273]) );
  BUFFD6BWP30P140LVT U660 ( .I(n4016), .Z(o_data_bus[272]) );
  BUFFD6BWP30P140LVT U661 ( .I(n4017), .Z(o_data_bus[271]) );
  BUFFD6BWP30P140LVT U662 ( .I(n4018), .Z(o_data_bus[270]) );
  BUFFD6BWP30P140LVT U663 ( .I(n4019), .Z(o_data_bus[269]) );
  BUFFD6BWP30P140LVT U664 ( .I(n4020), .Z(o_data_bus[268]) );
  BUFFD6BWP30P140LVT U665 ( .I(n4021), .Z(o_data_bus[267]) );
  BUFFD6BWP30P140LVT U666 ( .I(n4022), .Z(o_data_bus[266]) );
  BUFFD6BWP30P140LVT U667 ( .I(n4023), .Z(o_data_bus[265]) );
  BUFFD6BWP30P140LVT U668 ( .I(n4024), .Z(o_data_bus[264]) );
  BUFFD6BWP30P140LVT U669 ( .I(n4025), .Z(o_data_bus[263]) );
  BUFFD6BWP30P140LVT U670 ( .I(n4026), .Z(o_data_bus[262]) );
  BUFFD6BWP30P140LVT U671 ( .I(n4027), .Z(o_data_bus[261]) );
  BUFFD6BWP30P140LVT U672 ( .I(n4028), .Z(o_data_bus[260]) );
  BUFFD6BWP30P140LVT U673 ( .I(n4029), .Z(o_data_bus[259]) );
  BUFFD6BWP30P140LVT U674 ( .I(n4030), .Z(o_data_bus[258]) );
  BUFFD6BWP30P140LVT U675 ( .I(n4031), .Z(o_data_bus[257]) );
  BUFFD6BWP30P140LVT U676 ( .I(n4032), .Z(o_data_bus[256]) );
  BUFFD6BWP30P140LVT U677 ( .I(n4033), .Z(o_data_bus[255]) );
  BUFFD6BWP30P140LVT U678 ( .I(n4034), .Z(o_data_bus[254]) );
  BUFFD6BWP30P140LVT U679 ( .I(n4035), .Z(o_data_bus[253]) );
  BUFFD6BWP30P140LVT U680 ( .I(n4036), .Z(o_data_bus[252]) );
  BUFFD6BWP30P140LVT U681 ( .I(n4037), .Z(o_data_bus[251]) );
  BUFFD6BWP30P140LVT U682 ( .I(n4038), .Z(o_data_bus[250]) );
  BUFFD6BWP30P140LVT U683 ( .I(n4039), .Z(o_data_bus[249]) );
  BUFFD6BWP30P140LVT U684 ( .I(n4040), .Z(o_data_bus[248]) );
  BUFFD6BWP30P140LVT U685 ( .I(n4041), .Z(o_data_bus[247]) );
  BUFFD6BWP30P140LVT U686 ( .I(n4042), .Z(o_data_bus[246]) );
  BUFFD6BWP30P140LVT U687 ( .I(n4043), .Z(o_data_bus[245]) );
  BUFFD6BWP30P140LVT U688 ( .I(n4044), .Z(o_data_bus[244]) );
  BUFFD6BWP30P140LVT U689 ( .I(n4045), .Z(o_data_bus[243]) );
  BUFFD6BWP30P140LVT U690 ( .I(n4046), .Z(o_data_bus[242]) );
  BUFFD6BWP30P140LVT U691 ( .I(n4047), .Z(o_data_bus[241]) );
  BUFFD6BWP30P140LVT U692 ( .I(n4048), .Z(o_data_bus[240]) );
  BUFFD6BWP30P140LVT U693 ( .I(n4049), .Z(o_data_bus[239]) );
  BUFFD6BWP30P140LVT U694 ( .I(n4050), .Z(o_data_bus[238]) );
  BUFFD6BWP30P140LVT U695 ( .I(n4051), .Z(o_data_bus[237]) );
  BUFFD6BWP30P140LVT U696 ( .I(n4052), .Z(o_data_bus[236]) );
  BUFFD6BWP30P140LVT U697 ( .I(n4053), .Z(o_data_bus[235]) );
  BUFFD6BWP30P140LVT U698 ( .I(n4054), .Z(o_data_bus[234]) );
  BUFFD6BWP30P140LVT U699 ( .I(n4055), .Z(o_data_bus[233]) );
  BUFFD6BWP30P140LVT U700 ( .I(n4056), .Z(o_data_bus[232]) );
  BUFFD6BWP30P140LVT U701 ( .I(n4057), .Z(o_data_bus[231]) );
  BUFFD6BWP30P140LVT U702 ( .I(n4058), .Z(o_data_bus[230]) );
  BUFFD6BWP30P140LVT U703 ( .I(n4059), .Z(o_data_bus[229]) );
  BUFFD6BWP30P140LVT U704 ( .I(n4060), .Z(o_data_bus[228]) );
  BUFFD6BWP30P140LVT U705 ( .I(n4061), .Z(o_data_bus[227]) );
  BUFFD6BWP30P140LVT U706 ( .I(n4062), .Z(o_data_bus[226]) );
  BUFFD6BWP30P140LVT U707 ( .I(n4063), .Z(o_data_bus[225]) );
  BUFFD6BWP30P140LVT U708 ( .I(n4064), .Z(o_data_bus[224]) );
  BUFFD6BWP30P140LVT U709 ( .I(n4065), .Z(o_data_bus[223]) );
  BUFFD6BWP30P140LVT U710 ( .I(n4066), .Z(o_data_bus[222]) );
  BUFFD6BWP30P140LVT U711 ( .I(n4067), .Z(o_data_bus[221]) );
  BUFFD6BWP30P140LVT U712 ( .I(n4068), .Z(o_data_bus[220]) );
  BUFFD6BWP30P140LVT U713 ( .I(n4069), .Z(o_data_bus[219]) );
  BUFFD6BWP30P140LVT U714 ( .I(n4070), .Z(o_data_bus[218]) );
  BUFFD6BWP30P140LVT U715 ( .I(n4071), .Z(o_data_bus[217]) );
  BUFFD6BWP30P140LVT U716 ( .I(n4072), .Z(o_data_bus[216]) );
  BUFFD6BWP30P140LVT U717 ( .I(n4073), .Z(o_data_bus[215]) );
  BUFFD6BWP30P140LVT U718 ( .I(n4074), .Z(o_data_bus[214]) );
  BUFFD6BWP30P140LVT U719 ( .I(n4075), .Z(o_data_bus[213]) );
  BUFFD6BWP30P140LVT U720 ( .I(n4076), .Z(o_data_bus[212]) );
  BUFFD6BWP30P140LVT U721 ( .I(n4077), .Z(o_data_bus[211]) );
  BUFFD6BWP30P140LVT U722 ( .I(n4078), .Z(o_data_bus[210]) );
  BUFFD6BWP30P140LVT U723 ( .I(n4079), .Z(o_data_bus[209]) );
  BUFFD6BWP30P140LVT U724 ( .I(n4080), .Z(o_data_bus[208]) );
  BUFFD6BWP30P140LVT U725 ( .I(n3811), .Z(o_data_bus[477]) );
  BUFFD6BWP30P140LVT U726 ( .I(n3812), .Z(o_data_bus[476]) );
  BUFFD6BWP30P140LVT U727 ( .I(n3813), .Z(o_data_bus[475]) );
  BUFFD6BWP30P140LVT U728 ( .I(n3814), .Z(o_data_bus[474]) );
  BUFFD6BWP30P140LVT U729 ( .I(n3815), .Z(o_data_bus[473]) );
  BUFFD6BWP30P140LVT U730 ( .I(n3816), .Z(o_data_bus[472]) );
  BUFFD6BWP30P140LVT U731 ( .I(n3817), .Z(o_data_bus[471]) );
  BUFFD6BWP30P140LVT U732 ( .I(n3818), .Z(o_data_bus[470]) );
  BUFFD6BWP30P140LVT U733 ( .I(n3819), .Z(o_data_bus[469]) );
  BUFFD6BWP30P140LVT U734 ( .I(n3820), .Z(o_data_bus[468]) );
  BUFFD6BWP30P140LVT U735 ( .I(n3821), .Z(o_data_bus[467]) );
  BUFFD6BWP30P140LVT U736 ( .I(n3822), .Z(o_data_bus[466]) );
  BUFFD6BWP30P140LVT U737 ( .I(n3823), .Z(o_data_bus[465]) );
  BUFFD6BWP30P140LVT U738 ( .I(n3824), .Z(o_data_bus[464]) );
  BUFFD6BWP30P140LVT U739 ( .I(n3825), .Z(o_data_bus[463]) );
  BUFFD6BWP30P140LVT U740 ( .I(n3826), .Z(o_data_bus[462]) );
  BUFFD6BWP30P140LVT U741 ( .I(n3827), .Z(o_data_bus[461]) );
  BUFFD6BWP30P140LVT U742 ( .I(n3828), .Z(o_data_bus[460]) );
  BUFFD6BWP30P140LVT U743 ( .I(n3829), .Z(o_data_bus[459]) );
  BUFFD6BWP30P140LVT U744 ( .I(n3830), .Z(o_data_bus[458]) );
  BUFFD6BWP30P140LVT U745 ( .I(n3831), .Z(o_data_bus[457]) );
  BUFFD6BWP30P140LVT U746 ( .I(n3832), .Z(o_data_bus[456]) );
  BUFFD6BWP30P140LVT U747 ( .I(n3833), .Z(o_data_bus[455]) );
  BUFFD6BWP30P140LVT U748 ( .I(n3834), .Z(o_data_bus[454]) );
  BUFFD6BWP30P140LVT U749 ( .I(n3835), .Z(o_data_bus[453]) );
  BUFFD6BWP30P140LVT U750 ( .I(n3836), .Z(o_data_bus[452]) );
  BUFFD6BWP30P140LVT U751 ( .I(n3837), .Z(o_data_bus[451]) );
  BUFFD6BWP30P140LVT U752 ( .I(n3838), .Z(o_data_bus[450]) );
  BUFFD6BWP30P140LVT U753 ( .I(n3839), .Z(o_data_bus[449]) );
  BUFFD6BWP30P140LVT U754 ( .I(n3840), .Z(o_data_bus[448]) );
  BUFFD6BWP30P140LVT U755 ( .I(n3841), .Z(o_data_bus[447]) );
  BUFFD6BWP30P140LVT U756 ( .I(n3842), .Z(o_data_bus[446]) );
  BUFFD6BWP30P140LVT U757 ( .I(n3843), .Z(o_data_bus[445]) );
  BUFFD6BWP30P140LVT U758 ( .I(n3844), .Z(o_data_bus[444]) );
  BUFFD6BWP30P140LVT U759 ( .I(n3845), .Z(o_data_bus[443]) );
  BUFFD6BWP30P140LVT U760 ( .I(n3846), .Z(o_data_bus[442]) );
  BUFFD6BWP30P140LVT U761 ( .I(n3847), .Z(o_data_bus[441]) );
  BUFFD6BWP30P140LVT U762 ( .I(n3848), .Z(o_data_bus[440]) );
  BUFFD6BWP30P140LVT U763 ( .I(n3849), .Z(o_data_bus[439]) );
  BUFFD6BWP30P140LVT U764 ( .I(n3850), .Z(o_data_bus[438]) );
  BUFFD6BWP30P140LVT U765 ( .I(n3851), .Z(o_data_bus[437]) );
  BUFFD6BWP30P140LVT U766 ( .I(n3852), .Z(o_data_bus[436]) );
  BUFFD6BWP30P140LVT U767 ( .I(n3853), .Z(o_data_bus[435]) );
  BUFFD6BWP30P140LVT U768 ( .I(n3854), .Z(o_data_bus[434]) );
  BUFFD6BWP30P140LVT U769 ( .I(n3855), .Z(o_data_bus[433]) );
  BUFFD6BWP30P140LVT U770 ( .I(n3856), .Z(o_data_bus[432]) );
  BUFFD6BWP30P140LVT U771 ( .I(n3857), .Z(o_data_bus[431]) );
  BUFFD6BWP30P140LVT U772 ( .I(n3858), .Z(o_data_bus[430]) );
  BUFFD6BWP30P140LVT U773 ( .I(n3859), .Z(o_data_bus[429]) );
  BUFFD6BWP30P140LVT U774 ( .I(n3860), .Z(o_data_bus[428]) );
  BUFFD6BWP30P140LVT U775 ( .I(n3861), .Z(o_data_bus[427]) );
  BUFFD6BWP30P140LVT U776 ( .I(n3862), .Z(o_data_bus[426]) );
  BUFFD6BWP30P140LVT U777 ( .I(n3863), .Z(o_data_bus[425]) );
  BUFFD6BWP30P140LVT U778 ( .I(n3864), .Z(o_data_bus[424]) );
  BUFFD6BWP30P140LVT U779 ( .I(n3865), .Z(o_data_bus[423]) );
  BUFFD6BWP30P140LVT U780 ( .I(n3866), .Z(o_data_bus[422]) );
  BUFFD6BWP30P140LVT U781 ( .I(n3867), .Z(o_data_bus[421]) );
  BUFFD6BWP30P140LVT U782 ( .I(n3868), .Z(o_data_bus[420]) );
  BUFFD6BWP30P140LVT U783 ( .I(n3869), .Z(o_data_bus[419]) );
  BUFFD6BWP30P140LVT U784 ( .I(n3870), .Z(o_data_bus[418]) );
  BUFFD6BWP30P140LVT U785 ( .I(n3871), .Z(o_data_bus[417]) );
  BUFFD6BWP30P140LVT U786 ( .I(n3872), .Z(o_data_bus[416]) );
  BUFFD6BWP30P140LVT U787 ( .I(n3873), .Z(o_data_bus[415]) );
  BUFFD6BWP30P140LVT U788 ( .I(n3874), .Z(o_data_bus[414]) );
  BUFFD6BWP30P140LVT U789 ( .I(n3875), .Z(o_data_bus[413]) );
  BUFFD6BWP30P140LVT U790 ( .I(n3876), .Z(o_data_bus[412]) );
  BUFFD6BWP30P140LVT U791 ( .I(n3877), .Z(o_data_bus[411]) );
  BUFFD6BWP30P140LVT U792 ( .I(n3810), .Z(o_data_bus[478]) );
  BUFFD6BWP30P140LVT U793 ( .I(n3878), .Z(o_data_bus[410]) );
  BUFFD6BWP30P140LVT U794 ( .I(n3879), .Z(o_data_bus[409]) );
  BUFFD6BWP30P140LVT U795 ( .I(n3880), .Z(o_data_bus[408]) );
  BUFFD6BWP30P140LVT U796 ( .I(n3881), .Z(o_data_bus[407]) );
  BUFFD6BWP30P140LVT U797 ( .I(n3882), .Z(o_data_bus[406]) );
  BUFFD6BWP30P140LVT U798 ( .I(n3883), .Z(o_data_bus[405]) );
  BUFFD6BWP30P140LVT U799 ( .I(n3884), .Z(o_data_bus[404]) );
  BUFFD6BWP30P140LVT U800 ( .I(n3885), .Z(o_data_bus[403]) );
  BUFFD6BWP30P140LVT U801 ( .I(n3886), .Z(o_data_bus[402]) );
  BUFFD6BWP30P140LVT U802 ( .I(n3887), .Z(o_data_bus[401]) );
  BUFFD6BWP30P140LVT U803 ( .I(n3888), .Z(o_data_bus[400]) );
  BUFFD6BWP30P140LVT U804 ( .I(n3889), .Z(o_data_bus[399]) );
  BUFFD6BWP30P140LVT U805 ( .I(n3890), .Z(o_data_bus[398]) );
  BUFFD6BWP30P140LVT U806 ( .I(n3891), .Z(o_data_bus[397]) );
  BUFFD6BWP30P140LVT U807 ( .I(n3892), .Z(o_data_bus[396]) );
  BUFFD6BWP30P140LVT U808 ( .I(n3893), .Z(o_data_bus[395]) );
  BUFFD6BWP30P140LVT U809 ( .I(n3894), .Z(o_data_bus[394]) );
  BUFFD6BWP30P140LVT U810 ( .I(n3895), .Z(o_data_bus[393]) );
  BUFFD6BWP30P140LVT U811 ( .I(n3896), .Z(o_data_bus[392]) );
  BUFFD6BWP30P140LVT U812 ( .I(n3897), .Z(o_data_bus[391]) );
  BUFFD6BWP30P140LVT U813 ( .I(n3898), .Z(o_data_bus[390]) );
  BUFFD6BWP30P140LVT U814 ( .I(n3899), .Z(o_data_bus[389]) );
  BUFFD6BWP30P140LVT U815 ( .I(n3900), .Z(o_data_bus[388]) );
  BUFFD6BWP30P140LVT U816 ( .I(n3901), .Z(o_data_bus[387]) );
  BUFFD6BWP30P140LVT U817 ( .I(n3902), .Z(o_data_bus[386]) );
  BUFFD6BWP30P140LVT U818 ( .I(n3903), .Z(o_data_bus[385]) );
  BUFFD6BWP30P140LVT U819 ( .I(n3904), .Z(o_data_bus[384]) );
  BUFFD6BWP30P140LVT U820 ( .I(n3905), .Z(o_data_bus[383]) );
  BUFFD6BWP30P140LVT U821 ( .I(n3906), .Z(o_data_bus[382]) );
  BUFFD6BWP30P140LVT U822 ( .I(n3907), .Z(o_data_bus[381]) );
  BUFFD6BWP30P140LVT U823 ( .I(n3908), .Z(o_data_bus[380]) );
  BUFFD6BWP30P140LVT U824 ( .I(n3909), .Z(o_data_bus[379]) );
  BUFFD6BWP30P140LVT U825 ( .I(n3910), .Z(o_data_bus[378]) );
  BUFFD6BWP30P140LVT U826 ( .I(n3911), .Z(o_data_bus[377]) );
  BUFFD6BWP30P140LVT U827 ( .I(n3912), .Z(o_data_bus[376]) );
  BUFFD6BWP30P140LVT U828 ( .I(n3913), .Z(o_data_bus[375]) );
  BUFFD6BWP30P140LVT U829 ( .I(n3914), .Z(o_data_bus[374]) );
  BUFFD6BWP30P140LVT U830 ( .I(n3915), .Z(o_data_bus[373]) );
  BUFFD6BWP30P140LVT U831 ( .I(n3916), .Z(o_data_bus[372]) );
  BUFFD6BWP30P140LVT U832 ( .I(n3917), .Z(o_data_bus[371]) );
  BUFFD6BWP30P140LVT U833 ( .I(n3918), .Z(o_data_bus[370]) );
  BUFFD6BWP30P140LVT U834 ( .I(n3919), .Z(o_data_bus[369]) );
  BUFFD6BWP30P140LVT U835 ( .I(n3920), .Z(o_data_bus[368]) );
  BUFFD6BWP30P140LVT U836 ( .I(n3921), .Z(o_data_bus[367]) );
  BUFFD6BWP30P140LVT U837 ( .I(n3922), .Z(o_data_bus[366]) );
  BUFFD6BWP30P140LVT U838 ( .I(n3923), .Z(o_data_bus[365]) );
  BUFFD6BWP30P140LVT U839 ( .I(n3924), .Z(o_data_bus[364]) );
  BUFFD6BWP30P140LVT U840 ( .I(n3925), .Z(o_data_bus[363]) );
  BUFFD6BWP30P140LVT U841 ( .I(n3926), .Z(o_data_bus[362]) );
  BUFFD6BWP30P140LVT U842 ( .I(n3927), .Z(o_data_bus[361]) );
  BUFFD6BWP30P140LVT U843 ( .I(n3928), .Z(o_data_bus[360]) );
  BUFFD6BWP30P140LVT U844 ( .I(n3929), .Z(o_data_bus[359]) );
  BUFFD6BWP30P140LVT U845 ( .I(n3930), .Z(o_data_bus[358]) );
  BUFFD6BWP30P140LVT U846 ( .I(n3931), .Z(o_data_bus[357]) );
  BUFFD6BWP30P140LVT U847 ( .I(n3932), .Z(o_data_bus[356]) );
  BUFFD6BWP30P140LVT U848 ( .I(n3933), .Z(o_data_bus[355]) );
  BUFFD6BWP30P140LVT U849 ( .I(n3934), .Z(o_data_bus[354]) );
  BUFFD6BWP30P140LVT U850 ( .I(n3935), .Z(o_data_bus[353]) );
  BUFFD6BWP30P140LVT U851 ( .I(n3936), .Z(o_data_bus[352]) );
  BUFFD6BWP30P140LVT U852 ( .I(n3937), .Z(o_data_bus[351]) );
  BUFFD6BWP30P140LVT U853 ( .I(n3938), .Z(o_data_bus[350]) );
  BUFFD6BWP30P140LVT U854 ( .I(n3939), .Z(o_data_bus[349]) );
  BUFFD6BWP30P140LVT U855 ( .I(n3940), .Z(o_data_bus[348]) );
  BUFFD6BWP30P140LVT U856 ( .I(n3941), .Z(o_data_bus[347]) );
  BUFFD6BWP30P140LVT U857 ( .I(n3942), .Z(o_data_bus[346]) );
  BUFFD6BWP30P140LVT U858 ( .I(n3943), .Z(o_data_bus[345]) );
  BUFFD6BWP30P140LVT U859 ( .I(n3944), .Z(o_data_bus[344]) );
  BUFFD6BWP30P140LVT U860 ( .I(n3809), .Z(o_data_bus[479]) );
  BUFFD6BWP30P140LVT U861 ( .I(n4217), .Z(o_data_bus[71]) );
  BUFFD6BWP30P140LVT U862 ( .I(n4218), .Z(o_data_bus[70]) );
  BUFFD6BWP30P140LVT U863 ( .I(n4219), .Z(o_data_bus[69]) );
  BUFFD6BWP30P140LVT U864 ( .I(n4220), .Z(o_data_bus[68]) );
  BUFFD6BWP30P140LVT U865 ( .I(n4221), .Z(o_data_bus[67]) );
  BUFFD6BWP30P140LVT U866 ( .I(n4222), .Z(o_data_bus[66]) );
  BUFFD6BWP30P140LVT U867 ( .I(n4223), .Z(o_data_bus[65]) );
  BUFFD6BWP30P140LVT U868 ( .I(n4224), .Z(o_data_bus[64]) );
  BUFFD6BWP30P140LVT U869 ( .I(n4225), .Z(o_data_bus[63]) );
  BUFFD6BWP30P140LVT U870 ( .I(n4226), .Z(o_data_bus[62]) );
  BUFFD6BWP30P140LVT U871 ( .I(n4227), .Z(o_data_bus[61]) );
  BUFFD6BWP30P140LVT U872 ( .I(n4228), .Z(o_data_bus[60]) );
  BUFFD6BWP30P140LVT U873 ( .I(n4229), .Z(o_data_bus[59]) );
  BUFFD6BWP30P140LVT U874 ( .I(n4230), .Z(o_data_bus[58]) );
  BUFFD6BWP30P140LVT U875 ( .I(n4231), .Z(o_data_bus[57]) );
  BUFFD6BWP30P140LVT U876 ( .I(n4232), .Z(o_data_bus[56]) );
  BUFFD6BWP30P140LVT U877 ( .I(n4233), .Z(o_data_bus[55]) );
  BUFFD6BWP30P140LVT U878 ( .I(n4234), .Z(o_data_bus[54]) );
  BUFFD6BWP30P140LVT U879 ( .I(n4235), .Z(o_data_bus[53]) );
  BUFFD6BWP30P140LVT U880 ( .I(n4236), .Z(o_data_bus[52]) );
  BUFFD6BWP30P140LVT U881 ( .I(n4237), .Z(o_data_bus[51]) );
  BUFFD6BWP30P140LVT U882 ( .I(n4238), .Z(o_data_bus[50]) );
  BUFFD6BWP30P140LVT U883 ( .I(n4239), .Z(o_data_bus[49]) );
  BUFFD6BWP30P140LVT U884 ( .I(n4240), .Z(o_data_bus[48]) );
  BUFFD6BWP30P140LVT U885 ( .I(n4241), .Z(o_data_bus[47]) );
  BUFFD6BWP30P140LVT U886 ( .I(n4242), .Z(o_data_bus[46]) );
  BUFFD6BWP30P140LVT U887 ( .I(n4243), .Z(o_data_bus[45]) );
  BUFFD6BWP30P140LVT U888 ( .I(n4244), .Z(o_data_bus[44]) );
  BUFFD6BWP30P140LVT U889 ( .I(n4245), .Z(o_data_bus[43]) );
  BUFFD6BWP30P140LVT U890 ( .I(n4246), .Z(o_data_bus[42]) );
  BUFFD6BWP30P140LVT U891 ( .I(n4247), .Z(o_data_bus[41]) );
  BUFFD6BWP30P140LVT U892 ( .I(n4248), .Z(o_data_bus[40]) );
  BUFFD6BWP30P140LVT U893 ( .I(n4249), .Z(o_data_bus[39]) );
  BUFFD6BWP30P140LVT U894 ( .I(n4250), .Z(o_data_bus[38]) );
  BUFFD6BWP30P140LVT U895 ( .I(n4251), .Z(o_data_bus[37]) );
  BUFFD6BWP30P140LVT U896 ( .I(n4252), .Z(o_data_bus[36]) );
  BUFFD6BWP30P140LVT U897 ( .I(n4253), .Z(o_data_bus[35]) );
  BUFFD6BWP30P140LVT U898 ( .I(n4254), .Z(o_data_bus[34]) );
  BUFFD6BWP30P140LVT U899 ( .I(n4255), .Z(o_data_bus[33]) );
  BUFFD6BWP30P140LVT U900 ( .I(n4256), .Z(o_data_bus[32]) );
  BUFFD6BWP30P140LVT U901 ( .I(n4257), .Z(o_data_bus[31]) );
  BUFFD6BWP30P140LVT U902 ( .I(n4258), .Z(o_data_bus[30]) );
  BUFFD6BWP30P140LVT U903 ( .I(n4259), .Z(o_data_bus[29]) );
  BUFFD6BWP30P140LVT U904 ( .I(n4260), .Z(o_data_bus[28]) );
  BUFFD6BWP30P140LVT U905 ( .I(n4261), .Z(o_data_bus[27]) );
  BUFFD6BWP30P140LVT U906 ( .I(n4262), .Z(o_data_bus[26]) );
  BUFFD6BWP30P140LVT U907 ( .I(n4263), .Z(o_data_bus[25]) );
  BUFFD6BWP30P140LVT U908 ( .I(n4264), .Z(o_data_bus[24]) );
  BUFFD6BWP30P140LVT U909 ( .I(n4265), .Z(o_data_bus[23]) );
  BUFFD6BWP30P140LVT U910 ( .I(n4266), .Z(o_data_bus[22]) );
  BUFFD6BWP30P140LVT U911 ( .I(n4267), .Z(o_data_bus[21]) );
  BUFFD6BWP30P140LVT U912 ( .I(n4268), .Z(o_data_bus[20]) );
  BUFFD6BWP30P140LVT U913 ( .I(n4269), .Z(o_data_bus[19]) );
  BUFFD6BWP30P140LVT U914 ( .I(n4270), .Z(o_data_bus[18]) );
  BUFFD6BWP30P140LVT U915 ( .I(n4271), .Z(o_data_bus[17]) );
  BUFFD6BWP30P140LVT U916 ( .I(n4272), .Z(o_data_bus[16]) );
  BUFFD6BWP30P140LVT U917 ( .I(n4273), .Z(o_data_bus[15]) );
  BUFFD6BWP30P140LVT U918 ( .I(n4274), .Z(o_data_bus[14]) );
  BUFFD6BWP30P140LVT U919 ( .I(n4275), .Z(o_data_bus[13]) );
  BUFFD6BWP30P140LVT U920 ( .I(n4276), .Z(o_data_bus[12]) );
  BUFFD6BWP30P140LVT U921 ( .I(n4277), .Z(o_data_bus[11]) );
  BUFFD6BWP30P140LVT U922 ( .I(n4278), .Z(o_data_bus[10]) );
  BUFFD6BWP30P140LVT U923 ( .I(n4279), .Z(o_data_bus[9]) );
  BUFFD6BWP30P140LVT U924 ( .I(n4280), .Z(o_data_bus[8]) );
  BUFFD6BWP30P140LVT U925 ( .I(n4281), .Z(o_data_bus[7]) );
  BUFFD6BWP30P140LVT U926 ( .I(n4282), .Z(o_data_bus[6]) );
  BUFFD6BWP30P140LVT U927 ( .I(n4283), .Z(o_data_bus[5]) );
  BUFFD6BWP30P140LVT U928 ( .I(n4216), .Z(o_data_bus[72]) );
  BUFFD6BWP30P140LVT U929 ( .I(n4284), .Z(o_data_bus[4]) );
  BUFFD6BWP30P140LVT U930 ( .I(n4285), .Z(o_data_bus[3]) );
  BUFFD6BWP30P140LVT U931 ( .I(n4286), .Z(o_data_bus[2]) );
  BUFFD6BWP30P140LVT U932 ( .I(n4287), .Z(o_data_bus[1]) );
  BUFFD6BWP30P140LVT U933 ( .I(n4288), .Z(o_data_bus[0]) );
  BUFFD6BWP30P140LVT U934 ( .I(n4289), .Z(o_cmd[63]) );
  BUFFD6BWP30P140LVT U935 ( .I(n4290), .Z(o_cmd[62]) );
  BUFFD6BWP30P140LVT U936 ( .I(n4291), .Z(o_cmd[61]) );
  BUFFD6BWP30P140LVT U937 ( .I(n4292), .Z(o_cmd[60]) );
  BUFFD6BWP30P140LVT U938 ( .I(n4293), .Z(o_cmd[59]) );
  BUFFD6BWP30P140LVT U939 ( .I(n4294), .Z(o_cmd[58]) );
  BUFFD6BWP30P140LVT U940 ( .I(n4295), .Z(o_cmd[57]) );
  BUFFD6BWP30P140LVT U941 ( .I(n4296), .Z(o_cmd[56]) );
  BUFFD6BWP30P140LVT U942 ( .I(n4297), .Z(o_cmd[55]) );
  BUFFD6BWP30P140LVT U943 ( .I(n4298), .Z(o_cmd[54]) );
  BUFFD6BWP30P140LVT U944 ( .I(n4299), .Z(o_cmd[53]) );
  BUFFD6BWP30P140LVT U945 ( .I(n4300), .Z(o_cmd[52]) );
  BUFFD6BWP30P140LVT U946 ( .I(n4301), .Z(o_cmd[51]) );
  BUFFD6BWP30P140LVT U947 ( .I(n4302), .Z(o_cmd[50]) );
  BUFFD6BWP30P140LVT U948 ( .I(n4303), .Z(o_cmd[49]) );
  BUFFD6BWP30P140LVT U949 ( .I(n4304), .Z(o_cmd[48]) );
  BUFFD6BWP30P140LVT U950 ( .I(n4305), .Z(o_cmd[47]) );
  BUFFD6BWP30P140LVT U951 ( .I(n4306), .Z(o_cmd[46]) );
  BUFFD6BWP30P140LVT U952 ( .I(n4307), .Z(o_cmd[45]) );
  BUFFD6BWP30P140LVT U953 ( .I(n4308), .Z(o_cmd[44]) );
  BUFFD6BWP30P140LVT U954 ( .I(n4309), .Z(o_cmd[43]) );
  BUFFD6BWP30P140LVT U955 ( .I(n4310), .Z(o_cmd[42]) );
  BUFFD6BWP30P140LVT U956 ( .I(n4311), .Z(o_cmd[41]) );
  BUFFD6BWP30P140LVT U957 ( .I(n4312), .Z(o_cmd[40]) );
  BUFFD6BWP30P140LVT U958 ( .I(n4313), .Z(o_cmd[39]) );
  BUFFD6BWP30P140LVT U959 ( .I(n4314), .Z(o_cmd[38]) );
  BUFFD6BWP30P140LVT U960 ( .I(n4315), .Z(o_cmd[37]) );
  BUFFD6BWP30P140LVT U961 ( .I(n4316), .Z(o_cmd[36]) );
  BUFFD6BWP30P140LVT U962 ( .I(n4317), .Z(o_cmd[35]) );
  BUFFD6BWP30P140LVT U963 ( .I(n4318), .Z(o_cmd[34]) );
  BUFFD6BWP30P140LVT U964 ( .I(n4319), .Z(o_cmd[33]) );
  BUFFD6BWP30P140LVT U965 ( .I(n4320), .Z(o_cmd[32]) );
  BUFFD6BWP30P140LVT U966 ( .I(n4321), .Z(o_cmd[31]) );
  BUFFD6BWP30P140LVT U967 ( .I(n4322), .Z(o_cmd[30]) );
  BUFFD6BWP30P140LVT U968 ( .I(n4323), .Z(o_cmd[29]) );
  BUFFD6BWP30P140LVT U969 ( .I(n4324), .Z(o_cmd[28]) );
  BUFFD6BWP30P140LVT U970 ( .I(n4325), .Z(o_cmd[27]) );
  BUFFD6BWP30P140LVT U971 ( .I(n4326), .Z(o_cmd[26]) );
  BUFFD6BWP30P140LVT U972 ( .I(n4327), .Z(o_cmd[25]) );
  BUFFD6BWP30P140LVT U973 ( .I(n4328), .Z(o_cmd[24]) );
  BUFFD6BWP30P140LVT U974 ( .I(n4329), .Z(o_cmd[23]) );
  BUFFD6BWP30P140LVT U975 ( .I(n4330), .Z(o_cmd[22]) );
  BUFFD6BWP30P140LVT U976 ( .I(n4331), .Z(o_cmd[21]) );
  BUFFD6BWP30P140LVT U977 ( .I(n4332), .Z(o_cmd[20]) );
  BUFFD6BWP30P140LVT U978 ( .I(n4333), .Z(o_cmd[19]) );
  BUFFD6BWP30P140LVT U979 ( .I(n4334), .Z(o_cmd[18]) );
  BUFFD6BWP30P140LVT U980 ( .I(n4335), .Z(o_cmd[17]) );
  BUFFD6BWP30P140LVT U981 ( .I(n4336), .Z(o_cmd[16]) );
  BUFFD6BWP30P140LVT U982 ( .I(n4337), .Z(o_cmd[15]) );
  BUFFD6BWP30P140LVT U983 ( .I(n4338), .Z(o_cmd[14]) );
  BUFFD6BWP30P140LVT U984 ( .I(n4339), .Z(o_cmd[13]) );
  BUFFD6BWP30P140LVT U985 ( .I(n4340), .Z(o_cmd[12]) );
  BUFFD6BWP30P140LVT U986 ( .I(n4341), .Z(o_cmd[11]) );
  BUFFD6BWP30P140LVT U987 ( .I(n4342), .Z(o_cmd[10]) );
  BUFFD6BWP30P140LVT U988 ( .I(n4343), .Z(o_cmd[9]) );
  BUFFD6BWP30P140LVT U989 ( .I(n4344), .Z(o_cmd[8]) );
  BUFFD6BWP30P140LVT U990 ( .I(n4345), .Z(o_cmd[7]) );
  BUFFD6BWP30P140LVT U991 ( .I(n4346), .Z(o_cmd[6]) );
  BUFFD6BWP30P140LVT U992 ( .I(n4347), .Z(o_cmd[5]) );
  BUFFD6BWP30P140LVT U993 ( .I(n4348), .Z(o_cmd[4]) );
  BUFFD6BWP30P140LVT U994 ( .I(n4349), .Z(o_cmd[3]) );
  BUFFD6BWP30P140LVT U995 ( .I(n4350), .Z(o_cmd[2]) );
  BUFFD6BWP30P140LVT U996 ( .I(n4351), .Z(o_cmd[1]) );
  BUFFD6BWP30P140LVT U997 ( .I(n4082), .Z(o_data_bus[206]) );
  BUFFD6BWP30P140LVT U998 ( .I(n4083), .Z(o_data_bus[205]) );
  BUFFD6BWP30P140LVT U999 ( .I(n4084), .Z(o_data_bus[204]) );
  BUFFD6BWP30P140LVT U1000 ( .I(n4085), .Z(o_data_bus[203]) );
  BUFFD6BWP30P140LVT U1001 ( .I(n4086), .Z(o_data_bus[202]) );
  BUFFD6BWP30P140LVT U1002 ( .I(n4087), .Z(o_data_bus[201]) );
  BUFFD6BWP30P140LVT U1003 ( .I(n4088), .Z(o_data_bus[200]) );
  BUFFD6BWP30P140LVT U1004 ( .I(n4089), .Z(o_data_bus[199]) );
  BUFFD6BWP30P140LVT U1005 ( .I(n4090), .Z(o_data_bus[198]) );
  BUFFD6BWP30P140LVT U1006 ( .I(n4091), .Z(o_data_bus[197]) );
  BUFFD6BWP30P140LVT U1007 ( .I(n4092), .Z(o_data_bus[196]) );
  BUFFD6BWP30P140LVT U1008 ( .I(n4093), .Z(o_data_bus[195]) );
  BUFFD6BWP30P140LVT U1009 ( .I(n4094), .Z(o_data_bus[194]) );
  BUFFD6BWP30P140LVT U1010 ( .I(n4095), .Z(o_data_bus[193]) );
  BUFFD6BWP30P140LVT U1011 ( .I(n4096), .Z(o_data_bus[192]) );
  BUFFD6BWP30P140LVT U1012 ( .I(n4097), .Z(o_data_bus[191]) );
  BUFFD6BWP30P140LVT U1013 ( .I(n4098), .Z(o_data_bus[190]) );
  BUFFD6BWP30P140LVT U1014 ( .I(n4099), .Z(o_data_bus[189]) );
  BUFFD6BWP30P140LVT U1015 ( .I(n4100), .Z(o_data_bus[188]) );
  BUFFD6BWP30P140LVT U1016 ( .I(n4101), .Z(o_data_bus[187]) );
  BUFFD6BWP30P140LVT U1017 ( .I(n4102), .Z(o_data_bus[186]) );
  BUFFD6BWP30P140LVT U1018 ( .I(n4103), .Z(o_data_bus[185]) );
  BUFFD6BWP30P140LVT U1019 ( .I(n4104), .Z(o_data_bus[184]) );
  BUFFD6BWP30P140LVT U1020 ( .I(n4105), .Z(o_data_bus[183]) );
  BUFFD6BWP30P140LVT U1021 ( .I(n4106), .Z(o_data_bus[182]) );
  BUFFD6BWP30P140LVT U1022 ( .I(n4107), .Z(o_data_bus[181]) );
  BUFFD6BWP30P140LVT U1023 ( .I(n4108), .Z(o_data_bus[180]) );
  BUFFD6BWP30P140LVT U1024 ( .I(n4109), .Z(o_data_bus[179]) );
  BUFFD6BWP30P140LVT U1025 ( .I(n4110), .Z(o_data_bus[178]) );
  BUFFD6BWP30P140LVT U1026 ( .I(n4111), .Z(o_data_bus[177]) );
  BUFFD6BWP30P140LVT U1027 ( .I(n4112), .Z(o_data_bus[176]) );
  BUFFD6BWP30P140LVT U1028 ( .I(n4113), .Z(o_data_bus[175]) );
  BUFFD6BWP30P140LVT U1029 ( .I(n4114), .Z(o_data_bus[174]) );
  BUFFD6BWP30P140LVT U1030 ( .I(n4115), .Z(o_data_bus[173]) );
  BUFFD6BWP30P140LVT U1031 ( .I(n4116), .Z(o_data_bus[172]) );
  BUFFD6BWP30P140LVT U1032 ( .I(n4117), .Z(o_data_bus[171]) );
  BUFFD6BWP30P140LVT U1033 ( .I(n4118), .Z(o_data_bus[170]) );
  BUFFD6BWP30P140LVT U1034 ( .I(n4119), .Z(o_data_bus[169]) );
  BUFFD6BWP30P140LVT U1035 ( .I(n4120), .Z(o_data_bus[168]) );
  BUFFD6BWP30P140LVT U1036 ( .I(n4121), .Z(o_data_bus[167]) );
  BUFFD6BWP30P140LVT U1037 ( .I(n4122), .Z(o_data_bus[166]) );
  BUFFD6BWP30P140LVT U1038 ( .I(n4123), .Z(o_data_bus[165]) );
  BUFFD6BWP30P140LVT U1039 ( .I(n4124), .Z(o_data_bus[164]) );
  BUFFD6BWP30P140LVT U1040 ( .I(n4125), .Z(o_data_bus[163]) );
  BUFFD6BWP30P140LVT U1041 ( .I(n4126), .Z(o_data_bus[162]) );
  BUFFD6BWP30P140LVT U1042 ( .I(n4127), .Z(o_data_bus[161]) );
  BUFFD6BWP30P140LVT U1043 ( .I(n4128), .Z(o_data_bus[160]) );
  BUFFD6BWP30P140LVT U1044 ( .I(n4129), .Z(o_data_bus[159]) );
  BUFFD6BWP30P140LVT U1045 ( .I(n4130), .Z(o_data_bus[158]) );
  BUFFD6BWP30P140LVT U1046 ( .I(n4131), .Z(o_data_bus[157]) );
  BUFFD6BWP30P140LVT U1047 ( .I(n4132), .Z(o_data_bus[156]) );
  BUFFD6BWP30P140LVT U1048 ( .I(n4133), .Z(o_data_bus[155]) );
  BUFFD6BWP30P140LVT U1049 ( .I(n4134), .Z(o_data_bus[154]) );
  BUFFD6BWP30P140LVT U1050 ( .I(n4135), .Z(o_data_bus[153]) );
  BUFFD6BWP30P140LVT U1051 ( .I(n4136), .Z(o_data_bus[152]) );
  BUFFD6BWP30P140LVT U1052 ( .I(n4137), .Z(o_data_bus[151]) );
  BUFFD6BWP30P140LVT U1053 ( .I(n4138), .Z(o_data_bus[150]) );
  BUFFD6BWP30P140LVT U1054 ( .I(n4139), .Z(o_data_bus[149]) );
  BUFFD6BWP30P140LVT U1055 ( .I(n4140), .Z(o_data_bus[148]) );
  BUFFD6BWP30P140LVT U1056 ( .I(n4141), .Z(o_data_bus[147]) );
  BUFFD6BWP30P140LVT U1057 ( .I(n4142), .Z(o_data_bus[146]) );
  BUFFD6BWP30P140LVT U1058 ( .I(n4143), .Z(o_data_bus[145]) );
  BUFFD6BWP30P140LVT U1059 ( .I(n4144), .Z(o_data_bus[144]) );
  BUFFD6BWP30P140LVT U1060 ( .I(n4145), .Z(o_data_bus[143]) );
  BUFFD6BWP30P140LVT U1061 ( .I(n4146), .Z(o_data_bus[142]) );
  BUFFD6BWP30P140LVT U1062 ( .I(n4147), .Z(o_data_bus[141]) );
  BUFFD6BWP30P140LVT U1063 ( .I(n4148), .Z(o_data_bus[140]) );
  BUFFD6BWP30P140LVT U1064 ( .I(n4081), .Z(o_data_bus[207]) );
  BUFFD6BWP30P140LVT U1065 ( .I(n4149), .Z(o_data_bus[139]) );
  BUFFD6BWP30P140LVT U1066 ( .I(n4150), .Z(o_data_bus[138]) );
  BUFFD6BWP30P140LVT U1067 ( .I(n4151), .Z(o_data_bus[137]) );
  BUFFD6BWP30P140LVT U1068 ( .I(n4152), .Z(o_data_bus[136]) );
  BUFFD6BWP30P140LVT U1069 ( .I(n4153), .Z(o_data_bus[135]) );
  BUFFD6BWP30P140LVT U1070 ( .I(n4154), .Z(o_data_bus[134]) );
  BUFFD6BWP30P140LVT U1071 ( .I(n4155), .Z(o_data_bus[133]) );
  BUFFD6BWP30P140LVT U1072 ( .I(n4156), .Z(o_data_bus[132]) );
  BUFFD6BWP30P140LVT U1073 ( .I(n4157), .Z(o_data_bus[131]) );
  BUFFD6BWP30P140LVT U1074 ( .I(n4158), .Z(o_data_bus[130]) );
  BUFFD6BWP30P140LVT U1075 ( .I(n4159), .Z(o_data_bus[129]) );
  BUFFD6BWP30P140LVT U1076 ( .I(n4160), .Z(o_data_bus[128]) );
  BUFFD6BWP30P140LVT U1077 ( .I(n4161), .Z(o_data_bus[127]) );
  BUFFD6BWP30P140LVT U1078 ( .I(n4162), .Z(o_data_bus[126]) );
  BUFFD6BWP30P140LVT U1079 ( .I(n4163), .Z(o_data_bus[125]) );
  BUFFD6BWP30P140LVT U1080 ( .I(n4164), .Z(o_data_bus[124]) );
  BUFFD6BWP30P140LVT U1081 ( .I(n4165), .Z(o_data_bus[123]) );
  BUFFD6BWP30P140LVT U1082 ( .I(n4166), .Z(o_data_bus[122]) );
  BUFFD6BWP30P140LVT U1083 ( .I(n4167), .Z(o_data_bus[121]) );
  BUFFD6BWP30P140LVT U1084 ( .I(n4168), .Z(o_data_bus[120]) );
  BUFFD6BWP30P140LVT U1085 ( .I(n4169), .Z(o_data_bus[119]) );
  BUFFD6BWP30P140LVT U1086 ( .I(n4170), .Z(o_data_bus[118]) );
  BUFFD6BWP30P140LVT U1087 ( .I(n4171), .Z(o_data_bus[117]) );
  BUFFD6BWP30P140LVT U1088 ( .I(n4172), .Z(o_data_bus[116]) );
  BUFFD6BWP30P140LVT U1089 ( .I(n4173), .Z(o_data_bus[115]) );
  BUFFD6BWP30P140LVT U1090 ( .I(n4174), .Z(o_data_bus[114]) );
  BUFFD6BWP30P140LVT U1091 ( .I(n4175), .Z(o_data_bus[113]) );
  BUFFD6BWP30P140LVT U1092 ( .I(n4176), .Z(o_data_bus[112]) );
  BUFFD6BWP30P140LVT U1093 ( .I(n4177), .Z(o_data_bus[111]) );
  BUFFD6BWP30P140LVT U1094 ( .I(n4178), .Z(o_data_bus[110]) );
  BUFFD6BWP30P140LVT U1095 ( .I(n4179), .Z(o_data_bus[109]) );
  BUFFD6BWP30P140LVT U1096 ( .I(n4180), .Z(o_data_bus[108]) );
  BUFFD6BWP30P140LVT U1097 ( .I(n4181), .Z(o_data_bus[107]) );
  BUFFD6BWP30P140LVT U1098 ( .I(n4182), .Z(o_data_bus[106]) );
  BUFFD6BWP30P140LVT U1099 ( .I(n4183), .Z(o_data_bus[105]) );
  BUFFD6BWP30P140LVT U1100 ( .I(n4184), .Z(o_data_bus[104]) );
  BUFFD6BWP30P140LVT U1101 ( .I(n4185), .Z(o_data_bus[103]) );
  BUFFD6BWP30P140LVT U1102 ( .I(n4186), .Z(o_data_bus[102]) );
  BUFFD6BWP30P140LVT U1103 ( .I(n4187), .Z(o_data_bus[101]) );
  BUFFD6BWP30P140LVT U1104 ( .I(n4188), .Z(o_data_bus[100]) );
  BUFFD6BWP30P140LVT U1105 ( .I(n4189), .Z(o_data_bus[99]) );
  BUFFD6BWP30P140LVT U1106 ( .I(n4190), .Z(o_data_bus[98]) );
  BUFFD6BWP30P140LVT U1107 ( .I(n4191), .Z(o_data_bus[97]) );
  BUFFD6BWP30P140LVT U1108 ( .I(n4192), .Z(o_data_bus[96]) );
  BUFFD6BWP30P140LVT U1109 ( .I(n4193), .Z(o_data_bus[95]) );
  BUFFD6BWP30P140LVT U1110 ( .I(n4194), .Z(o_data_bus[94]) );
  BUFFD6BWP30P140LVT U1111 ( .I(n4195), .Z(o_data_bus[93]) );
  BUFFD6BWP30P140LVT U1112 ( .I(n4196), .Z(o_data_bus[92]) );
  BUFFD6BWP30P140LVT U1113 ( .I(n4197), .Z(o_data_bus[91]) );
  BUFFD6BWP30P140LVT U1114 ( .I(n4198), .Z(o_data_bus[90]) );
  BUFFD6BWP30P140LVT U1115 ( .I(n4199), .Z(o_data_bus[89]) );
  BUFFD6BWP30P140LVT U1116 ( .I(n4200), .Z(o_data_bus[88]) );
  BUFFD6BWP30P140LVT U1117 ( .I(n4201), .Z(o_data_bus[87]) );
  BUFFD6BWP30P140LVT U1118 ( .I(n4202), .Z(o_data_bus[86]) );
  BUFFD6BWP30P140LVT U1119 ( .I(n4203), .Z(o_data_bus[85]) );
  BUFFD6BWP30P140LVT U1120 ( .I(n4204), .Z(o_data_bus[84]) );
  BUFFD6BWP30P140LVT U1121 ( .I(n4205), .Z(o_data_bus[83]) );
  BUFFD6BWP30P140LVT U1122 ( .I(n4206), .Z(o_data_bus[82]) );
  BUFFD6BWP30P140LVT U1123 ( .I(n4207), .Z(o_data_bus[81]) );
  BUFFD6BWP30P140LVT U1124 ( .I(n4208), .Z(o_data_bus[80]) );
  BUFFD6BWP30P140LVT U1125 ( .I(n4209), .Z(o_data_bus[79]) );
  BUFFD6BWP30P140LVT U1126 ( .I(n4210), .Z(o_data_bus[78]) );
  BUFFD6BWP30P140LVT U1127 ( .I(n4211), .Z(o_data_bus[77]) );
  BUFFD6BWP30P140LVT U1128 ( .I(n4212), .Z(o_data_bus[76]) );
  BUFFD6BWP30P140LVT U1129 ( .I(n4213), .Z(o_data_bus[75]) );
  BUFFD6BWP30P140LVT U1130 ( .I(n4214), .Z(o_data_bus[74]) );
  BUFFD6BWP30P140LVT U1131 ( .I(n4215), .Z(o_data_bus[73]) );
  BUFFD6BWP30P140LVT U1132 ( .I(n3808), .Z(o_data_bus[480]) );
  BUFFD6BWP30P140LVT U1133 ( .I(n3402), .Z(o_data_bus[886]) );
  BUFFD6BWP30P140LVT U1134 ( .I(n3403), .Z(o_data_bus[885]) );
  BUFFD6BWP30P140LVT U1135 ( .I(n3404), .Z(o_data_bus[884]) );
  BUFFD6BWP30P140LVT U1136 ( .I(n3405), .Z(o_data_bus[883]) );
  BUFFD6BWP30P140LVT U1137 ( .I(n3406), .Z(o_data_bus[882]) );
  BUFFD6BWP30P140LVT U1138 ( .I(n3407), .Z(o_data_bus[881]) );
  BUFFD6BWP30P140LVT U1139 ( .I(n3408), .Z(o_data_bus[880]) );
  BUFFD6BWP30P140LVT U1140 ( .I(n3409), .Z(o_data_bus[879]) );
  BUFFD6BWP30P140LVT U1141 ( .I(n3410), .Z(o_data_bus[878]) );
  BUFFD6BWP30P140LVT U1142 ( .I(n3411), .Z(o_data_bus[877]) );
  BUFFD6BWP30P140LVT U1143 ( .I(n3412), .Z(o_data_bus[876]) );
  BUFFD6BWP30P140LVT U1144 ( .I(n3413), .Z(o_data_bus[875]) );
  BUFFD6BWP30P140LVT U1145 ( .I(n3414), .Z(o_data_bus[874]) );
  BUFFD6BWP30P140LVT U1146 ( .I(n3415), .Z(o_data_bus[873]) );
  BUFFD6BWP30P140LVT U1147 ( .I(n3416), .Z(o_data_bus[872]) );
  BUFFD6BWP30P140LVT U1148 ( .I(n3417), .Z(o_data_bus[871]) );
  BUFFD6BWP30P140LVT U1149 ( .I(n3418), .Z(o_data_bus[870]) );
  BUFFD6BWP30P140LVT U1150 ( .I(n3419), .Z(o_data_bus[869]) );
  BUFFD6BWP30P140LVT U1151 ( .I(n3420), .Z(o_data_bus[868]) );
  BUFFD6BWP30P140LVT U1152 ( .I(n3421), .Z(o_data_bus[867]) );
  BUFFD6BWP30P140LVT U1153 ( .I(n3422), .Z(o_data_bus[866]) );
  BUFFD6BWP30P140LVT U1154 ( .I(n3423), .Z(o_data_bus[865]) );
  BUFFD6BWP30P140LVT U1155 ( .I(n3424), .Z(o_data_bus[864]) );
  BUFFD6BWP30P140LVT U1156 ( .I(n3425), .Z(o_data_bus[863]) );
  BUFFD6BWP30P140LVT U1157 ( .I(n3426), .Z(o_data_bus[862]) );
  BUFFD6BWP30P140LVT U1158 ( .I(n3427), .Z(o_data_bus[861]) );
  BUFFD6BWP30P140LVT U1159 ( .I(n3428), .Z(o_data_bus[860]) );
  BUFFD6BWP30P140LVT U1160 ( .I(n3429), .Z(o_data_bus[859]) );
  BUFFD6BWP30P140LVT U1161 ( .I(n3430), .Z(o_data_bus[858]) );
  BUFFD6BWP30P140LVT U1162 ( .I(n3431), .Z(o_data_bus[857]) );
  BUFFD6BWP30P140LVT U1163 ( .I(n3432), .Z(o_data_bus[856]) );
  BUFFD6BWP30P140LVT U1164 ( .I(n3433), .Z(o_data_bus[855]) );
  BUFFD6BWP30P140LVT U1165 ( .I(n3434), .Z(o_data_bus[854]) );
  BUFFD6BWP30P140LVT U1166 ( .I(n3435), .Z(o_data_bus[853]) );
  BUFFD6BWP30P140LVT U1167 ( .I(n3436), .Z(o_data_bus[852]) );
  BUFFD6BWP30P140LVT U1168 ( .I(n3437), .Z(o_data_bus[851]) );
  BUFFD6BWP30P140LVT U1169 ( .I(n3438), .Z(o_data_bus[850]) );
  BUFFD6BWP30P140LVT U1170 ( .I(n3439), .Z(o_data_bus[849]) );
  BUFFD6BWP30P140LVT U1171 ( .I(n3440), .Z(o_data_bus[848]) );
  BUFFD6BWP30P140LVT U1172 ( .I(n3441), .Z(o_data_bus[847]) );
  BUFFD6BWP30P140LVT U1173 ( .I(n3442), .Z(o_data_bus[846]) );
  BUFFD6BWP30P140LVT U1174 ( .I(n3443), .Z(o_data_bus[845]) );
  BUFFD6BWP30P140LVT U1175 ( .I(n3444), .Z(o_data_bus[844]) );
  BUFFD6BWP30P140LVT U1176 ( .I(n3445), .Z(o_data_bus[843]) );
  BUFFD6BWP30P140LVT U1177 ( .I(n3446), .Z(o_data_bus[842]) );
  BUFFD6BWP30P140LVT U1178 ( .I(n3447), .Z(o_data_bus[841]) );
  BUFFD6BWP30P140LVT U1179 ( .I(n3448), .Z(o_data_bus[840]) );
  BUFFD6BWP30P140LVT U1180 ( .I(n3449), .Z(o_data_bus[839]) );
  BUFFD6BWP30P140LVT U1181 ( .I(n3450), .Z(o_data_bus[838]) );
  BUFFD6BWP30P140LVT U1182 ( .I(n3451), .Z(o_data_bus[837]) );
  BUFFD6BWP30P140LVT U1183 ( .I(n3452), .Z(o_data_bus[836]) );
  BUFFD6BWP30P140LVT U1184 ( .I(n3453), .Z(o_data_bus[835]) );
  BUFFD6BWP30P140LVT U1185 ( .I(n3454), .Z(o_data_bus[834]) );
  BUFFD6BWP30P140LVT U1186 ( .I(n3455), .Z(o_data_bus[833]) );
  BUFFD6BWP30P140LVT U1187 ( .I(n3456), .Z(o_data_bus[832]) );
  BUFFD6BWP30P140LVT U1188 ( .I(n3457), .Z(o_data_bus[831]) );
  BUFFD6BWP30P140LVT U1189 ( .I(n3458), .Z(o_data_bus[830]) );
  BUFFD6BWP30P140LVT U1190 ( .I(n3459), .Z(o_data_bus[829]) );
  BUFFD6BWP30P140LVT U1191 ( .I(n3460), .Z(o_data_bus[828]) );
  BUFFD6BWP30P140LVT U1192 ( .I(n3461), .Z(o_data_bus[827]) );
  BUFFD6BWP30P140LVT U1193 ( .I(n3462), .Z(o_data_bus[826]) );
  BUFFD6BWP30P140LVT U1194 ( .I(n3463), .Z(o_data_bus[825]) );
  BUFFD6BWP30P140LVT U1195 ( .I(n3464), .Z(o_data_bus[824]) );
  BUFFD6BWP30P140LVT U1196 ( .I(n3465), .Z(o_data_bus[823]) );
  BUFFD6BWP30P140LVT U1197 ( .I(n3466), .Z(o_data_bus[822]) );
  BUFFD6BWP30P140LVT U1198 ( .I(n3467), .Z(o_data_bus[821]) );
  BUFFD6BWP30P140LVT U1199 ( .I(n3468), .Z(o_data_bus[820]) );
  BUFFD6BWP30P140LVT U1200 ( .I(n3401), .Z(o_data_bus[887]) );
  BUFFD6BWP30P140LVT U1201 ( .I(n3469), .Z(o_data_bus[819]) );
  BUFFD6BWP30P140LVT U1202 ( .I(n3470), .Z(o_data_bus[818]) );
  BUFFD6BWP30P140LVT U1203 ( .I(n3471), .Z(o_data_bus[817]) );
  BUFFD6BWP30P140LVT U1204 ( .I(n3472), .Z(o_data_bus[816]) );
  BUFFD6BWP30P140LVT U1205 ( .I(n3473), .Z(o_data_bus[815]) );
  BUFFD6BWP30P140LVT U1206 ( .I(n3474), .Z(o_data_bus[814]) );
  BUFFD6BWP30P140LVT U1207 ( .I(n3475), .Z(o_data_bus[813]) );
  BUFFD6BWP30P140LVT U1208 ( .I(n3476), .Z(o_data_bus[812]) );
  BUFFD6BWP30P140LVT U1209 ( .I(n3477), .Z(o_data_bus[811]) );
  BUFFD6BWP30P140LVT U1210 ( .I(n3478), .Z(o_data_bus[810]) );
  BUFFD6BWP30P140LVT U1211 ( .I(n3479), .Z(o_data_bus[809]) );
  BUFFD6BWP30P140LVT U1212 ( .I(n3480), .Z(o_data_bus[808]) );
  BUFFD6BWP30P140LVT U1213 ( .I(n3481), .Z(o_data_bus[807]) );
  BUFFD6BWP30P140LVT U1214 ( .I(n3482), .Z(o_data_bus[806]) );
  BUFFD6BWP30P140LVT U1215 ( .I(n3483), .Z(o_data_bus[805]) );
  BUFFD6BWP30P140LVT U1216 ( .I(n3484), .Z(o_data_bus[804]) );
  BUFFD6BWP30P140LVT U1217 ( .I(n3485), .Z(o_data_bus[803]) );
  BUFFD6BWP30P140LVT U1218 ( .I(n3486), .Z(o_data_bus[802]) );
  BUFFD6BWP30P140LVT U1219 ( .I(n3487), .Z(o_data_bus[801]) );
  BUFFD6BWP30P140LVT U1220 ( .I(n3488), .Z(o_data_bus[800]) );
  BUFFD6BWP30P140LVT U1221 ( .I(n3489), .Z(o_data_bus[799]) );
  BUFFD6BWP30P140LVT U1222 ( .I(n3490), .Z(o_data_bus[798]) );
  BUFFD6BWP30P140LVT U1223 ( .I(n3491), .Z(o_data_bus[797]) );
  BUFFD6BWP30P140LVT U1224 ( .I(n3492), .Z(o_data_bus[796]) );
  BUFFD6BWP30P140LVT U1225 ( .I(n3493), .Z(o_data_bus[795]) );
  BUFFD6BWP30P140LVT U1226 ( .I(n3494), .Z(o_data_bus[794]) );
  BUFFD6BWP30P140LVT U1227 ( .I(n3495), .Z(o_data_bus[793]) );
  BUFFD6BWP30P140LVT U1228 ( .I(n3496), .Z(o_data_bus[792]) );
  BUFFD6BWP30P140LVT U1229 ( .I(n3497), .Z(o_data_bus[791]) );
  BUFFD6BWP30P140LVT U1230 ( .I(n3498), .Z(o_data_bus[790]) );
  BUFFD6BWP30P140LVT U1231 ( .I(n3499), .Z(o_data_bus[789]) );
  BUFFD6BWP30P140LVT U1232 ( .I(n3500), .Z(o_data_bus[788]) );
  BUFFD6BWP30P140LVT U1233 ( .I(n3501), .Z(o_data_bus[787]) );
  BUFFD6BWP30P140LVT U1234 ( .I(n3502), .Z(o_data_bus[786]) );
  BUFFD6BWP30P140LVT U1235 ( .I(n3503), .Z(o_data_bus[785]) );
  BUFFD6BWP30P140LVT U1236 ( .I(n3504), .Z(o_data_bus[784]) );
  BUFFD6BWP30P140LVT U1237 ( .I(n3505), .Z(o_data_bus[783]) );
  BUFFD6BWP30P140LVT U1238 ( .I(n3506), .Z(o_data_bus[782]) );
  BUFFD6BWP30P140LVT U1239 ( .I(n3507), .Z(o_data_bus[781]) );
  BUFFD6BWP30P140LVT U1240 ( .I(n3508), .Z(o_data_bus[780]) );
  BUFFD6BWP30P140LVT U1241 ( .I(n3509), .Z(o_data_bus[779]) );
  BUFFD6BWP30P140LVT U1242 ( .I(n3510), .Z(o_data_bus[778]) );
  BUFFD6BWP30P140LVT U1243 ( .I(n3511), .Z(o_data_bus[777]) );
  BUFFD6BWP30P140LVT U1244 ( .I(n3512), .Z(o_data_bus[776]) );
  BUFFD6BWP30P140LVT U1245 ( .I(n3513), .Z(o_data_bus[775]) );
  BUFFD6BWP30P140LVT U1246 ( .I(n3514), .Z(o_data_bus[774]) );
  BUFFD6BWP30P140LVT U1247 ( .I(n3515), .Z(o_data_bus[773]) );
  BUFFD6BWP30P140LVT U1248 ( .I(n3516), .Z(o_data_bus[772]) );
  BUFFD6BWP30P140LVT U1249 ( .I(n3517), .Z(o_data_bus[771]) );
  BUFFD6BWP30P140LVT U1250 ( .I(n3518), .Z(o_data_bus[770]) );
  BUFFD6BWP30P140LVT U1251 ( .I(n3519), .Z(o_data_bus[769]) );
  BUFFD6BWP30P140LVT U1252 ( .I(n3520), .Z(o_data_bus[768]) );
  BUFFD6BWP30P140LVT U1253 ( .I(n3521), .Z(o_data_bus[767]) );
  BUFFD6BWP30P140LVT U1254 ( .I(n3522), .Z(o_data_bus[766]) );
  BUFFD6BWP30P140LVT U1255 ( .I(n3523), .Z(o_data_bus[765]) );
  BUFFD6BWP30P140LVT U1256 ( .I(n3524), .Z(o_data_bus[764]) );
  BUFFD6BWP30P140LVT U1257 ( .I(n3525), .Z(o_data_bus[763]) );
  BUFFD6BWP30P140LVT U1258 ( .I(n3526), .Z(o_data_bus[762]) );
  BUFFD6BWP30P140LVT U1259 ( .I(n3527), .Z(o_data_bus[761]) );
  BUFFD6BWP30P140LVT U1260 ( .I(n3528), .Z(o_data_bus[760]) );
  BUFFD6BWP30P140LVT U1261 ( .I(n3529), .Z(o_data_bus[759]) );
  BUFFD6BWP30P140LVT U1262 ( .I(n3530), .Z(o_data_bus[758]) );
  BUFFD6BWP30P140LVT U1263 ( .I(n3531), .Z(o_data_bus[757]) );
  BUFFD6BWP30P140LVT U1264 ( .I(n3532), .Z(o_data_bus[756]) );
  BUFFD6BWP30P140LVT U1265 ( .I(n3533), .Z(o_data_bus[755]) );
  BUFFD6BWP30P140LVT U1266 ( .I(n3534), .Z(o_data_bus[754]) );
  BUFFD6BWP30P140LVT U1267 ( .I(n3535), .Z(o_data_bus[753]) );
  BUFFD6BWP30P140LVT U1268 ( .I(n3536), .Z(o_data_bus[752]) );
  BUFFD6BWP30P140LVT U1269 ( .I(n3267), .Z(o_data_bus[1021]) );
  BUFFD6BWP30P140LVT U1270 ( .I(n3268), .Z(o_data_bus[1020]) );
  BUFFD6BWP30P140LVT U1271 ( .I(n3269), .Z(o_data_bus[1019]) );
  BUFFD6BWP30P140LVT U1272 ( .I(n3270), .Z(o_data_bus[1018]) );
  BUFFD6BWP30P140LVT U1273 ( .I(n3271), .Z(o_data_bus[1017]) );
  BUFFD6BWP30P140LVT U1274 ( .I(n3272), .Z(o_data_bus[1016]) );
  BUFFD6BWP30P140LVT U1275 ( .I(n3273), .Z(o_data_bus[1015]) );
  BUFFD6BWP30P140LVT U1276 ( .I(n3274), .Z(o_data_bus[1014]) );
  BUFFD6BWP30P140LVT U1277 ( .I(n3275), .Z(o_data_bus[1013]) );
  BUFFD6BWP30P140LVT U1278 ( .I(n3276), .Z(o_data_bus[1012]) );
  BUFFD6BWP30P140LVT U1279 ( .I(n3277), .Z(o_data_bus[1011]) );
  BUFFD6BWP30P140LVT U1280 ( .I(n3278), .Z(o_data_bus[1010]) );
  BUFFD6BWP30P140LVT U1281 ( .I(n3279), .Z(o_data_bus[1009]) );
  BUFFD6BWP30P140LVT U1282 ( .I(n3280), .Z(o_data_bus[1008]) );
  BUFFD6BWP30P140LVT U1283 ( .I(n3281), .Z(o_data_bus[1007]) );
  BUFFD6BWP30P140LVT U1284 ( .I(n3282), .Z(o_data_bus[1006]) );
  BUFFD6BWP30P140LVT U1285 ( .I(n3283), .Z(o_data_bus[1005]) );
  BUFFD6BWP30P140LVT U1286 ( .I(n3284), .Z(o_data_bus[1004]) );
  BUFFD6BWP30P140LVT U1287 ( .I(n3285), .Z(o_data_bus[1003]) );
  BUFFD6BWP30P140LVT U1288 ( .I(n3286), .Z(o_data_bus[1002]) );
  BUFFD6BWP30P140LVT U1289 ( .I(n3287), .Z(o_data_bus[1001]) );
  BUFFD6BWP30P140LVT U1290 ( .I(n3288), .Z(o_data_bus[1000]) );
  BUFFD6BWP30P140LVT U1291 ( .I(n3289), .Z(o_data_bus[999]) );
  BUFFD6BWP30P140LVT U1292 ( .I(n3290), .Z(o_data_bus[998]) );
  BUFFD6BWP30P140LVT U1293 ( .I(n3291), .Z(o_data_bus[997]) );
  BUFFD6BWP30P140LVT U1294 ( .I(n3292), .Z(o_data_bus[996]) );
  BUFFD6BWP30P140LVT U1295 ( .I(n3293), .Z(o_data_bus[995]) );
  BUFFD6BWP30P140LVT U1296 ( .I(n3294), .Z(o_data_bus[994]) );
  BUFFD6BWP30P140LVT U1297 ( .I(n3295), .Z(o_data_bus[993]) );
  BUFFD6BWP30P140LVT U1298 ( .I(n3296), .Z(o_data_bus[992]) );
  BUFFD6BWP30P140LVT U1299 ( .I(n3297), .Z(o_data_bus[991]) );
  BUFFD6BWP30P140LVT U1300 ( .I(n3298), .Z(o_data_bus[990]) );
  BUFFD6BWP30P140LVT U1301 ( .I(n3299), .Z(o_data_bus[989]) );
  BUFFD6BWP30P140LVT U1302 ( .I(n3300), .Z(o_data_bus[988]) );
  BUFFD6BWP30P140LVT U1303 ( .I(n3301), .Z(o_data_bus[987]) );
  BUFFD6BWP30P140LVT U1304 ( .I(n3302), .Z(o_data_bus[986]) );
  BUFFD6BWP30P140LVT U1305 ( .I(n3303), .Z(o_data_bus[985]) );
  BUFFD6BWP30P140LVT U1306 ( .I(n3304), .Z(o_data_bus[984]) );
  BUFFD6BWP30P140LVT U1307 ( .I(n3305), .Z(o_data_bus[983]) );
  BUFFD6BWP30P140LVT U1308 ( .I(n3306), .Z(o_data_bus[982]) );
  BUFFD6BWP30P140LVT U1309 ( .I(n3307), .Z(o_data_bus[981]) );
  BUFFD6BWP30P140LVT U1310 ( .I(n3308), .Z(o_data_bus[980]) );
  BUFFD6BWP30P140LVT U1311 ( .I(n3309), .Z(o_data_bus[979]) );
  BUFFD6BWP30P140LVT U1312 ( .I(n3310), .Z(o_data_bus[978]) );
  BUFFD6BWP30P140LVT U1313 ( .I(n3311), .Z(o_data_bus[977]) );
  BUFFD6BWP30P140LVT U1314 ( .I(n3312), .Z(o_data_bus[976]) );
  BUFFD6BWP30P140LVT U1315 ( .I(n3313), .Z(o_data_bus[975]) );
  BUFFD6BWP30P140LVT U1316 ( .I(n3314), .Z(o_data_bus[974]) );
  BUFFD6BWP30P140LVT U1317 ( .I(n3315), .Z(o_data_bus[973]) );
  BUFFD6BWP30P140LVT U1318 ( .I(n3316), .Z(o_data_bus[972]) );
  BUFFD6BWP30P140LVT U1319 ( .I(n3317), .Z(o_data_bus[971]) );
  BUFFD6BWP30P140LVT U1320 ( .I(n3318), .Z(o_data_bus[970]) );
  BUFFD6BWP30P140LVT U1321 ( .I(n3319), .Z(o_data_bus[969]) );
  BUFFD6BWP30P140LVT U1322 ( .I(n3320), .Z(o_data_bus[968]) );
  BUFFD6BWP30P140LVT U1323 ( .I(n3321), .Z(o_data_bus[967]) );
  BUFFD6BWP30P140LVT U1324 ( .I(n3322), .Z(o_data_bus[966]) );
  BUFFD6BWP30P140LVT U1325 ( .I(n3323), .Z(o_data_bus[965]) );
  BUFFD6BWP30P140LVT U1326 ( .I(n3324), .Z(o_data_bus[964]) );
  BUFFD6BWP30P140LVT U1327 ( .I(n3325), .Z(o_data_bus[963]) );
  BUFFD6BWP30P140LVT U1328 ( .I(n3326), .Z(o_data_bus[962]) );
  BUFFD6BWP30P140LVT U1329 ( .I(n3327), .Z(o_data_bus[961]) );
  BUFFD6BWP30P140LVT U1330 ( .I(n3328), .Z(o_data_bus[960]) );
  BUFFD6BWP30P140LVT U1331 ( .I(n3329), .Z(o_data_bus[959]) );
  BUFFD6BWP30P140LVT U1332 ( .I(n3330), .Z(o_data_bus[958]) );
  BUFFD6BWP30P140LVT U1333 ( .I(n3331), .Z(o_data_bus[957]) );
  BUFFD6BWP30P140LVT U1334 ( .I(n3332), .Z(o_data_bus[956]) );
  BUFFD6BWP30P140LVT U1335 ( .I(n3333), .Z(o_data_bus[955]) );
  BUFFD6BWP30P140LVT U1336 ( .I(n3266), .Z(o_data_bus[1022]) );
  BUFFD6BWP30P140LVT U1337 ( .I(n3334), .Z(o_data_bus[954]) );
  BUFFD6BWP30P140LVT U1338 ( .I(n3335), .Z(o_data_bus[953]) );
  BUFFD6BWP30P140LVT U1339 ( .I(n3336), .Z(o_data_bus[952]) );
  BUFFD6BWP30P140LVT U1340 ( .I(n3337), .Z(o_data_bus[951]) );
  BUFFD6BWP30P140LVT U1341 ( .I(n3338), .Z(o_data_bus[950]) );
  BUFFD6BWP30P140LVT U1342 ( .I(n3339), .Z(o_data_bus[949]) );
  BUFFD6BWP30P140LVT U1343 ( .I(n3340), .Z(o_data_bus[948]) );
  BUFFD6BWP30P140LVT U1344 ( .I(n3341), .Z(o_data_bus[947]) );
  BUFFD6BWP30P140LVT U1345 ( .I(n3342), .Z(o_data_bus[946]) );
  BUFFD6BWP30P140LVT U1346 ( .I(n3343), .Z(o_data_bus[945]) );
  BUFFD6BWP30P140LVT U1347 ( .I(n3344), .Z(o_data_bus[944]) );
  BUFFD6BWP30P140LVT U1348 ( .I(n3345), .Z(o_data_bus[943]) );
  BUFFD6BWP30P140LVT U1349 ( .I(n3346), .Z(o_data_bus[942]) );
  BUFFD6BWP30P140LVT U1350 ( .I(n3347), .Z(o_data_bus[941]) );
  BUFFD6BWP30P140LVT U1351 ( .I(n3348), .Z(o_data_bus[940]) );
  BUFFD6BWP30P140LVT U1352 ( .I(n3349), .Z(o_data_bus[939]) );
  BUFFD6BWP30P140LVT U1353 ( .I(n3350), .Z(o_data_bus[938]) );
  BUFFD6BWP30P140LVT U1354 ( .I(n3351), .Z(o_data_bus[937]) );
  BUFFD6BWP30P140LVT U1355 ( .I(n3352), .Z(o_data_bus[936]) );
  BUFFD6BWP30P140LVT U1356 ( .I(n3353), .Z(o_data_bus[935]) );
  BUFFD6BWP30P140LVT U1357 ( .I(n3354), .Z(o_data_bus[934]) );
  BUFFD6BWP30P140LVT U1358 ( .I(n3355), .Z(o_data_bus[933]) );
  BUFFD6BWP30P140LVT U1359 ( .I(n3356), .Z(o_data_bus[932]) );
  BUFFD6BWP30P140LVT U1360 ( .I(n3357), .Z(o_data_bus[931]) );
  BUFFD6BWP30P140LVT U1361 ( .I(n3358), .Z(o_data_bus[930]) );
  BUFFD6BWP30P140LVT U1362 ( .I(n3359), .Z(o_data_bus[929]) );
  BUFFD6BWP30P140LVT U1363 ( .I(n3360), .Z(o_data_bus[928]) );
  BUFFD6BWP30P140LVT U1364 ( .I(n3361), .Z(o_data_bus[927]) );
  BUFFD6BWP30P140LVT U1365 ( .I(n3362), .Z(o_data_bus[926]) );
  BUFFD6BWP30P140LVT U1366 ( .I(n3363), .Z(o_data_bus[925]) );
  BUFFD6BWP30P140LVT U1367 ( .I(n3364), .Z(o_data_bus[924]) );
  BUFFD6BWP30P140LVT U1368 ( .I(n3365), .Z(o_data_bus[923]) );
  BUFFD6BWP30P140LVT U1369 ( .I(n3366), .Z(o_data_bus[922]) );
  BUFFD6BWP30P140LVT U1370 ( .I(n3367), .Z(o_data_bus[921]) );
  BUFFD6BWP30P140LVT U1371 ( .I(n3368), .Z(o_data_bus[920]) );
  BUFFD6BWP30P140LVT U1372 ( .I(n3369), .Z(o_data_bus[919]) );
  BUFFD6BWP30P140LVT U1373 ( .I(n3370), .Z(o_data_bus[918]) );
  BUFFD6BWP30P140LVT U1374 ( .I(n3371), .Z(o_data_bus[917]) );
  BUFFD6BWP30P140LVT U1375 ( .I(n3372), .Z(o_data_bus[916]) );
  BUFFD6BWP30P140LVT U1376 ( .I(n3373), .Z(o_data_bus[915]) );
  BUFFD6BWP30P140LVT U1377 ( .I(n3374), .Z(o_data_bus[914]) );
  BUFFD6BWP30P140LVT U1378 ( .I(n3375), .Z(o_data_bus[913]) );
  BUFFD6BWP30P140LVT U1379 ( .I(n3376), .Z(o_data_bus[912]) );
  BUFFD6BWP30P140LVT U1380 ( .I(n3377), .Z(o_data_bus[911]) );
  BUFFD6BWP30P140LVT U1381 ( .I(n3378), .Z(o_data_bus[910]) );
  BUFFD6BWP30P140LVT U1382 ( .I(n3379), .Z(o_data_bus[909]) );
  BUFFD6BWP30P140LVT U1383 ( .I(n3380), .Z(o_data_bus[908]) );
  BUFFD6BWP30P140LVT U1384 ( .I(n3381), .Z(o_data_bus[907]) );
  BUFFD6BWP30P140LVT U1385 ( .I(n3382), .Z(o_data_bus[906]) );
  BUFFD6BWP30P140LVT U1386 ( .I(n3383), .Z(o_data_bus[905]) );
  BUFFD6BWP30P140LVT U1387 ( .I(n3384), .Z(o_data_bus[904]) );
  BUFFD6BWP30P140LVT U1388 ( .I(n3385), .Z(o_data_bus[903]) );
  BUFFD6BWP30P140LVT U1389 ( .I(n3386), .Z(o_data_bus[902]) );
  BUFFD6BWP30P140LVT U1390 ( .I(n3387), .Z(o_data_bus[901]) );
  BUFFD6BWP30P140LVT U1391 ( .I(n3388), .Z(o_data_bus[900]) );
  BUFFD6BWP30P140LVT U1392 ( .I(n3389), .Z(o_data_bus[899]) );
  BUFFD6BWP30P140LVT U1393 ( .I(n3390), .Z(o_data_bus[898]) );
  BUFFD6BWP30P140LVT U1394 ( .I(n3391), .Z(o_data_bus[897]) );
  BUFFD6BWP30P140LVT U1395 ( .I(n3392), .Z(o_data_bus[896]) );
  BUFFD6BWP30P140LVT U1396 ( .I(n3393), .Z(o_data_bus[895]) );
  BUFFD6BWP30P140LVT U1397 ( .I(n3394), .Z(o_data_bus[894]) );
  BUFFD6BWP30P140LVT U1398 ( .I(n3395), .Z(o_data_bus[893]) );
  BUFFD6BWP30P140LVT U1399 ( .I(n3396), .Z(o_data_bus[892]) );
  BUFFD6BWP30P140LVT U1400 ( .I(n3397), .Z(o_data_bus[891]) );
  BUFFD6BWP30P140LVT U1401 ( .I(n3398), .Z(o_data_bus[890]) );
  BUFFD6BWP30P140LVT U1402 ( .I(n3399), .Z(o_data_bus[889]) );
  BUFFD6BWP30P140LVT U1403 ( .I(n3400), .Z(o_data_bus[888]) );
  BUFFD6BWP30P140LVT U1404 ( .I(n3537), .Z(o_data_bus[751]) );
  BUFFD6BWP30P140LVT U1405 ( .I(n3674), .Z(o_data_bus[614]) );
  BUFFD6BWP30P140LVT U1406 ( .I(n3675), .Z(o_data_bus[613]) );
  BUFFD6BWP30P140LVT U1407 ( .I(n3676), .Z(o_data_bus[612]) );
  BUFFD6BWP30P140LVT U1408 ( .I(n3677), .Z(o_data_bus[611]) );
  BUFFD6BWP30P140LVT U1409 ( .I(n3678), .Z(o_data_bus[610]) );
  BUFFD6BWP30P140LVT U1410 ( .I(n3679), .Z(o_data_bus[609]) );
  BUFFD6BWP30P140LVT U1411 ( .I(n3680), .Z(o_data_bus[608]) );
  BUFFD6BWP30P140LVT U1412 ( .I(n3681), .Z(o_data_bus[607]) );
  BUFFD6BWP30P140LVT U1413 ( .I(n3682), .Z(o_data_bus[606]) );
  BUFFD6BWP30P140LVT U1414 ( .I(n3683), .Z(o_data_bus[605]) );
  BUFFD6BWP30P140LVT U1415 ( .I(n3684), .Z(o_data_bus[604]) );
  BUFFD6BWP30P140LVT U1416 ( .I(n3685), .Z(o_data_bus[603]) );
  BUFFD6BWP30P140LVT U1417 ( .I(n3686), .Z(o_data_bus[602]) );
  BUFFD6BWP30P140LVT U1418 ( .I(n3687), .Z(o_data_bus[601]) );
  BUFFD6BWP30P140LVT U1419 ( .I(n3688), .Z(o_data_bus[600]) );
  BUFFD6BWP30P140LVT U1420 ( .I(n3689), .Z(o_data_bus[599]) );
  BUFFD6BWP30P140LVT U1421 ( .I(n3690), .Z(o_data_bus[598]) );
  BUFFD6BWP30P140LVT U1422 ( .I(n3691), .Z(o_data_bus[597]) );
  BUFFD6BWP30P140LVT U1423 ( .I(n3692), .Z(o_data_bus[596]) );
  BUFFD6BWP30P140LVT U1424 ( .I(n3693), .Z(o_data_bus[595]) );
  BUFFD6BWP30P140LVT U1425 ( .I(n3694), .Z(o_data_bus[594]) );
  BUFFD6BWP30P140LVT U1426 ( .I(n3695), .Z(o_data_bus[593]) );
  BUFFD6BWP30P140LVT U1427 ( .I(n3696), .Z(o_data_bus[592]) );
  BUFFD6BWP30P140LVT U1428 ( .I(n3697), .Z(o_data_bus[591]) );
  BUFFD6BWP30P140LVT U1429 ( .I(n3698), .Z(o_data_bus[590]) );
  BUFFD6BWP30P140LVT U1430 ( .I(n3699), .Z(o_data_bus[589]) );
  BUFFD6BWP30P140LVT U1431 ( .I(n3700), .Z(o_data_bus[588]) );
  BUFFD6BWP30P140LVT U1432 ( .I(n3701), .Z(o_data_bus[587]) );
  BUFFD6BWP30P140LVT U1433 ( .I(n3702), .Z(o_data_bus[586]) );
  BUFFD6BWP30P140LVT U1434 ( .I(n3703), .Z(o_data_bus[585]) );
  BUFFD6BWP30P140LVT U1435 ( .I(n3704), .Z(o_data_bus[584]) );
  BUFFD6BWP30P140LVT U1436 ( .I(n3705), .Z(o_data_bus[583]) );
  BUFFD6BWP30P140LVT U1437 ( .I(n3706), .Z(o_data_bus[582]) );
  BUFFD6BWP30P140LVT U1438 ( .I(n3707), .Z(o_data_bus[581]) );
  BUFFD6BWP30P140LVT U1439 ( .I(n3708), .Z(o_data_bus[580]) );
  BUFFD6BWP30P140LVT U1440 ( .I(n3709), .Z(o_data_bus[579]) );
  BUFFD6BWP30P140LVT U1441 ( .I(n3710), .Z(o_data_bus[578]) );
  BUFFD6BWP30P140LVT U1442 ( .I(n3711), .Z(o_data_bus[577]) );
  BUFFD6BWP30P140LVT U1443 ( .I(n3712), .Z(o_data_bus[576]) );
  BUFFD6BWP30P140LVT U1444 ( .I(n3713), .Z(o_data_bus[575]) );
  BUFFD6BWP30P140LVT U1445 ( .I(n3714), .Z(o_data_bus[574]) );
  BUFFD6BWP30P140LVT U1446 ( .I(n3715), .Z(o_data_bus[573]) );
  BUFFD6BWP30P140LVT U1447 ( .I(n3716), .Z(o_data_bus[572]) );
  BUFFD6BWP30P140LVT U1448 ( .I(n3717), .Z(o_data_bus[571]) );
  BUFFD6BWP30P140LVT U1449 ( .I(n3718), .Z(o_data_bus[570]) );
  BUFFD6BWP30P140LVT U1450 ( .I(n3719), .Z(o_data_bus[569]) );
  BUFFD6BWP30P140LVT U1451 ( .I(n3720), .Z(o_data_bus[568]) );
  BUFFD6BWP30P140LVT U1452 ( .I(n3721), .Z(o_data_bus[567]) );
  BUFFD6BWP30P140LVT U1453 ( .I(n3722), .Z(o_data_bus[566]) );
  BUFFD6BWP30P140LVT U1454 ( .I(n3723), .Z(o_data_bus[565]) );
  BUFFD6BWP30P140LVT U1455 ( .I(n3724), .Z(o_data_bus[564]) );
  BUFFD6BWP30P140LVT U1456 ( .I(n3725), .Z(o_data_bus[563]) );
  BUFFD6BWP30P140LVT U1457 ( .I(n3726), .Z(o_data_bus[562]) );
  BUFFD6BWP30P140LVT U1458 ( .I(n3727), .Z(o_data_bus[561]) );
  BUFFD6BWP30P140LVT U1459 ( .I(n3728), .Z(o_data_bus[560]) );
  BUFFD6BWP30P140LVT U1460 ( .I(n3729), .Z(o_data_bus[559]) );
  BUFFD6BWP30P140LVT U1461 ( .I(n3730), .Z(o_data_bus[558]) );
  BUFFD6BWP30P140LVT U1462 ( .I(n3731), .Z(o_data_bus[557]) );
  BUFFD6BWP30P140LVT U1463 ( .I(n3732), .Z(o_data_bus[556]) );
  BUFFD6BWP30P140LVT U1464 ( .I(n3733), .Z(o_data_bus[555]) );
  BUFFD6BWP30P140LVT U1465 ( .I(n3734), .Z(o_data_bus[554]) );
  BUFFD6BWP30P140LVT U1466 ( .I(n3735), .Z(o_data_bus[553]) );
  BUFFD6BWP30P140LVT U1467 ( .I(n3736), .Z(o_data_bus[552]) );
  BUFFD6BWP30P140LVT U1468 ( .I(n3737), .Z(o_data_bus[551]) );
  BUFFD6BWP30P140LVT U1469 ( .I(n3738), .Z(o_data_bus[550]) );
  BUFFD6BWP30P140LVT U1470 ( .I(n3739), .Z(o_data_bus[549]) );
  BUFFD6BWP30P140LVT U1471 ( .I(n3740), .Z(o_data_bus[548]) );
  BUFFD6BWP30P140LVT U1472 ( .I(n3673), .Z(o_data_bus[615]) );
  BUFFD6BWP30P140LVT U1473 ( .I(n3741), .Z(o_data_bus[547]) );
  BUFFD6BWP30P140LVT U1474 ( .I(n3742), .Z(o_data_bus[546]) );
  BUFFD6BWP30P140LVT U1475 ( .I(n3743), .Z(o_data_bus[545]) );
  BUFFD6BWP30P140LVT U1476 ( .I(n3744), .Z(o_data_bus[544]) );
  BUFFD6BWP30P140LVT U1477 ( .I(n3745), .Z(o_data_bus[543]) );
  BUFFD6BWP30P140LVT U1478 ( .I(n3746), .Z(o_data_bus[542]) );
  BUFFD6BWP30P140LVT U1479 ( .I(n3747), .Z(o_data_bus[541]) );
  BUFFD6BWP30P140LVT U1480 ( .I(n3748), .Z(o_data_bus[540]) );
  BUFFD6BWP30P140LVT U1481 ( .I(n3749), .Z(o_data_bus[539]) );
  BUFFD6BWP30P140LVT U1482 ( .I(n3750), .Z(o_data_bus[538]) );
  BUFFD6BWP30P140LVT U1483 ( .I(n3751), .Z(o_data_bus[537]) );
  BUFFD6BWP30P140LVT U1484 ( .I(n3752), .Z(o_data_bus[536]) );
  BUFFD6BWP30P140LVT U1485 ( .I(n3753), .Z(o_data_bus[535]) );
  BUFFD6BWP30P140LVT U1486 ( .I(n3754), .Z(o_data_bus[534]) );
  BUFFD6BWP30P140LVT U1487 ( .I(n3755), .Z(o_data_bus[533]) );
  BUFFD6BWP30P140LVT U1488 ( .I(n3756), .Z(o_data_bus[532]) );
  BUFFD6BWP30P140LVT U1489 ( .I(n3757), .Z(o_data_bus[531]) );
  BUFFD6BWP30P140LVT U1490 ( .I(n3758), .Z(o_data_bus[530]) );
  BUFFD6BWP30P140LVT U1491 ( .I(n3759), .Z(o_data_bus[529]) );
  BUFFD6BWP30P140LVT U1492 ( .I(n3760), .Z(o_data_bus[528]) );
  BUFFD6BWP30P140LVT U1493 ( .I(n3761), .Z(o_data_bus[527]) );
  BUFFD6BWP30P140LVT U1494 ( .I(n3762), .Z(o_data_bus[526]) );
  BUFFD6BWP30P140LVT U1495 ( .I(n3763), .Z(o_data_bus[525]) );
  BUFFD6BWP30P140LVT U1496 ( .I(n3764), .Z(o_data_bus[524]) );
  BUFFD6BWP30P140LVT U1497 ( .I(n3765), .Z(o_data_bus[523]) );
  BUFFD6BWP30P140LVT U1498 ( .I(n3766), .Z(o_data_bus[522]) );
  BUFFD6BWP30P140LVT U1499 ( .I(n3767), .Z(o_data_bus[521]) );
  BUFFD6BWP30P140LVT U1500 ( .I(n3768), .Z(o_data_bus[520]) );
  BUFFD6BWP30P140LVT U1501 ( .I(n3769), .Z(o_data_bus[519]) );
  BUFFD6BWP30P140LVT U1502 ( .I(n3770), .Z(o_data_bus[518]) );
  BUFFD6BWP30P140LVT U1503 ( .I(n3771), .Z(o_data_bus[517]) );
  BUFFD6BWP30P140LVT U1504 ( .I(n3772), .Z(o_data_bus[516]) );
  BUFFD6BWP30P140LVT U1505 ( .I(n3773), .Z(o_data_bus[515]) );
  BUFFD6BWP30P140LVT U1506 ( .I(n3774), .Z(o_data_bus[514]) );
  BUFFD6BWP30P140LVT U1507 ( .I(n3775), .Z(o_data_bus[513]) );
  BUFFD6BWP30P140LVT U1508 ( .I(n3776), .Z(o_data_bus[512]) );
  BUFFD6BWP30P140LVT U1509 ( .I(n3777), .Z(o_data_bus[511]) );
  BUFFD6BWP30P140LVT U1510 ( .I(n3778), .Z(o_data_bus[510]) );
  BUFFD6BWP30P140LVT U1511 ( .I(n3779), .Z(o_data_bus[509]) );
  BUFFD6BWP30P140LVT U1512 ( .I(n3780), .Z(o_data_bus[508]) );
  BUFFD6BWP30P140LVT U1513 ( .I(n3781), .Z(o_data_bus[507]) );
  BUFFD6BWP30P140LVT U1514 ( .I(n3782), .Z(o_data_bus[506]) );
  BUFFD6BWP30P140LVT U1515 ( .I(n3783), .Z(o_data_bus[505]) );
  BUFFD6BWP30P140LVT U1516 ( .I(n3784), .Z(o_data_bus[504]) );
  BUFFD6BWP30P140LVT U1517 ( .I(n3785), .Z(o_data_bus[503]) );
  BUFFD6BWP30P140LVT U1518 ( .I(n3786), .Z(o_data_bus[502]) );
  BUFFD6BWP30P140LVT U1519 ( .I(n3787), .Z(o_data_bus[501]) );
  BUFFD6BWP30P140LVT U1520 ( .I(n3788), .Z(o_data_bus[500]) );
  BUFFD6BWP30P140LVT U1521 ( .I(n3789), .Z(o_data_bus[499]) );
  BUFFD6BWP30P140LVT U1522 ( .I(n3790), .Z(o_data_bus[498]) );
  BUFFD6BWP30P140LVT U1523 ( .I(n3791), .Z(o_data_bus[497]) );
  BUFFD6BWP30P140LVT U1524 ( .I(n3792), .Z(o_data_bus[496]) );
  BUFFD6BWP30P140LVT U1525 ( .I(n3793), .Z(o_data_bus[495]) );
  BUFFD6BWP30P140LVT U1526 ( .I(n3794), .Z(o_data_bus[494]) );
  BUFFD6BWP30P140LVT U1527 ( .I(n3795), .Z(o_data_bus[493]) );
  BUFFD6BWP30P140LVT U1528 ( .I(n3796), .Z(o_data_bus[492]) );
  BUFFD6BWP30P140LVT U1529 ( .I(n3797), .Z(o_data_bus[491]) );
  BUFFD6BWP30P140LVT U1530 ( .I(n3798), .Z(o_data_bus[490]) );
  BUFFD6BWP30P140LVT U1531 ( .I(n3799), .Z(o_data_bus[489]) );
  BUFFD6BWP30P140LVT U1532 ( .I(n3800), .Z(o_data_bus[488]) );
  BUFFD6BWP30P140LVT U1533 ( .I(n3801), .Z(o_data_bus[487]) );
  BUFFD6BWP30P140LVT U1534 ( .I(n3802), .Z(o_data_bus[486]) );
  BUFFD6BWP30P140LVT U1535 ( .I(n3803), .Z(o_data_bus[485]) );
  BUFFD6BWP30P140LVT U1536 ( .I(n3804), .Z(o_data_bus[484]) );
  BUFFD6BWP30P140LVT U1537 ( .I(n3805), .Z(o_data_bus[483]) );
  BUFFD6BWP30P140LVT U1538 ( .I(n3806), .Z(o_data_bus[482]) );
  BUFFD6BWP30P140LVT U1539 ( .I(n3807), .Z(o_data_bus[481]) );
  BUFFD6BWP30P140LVT U1540 ( .I(n3672), .Z(o_data_bus[616]) );
  BUFFD6BWP30P140LVT U1541 ( .I(n3538), .Z(o_data_bus[750]) );
  BUFFD6BWP30P140LVT U1542 ( .I(n3539), .Z(o_data_bus[749]) );
  BUFFD6BWP30P140LVT U1543 ( .I(n3540), .Z(o_data_bus[748]) );
  BUFFD6BWP30P140LVT U1544 ( .I(n3541), .Z(o_data_bus[747]) );
  BUFFD6BWP30P140LVT U1545 ( .I(n3542), .Z(o_data_bus[746]) );
  BUFFD6BWP30P140LVT U1546 ( .I(n3543), .Z(o_data_bus[745]) );
  BUFFD6BWP30P140LVT U1547 ( .I(n3544), .Z(o_data_bus[744]) );
  BUFFD6BWP30P140LVT U1548 ( .I(n3545), .Z(o_data_bus[743]) );
  BUFFD6BWP30P140LVT U1549 ( .I(n3546), .Z(o_data_bus[742]) );
  BUFFD6BWP30P140LVT U1550 ( .I(n3547), .Z(o_data_bus[741]) );
  BUFFD6BWP30P140LVT U1551 ( .I(n3548), .Z(o_data_bus[740]) );
  BUFFD6BWP30P140LVT U1552 ( .I(n3549), .Z(o_data_bus[739]) );
  BUFFD6BWP30P140LVT U1553 ( .I(n3550), .Z(o_data_bus[738]) );
  BUFFD6BWP30P140LVT U1554 ( .I(n3551), .Z(o_data_bus[737]) );
  BUFFD6BWP30P140LVT U1555 ( .I(n3552), .Z(o_data_bus[736]) );
  BUFFD6BWP30P140LVT U1556 ( .I(n3553), .Z(o_data_bus[735]) );
  BUFFD6BWP30P140LVT U1557 ( .I(n3554), .Z(o_data_bus[734]) );
  BUFFD6BWP30P140LVT U1558 ( .I(n3555), .Z(o_data_bus[733]) );
  BUFFD6BWP30P140LVT U1559 ( .I(n3556), .Z(o_data_bus[732]) );
  BUFFD6BWP30P140LVT U1560 ( .I(n3557), .Z(o_data_bus[731]) );
  BUFFD6BWP30P140LVT U1561 ( .I(n3558), .Z(o_data_bus[730]) );
  BUFFD6BWP30P140LVT U1562 ( .I(n3559), .Z(o_data_bus[729]) );
  BUFFD6BWP30P140LVT U1563 ( .I(n3560), .Z(o_data_bus[728]) );
  BUFFD6BWP30P140LVT U1564 ( .I(n3561), .Z(o_data_bus[727]) );
  BUFFD6BWP30P140LVT U1565 ( .I(n3562), .Z(o_data_bus[726]) );
  BUFFD6BWP30P140LVT U1566 ( .I(n3563), .Z(o_data_bus[725]) );
  BUFFD6BWP30P140LVT U1567 ( .I(n3564), .Z(o_data_bus[724]) );
  BUFFD6BWP30P140LVT U1568 ( .I(n3565), .Z(o_data_bus[723]) );
  BUFFD6BWP30P140LVT U1569 ( .I(n3566), .Z(o_data_bus[722]) );
  BUFFD6BWP30P140LVT U1570 ( .I(n3567), .Z(o_data_bus[721]) );
  BUFFD6BWP30P140LVT U1571 ( .I(n3568), .Z(o_data_bus[720]) );
  BUFFD6BWP30P140LVT U1572 ( .I(n3569), .Z(o_data_bus[719]) );
  BUFFD6BWP30P140LVT U1573 ( .I(n3570), .Z(o_data_bus[718]) );
  BUFFD6BWP30P140LVT U1574 ( .I(n3571), .Z(o_data_bus[717]) );
  BUFFD6BWP30P140LVT U1575 ( .I(n3572), .Z(o_data_bus[716]) );
  BUFFD6BWP30P140LVT U1576 ( .I(n3573), .Z(o_data_bus[715]) );
  BUFFD6BWP30P140LVT U1577 ( .I(n3574), .Z(o_data_bus[714]) );
  BUFFD6BWP30P140LVT U1578 ( .I(n3575), .Z(o_data_bus[713]) );
  BUFFD6BWP30P140LVT U1579 ( .I(n3576), .Z(o_data_bus[712]) );
  BUFFD6BWP30P140LVT U1580 ( .I(n3577), .Z(o_data_bus[711]) );
  BUFFD6BWP30P140LVT U1581 ( .I(n3578), .Z(o_data_bus[710]) );
  BUFFD6BWP30P140LVT U1582 ( .I(n3579), .Z(o_data_bus[709]) );
  BUFFD6BWP30P140LVT U1583 ( .I(n3580), .Z(o_data_bus[708]) );
  BUFFD6BWP30P140LVT U1584 ( .I(n3581), .Z(o_data_bus[707]) );
  BUFFD6BWP30P140LVT U1585 ( .I(n3582), .Z(o_data_bus[706]) );
  BUFFD6BWP30P140LVT U1586 ( .I(n3583), .Z(o_data_bus[705]) );
  BUFFD6BWP30P140LVT U1587 ( .I(n3584), .Z(o_data_bus[704]) );
  BUFFD6BWP30P140LVT U1588 ( .I(n3585), .Z(o_data_bus[703]) );
  BUFFD6BWP30P140LVT U1589 ( .I(n3586), .Z(o_data_bus[702]) );
  BUFFD6BWP30P140LVT U1590 ( .I(n3587), .Z(o_data_bus[701]) );
  BUFFD6BWP30P140LVT U1591 ( .I(n3588), .Z(o_data_bus[700]) );
  BUFFD6BWP30P140LVT U1592 ( .I(n3589), .Z(o_data_bus[699]) );
  BUFFD6BWP30P140LVT U1593 ( .I(n3590), .Z(o_data_bus[698]) );
  BUFFD6BWP30P140LVT U1594 ( .I(n3591), .Z(o_data_bus[697]) );
  BUFFD6BWP30P140LVT U1595 ( .I(n3592), .Z(o_data_bus[696]) );
  BUFFD6BWP30P140LVT U1596 ( .I(n3593), .Z(o_data_bus[695]) );
  BUFFD6BWP30P140LVT U1597 ( .I(n3594), .Z(o_data_bus[694]) );
  BUFFD6BWP30P140LVT U1598 ( .I(n3595), .Z(o_data_bus[693]) );
  BUFFD6BWP30P140LVT U1599 ( .I(n3596), .Z(o_data_bus[692]) );
  BUFFD6BWP30P140LVT U1600 ( .I(n3597), .Z(o_data_bus[691]) );
  BUFFD6BWP30P140LVT U1601 ( .I(n3598), .Z(o_data_bus[690]) );
  BUFFD6BWP30P140LVT U1602 ( .I(n3599), .Z(o_data_bus[689]) );
  BUFFD6BWP30P140LVT U1603 ( .I(n3600), .Z(o_data_bus[688]) );
  BUFFD6BWP30P140LVT U1604 ( .I(n3601), .Z(o_data_bus[687]) );
  BUFFD6BWP30P140LVT U1605 ( .I(n3602), .Z(o_data_bus[686]) );
  BUFFD6BWP30P140LVT U1606 ( .I(n3603), .Z(o_data_bus[685]) );
  BUFFD6BWP30P140LVT U1607 ( .I(n3604), .Z(o_data_bus[684]) );
  BUFFD6BWP30P140LVT U1608 ( .I(n3605), .Z(o_data_bus[683]) );
  BUFFD6BWP30P140LVT U1609 ( .I(n3081), .Z(o_data_bus[1207]) );
  BUFFD6BWP30P140LVT U1610 ( .I(n3606), .Z(o_data_bus[682]) );
  BUFFD6BWP30P140LVT U1611 ( .I(n3607), .Z(o_data_bus[681]) );
  BUFFD6BWP30P140LVT U1612 ( .I(n3608), .Z(o_data_bus[680]) );
  BUFFD6BWP30P140LVT U1613 ( .I(n3609), .Z(o_data_bus[679]) );
  BUFFD6BWP30P140LVT U1614 ( .I(n3610), .Z(o_data_bus[678]) );
  BUFFD6BWP30P140LVT U1615 ( .I(n3611), .Z(o_data_bus[677]) );
  BUFFD6BWP30P140LVT U1616 ( .I(n3612), .Z(o_data_bus[676]) );
  BUFFD6BWP30P140LVT U1617 ( .I(n3613), .Z(o_data_bus[675]) );
  BUFFD6BWP30P140LVT U1618 ( .I(n3614), .Z(o_data_bus[674]) );
  BUFFD6BWP30P140LVT U1619 ( .I(n3615), .Z(o_data_bus[673]) );
  BUFFD6BWP30P140LVT U1620 ( .I(n3616), .Z(o_data_bus[672]) );
  BUFFD6BWP30P140LVT U1621 ( .I(n3617), .Z(o_data_bus[671]) );
  BUFFD6BWP30P140LVT U1622 ( .I(n3618), .Z(o_data_bus[670]) );
  BUFFD6BWP30P140LVT U1623 ( .I(n3619), .Z(o_data_bus[669]) );
  BUFFD6BWP30P140LVT U1624 ( .I(n3620), .Z(o_data_bus[668]) );
  BUFFD6BWP30P140LVT U1625 ( .I(n3621), .Z(o_data_bus[667]) );
  BUFFD6BWP30P140LVT U1626 ( .I(n3622), .Z(o_data_bus[666]) );
  BUFFD6BWP30P140LVT U1627 ( .I(n3623), .Z(o_data_bus[665]) );
  BUFFD6BWP30P140LVT U1628 ( .I(n3624), .Z(o_data_bus[664]) );
  BUFFD6BWP30P140LVT U1629 ( .I(n3625), .Z(o_data_bus[663]) );
  BUFFD6BWP30P140LVT U1630 ( .I(n3626), .Z(o_data_bus[662]) );
  BUFFD6BWP30P140LVT U1631 ( .I(n3627), .Z(o_data_bus[661]) );
  BUFFD6BWP30P140LVT U1632 ( .I(n3628), .Z(o_data_bus[660]) );
  BUFFD6BWP30P140LVT U1633 ( .I(n3629), .Z(o_data_bus[659]) );
  BUFFD6BWP30P140LVT U1634 ( .I(n3630), .Z(o_data_bus[658]) );
  BUFFD6BWP30P140LVT U1635 ( .I(n3631), .Z(o_data_bus[657]) );
  BUFFD6BWP30P140LVT U1636 ( .I(n3632), .Z(o_data_bus[656]) );
  BUFFD6BWP30P140LVT U1637 ( .I(n3633), .Z(o_data_bus[655]) );
  BUFFD6BWP30P140LVT U1638 ( .I(n3634), .Z(o_data_bus[654]) );
  BUFFD6BWP30P140LVT U1639 ( .I(n3635), .Z(o_data_bus[653]) );
  BUFFD6BWP30P140LVT U1640 ( .I(n3636), .Z(o_data_bus[652]) );
  BUFFD6BWP30P140LVT U1641 ( .I(n3637), .Z(o_data_bus[651]) );
  BUFFD6BWP30P140LVT U1642 ( .I(n3638), .Z(o_data_bus[650]) );
  BUFFD6BWP30P140LVT U1643 ( .I(n3639), .Z(o_data_bus[649]) );
  BUFFD6BWP30P140LVT U1644 ( .I(n3640), .Z(o_data_bus[648]) );
  BUFFD6BWP30P140LVT U1645 ( .I(n3641), .Z(o_data_bus[647]) );
  BUFFD6BWP30P140LVT U1646 ( .I(n3642), .Z(o_data_bus[646]) );
  BUFFD6BWP30P140LVT U1647 ( .I(n3643), .Z(o_data_bus[645]) );
  BUFFD6BWP30P140LVT U1648 ( .I(n3644), .Z(o_data_bus[644]) );
  BUFFD6BWP30P140LVT U1649 ( .I(n3645), .Z(o_data_bus[643]) );
  BUFFD6BWP30P140LVT U1650 ( .I(n3646), .Z(o_data_bus[642]) );
  BUFFD6BWP30P140LVT U1651 ( .I(n3647), .Z(o_data_bus[641]) );
  BUFFD6BWP30P140LVT U1652 ( .I(n3648), .Z(o_data_bus[640]) );
  BUFFD6BWP30P140LVT U1653 ( .I(n3649), .Z(o_data_bus[639]) );
  BUFFD6BWP30P140LVT U1654 ( .I(n3650), .Z(o_data_bus[638]) );
  BUFFD6BWP30P140LVT U1655 ( .I(n3651), .Z(o_data_bus[637]) );
  BUFFD6BWP30P140LVT U1656 ( .I(n3652), .Z(o_data_bus[636]) );
  BUFFD6BWP30P140LVT U1657 ( .I(n3653), .Z(o_data_bus[635]) );
  BUFFD6BWP30P140LVT U1658 ( .I(n3654), .Z(o_data_bus[634]) );
  BUFFD6BWP30P140LVT U1659 ( .I(n3655), .Z(o_data_bus[633]) );
  BUFFD6BWP30P140LVT U1660 ( .I(n3656), .Z(o_data_bus[632]) );
  BUFFD6BWP30P140LVT U1661 ( .I(n3657), .Z(o_data_bus[631]) );
  BUFFD6BWP30P140LVT U1662 ( .I(n3658), .Z(o_data_bus[630]) );
  BUFFD6BWP30P140LVT U1663 ( .I(n3659), .Z(o_data_bus[629]) );
  BUFFD6BWP30P140LVT U1664 ( .I(n3660), .Z(o_data_bus[628]) );
  BUFFD6BWP30P140LVT U1665 ( .I(n3661), .Z(o_data_bus[627]) );
  BUFFD6BWP30P140LVT U1666 ( .I(n3662), .Z(o_data_bus[626]) );
  BUFFD6BWP30P140LVT U1667 ( .I(n3663), .Z(o_data_bus[625]) );
  BUFFD6BWP30P140LVT U1668 ( .I(n3664), .Z(o_data_bus[624]) );
  BUFFD6BWP30P140LVT U1669 ( .I(n3665), .Z(o_data_bus[623]) );
  BUFFD6BWP30P140LVT U1670 ( .I(n3666), .Z(o_data_bus[622]) );
  BUFFD6BWP30P140LVT U1671 ( .I(n3667), .Z(o_data_bus[621]) );
  BUFFD6BWP30P140LVT U1672 ( .I(n3668), .Z(o_data_bus[620]) );
  BUFFD6BWP30P140LVT U1673 ( .I(n3669), .Z(o_data_bus[619]) );
  BUFFD6BWP30P140LVT U1674 ( .I(n3670), .Z(o_data_bus[618]) );
  BUFFD6BWP30P140LVT U1675 ( .I(n3671), .Z(o_data_bus[617]) );
  BUFFD6BWP30P140LVT U1676 ( .I(n4352), .Z(o_cmd[0]) );
  BUFFD6BWP30P140LVT U1677 ( .I(n2676), .Z(o_data_bus[1612]) );
  BUFFD6BWP30P140LVT U1678 ( .I(n2675), .Z(o_data_bus[1613]) );
  BUFFD6BWP30P140LVT U1679 ( .I(n2674), .Z(o_data_bus[1614]) );
  BUFFD6BWP30P140LVT U1680 ( .I(n2673), .Z(o_data_bus[1615]) );
  BUFFD6BWP30P140LVT U1681 ( .I(n2672), .Z(o_data_bus[1616]) );
  BUFFD6BWP30P140LVT U1682 ( .I(n2671), .Z(o_data_bus[1617]) );
  BUFFD6BWP30P140LVT U1683 ( .I(n2670), .Z(o_data_bus[1618]) );
  BUFFD6BWP30P140LVT U1684 ( .I(n2669), .Z(o_data_bus[1619]) );
  BUFFD6BWP30P140LVT U1685 ( .I(n2668), .Z(o_data_bus[1620]) );
  BUFFD6BWP30P140LVT U1686 ( .I(n2667), .Z(o_data_bus[1621]) );
  BUFFD6BWP30P140LVT U1687 ( .I(n2666), .Z(o_data_bus[1622]) );
  BUFFD6BWP30P140LVT U1688 ( .I(n2665), .Z(o_data_bus[1623]) );
  BUFFD6BWP30P140LVT U1689 ( .I(n2664), .Z(o_data_bus[1624]) );
  BUFFD6BWP30P140LVT U1690 ( .I(n2663), .Z(o_data_bus[1625]) );
  BUFFD6BWP30P140LVT U1691 ( .I(n2662), .Z(o_data_bus[1626]) );
  BUFFD6BWP30P140LVT U1692 ( .I(n2661), .Z(o_data_bus[1627]) );
  BUFFD6BWP30P140LVT U1693 ( .I(n2660), .Z(o_data_bus[1628]) );
  BUFFD6BWP30P140LVT U1694 ( .I(n2659), .Z(o_data_bus[1629]) );
  BUFFD6BWP30P140LVT U1695 ( .I(n2658), .Z(o_data_bus[1630]) );
  BUFFD6BWP30P140LVT U1696 ( .I(n2657), .Z(o_data_bus[1631]) );
  BUFFD6BWP30P140LVT U1697 ( .I(n2656), .Z(o_data_bus[1632]) );
  BUFFD6BWP30P140LVT U1698 ( .I(n2655), .Z(o_data_bus[1633]) );
  BUFFD6BWP30P140LVT U1699 ( .I(n2654), .Z(o_data_bus[1634]) );
  BUFFD6BWP30P140LVT U1700 ( .I(n2653), .Z(o_data_bus[1635]) );
  BUFFD6BWP30P140LVT U1701 ( .I(n2652), .Z(o_data_bus[1636]) );
  BUFFD6BWP30P140LVT U1702 ( .I(n2651), .Z(o_data_bus[1637]) );
  BUFFD6BWP30P140LVT U1703 ( .I(n2650), .Z(o_data_bus[1638]) );
  BUFFD6BWP30P140LVT U1704 ( .I(n2649), .Z(o_data_bus[1639]) );
  BUFFD6BWP30P140LVT U1705 ( .I(n2648), .Z(o_data_bus[1640]) );
  BUFFD6BWP30P140LVT U1706 ( .I(n2647), .Z(o_data_bus[1641]) );
  BUFFD6BWP30P140LVT U1707 ( .I(n2646), .Z(o_data_bus[1642]) );
  BUFFD6BWP30P140LVT U1708 ( .I(n2645), .Z(o_data_bus[1643]) );
  BUFFD6BWP30P140LVT U1709 ( .I(n2644), .Z(o_data_bus[1644]) );
  BUFFD6BWP30P140LVT U1710 ( .I(n2643), .Z(o_data_bus[1645]) );
  BUFFD6BWP30P140LVT U1711 ( .I(n2642), .Z(o_data_bus[1646]) );
  BUFFD6BWP30P140LVT U1712 ( .I(n2641), .Z(o_data_bus[1647]) );
  BUFFD6BWP30P140LVT U1713 ( .I(n2640), .Z(o_data_bus[1648]) );
  BUFFD6BWP30P140LVT U1714 ( .I(n2639), .Z(o_data_bus[1649]) );
  BUFFD6BWP30P140LVT U1715 ( .I(n2638), .Z(o_data_bus[1650]) );
  BUFFD6BWP30P140LVT U1716 ( .I(n2637), .Z(o_data_bus[1651]) );
  BUFFD6BWP30P140LVT U1717 ( .I(n2636), .Z(o_data_bus[1652]) );
  BUFFD6BWP30P140LVT U1718 ( .I(n2635), .Z(o_data_bus[1653]) );
  BUFFD6BWP30P140LVT U1719 ( .I(n2634), .Z(o_data_bus[1654]) );
  BUFFD6BWP30P140LVT U1720 ( .I(n2633), .Z(o_data_bus[1655]) );
  BUFFD6BWP30P140LVT U1721 ( .I(n2632), .Z(o_data_bus[1656]) );
  BUFFD6BWP30P140LVT U1722 ( .I(n2631), .Z(o_data_bus[1657]) );
  BUFFD6BWP30P140LVT U1723 ( .I(n2630), .Z(o_data_bus[1658]) );
  BUFFD6BWP30P140LVT U1724 ( .I(n2629), .Z(o_data_bus[1659]) );
  BUFFD6BWP30P140LVT U1725 ( .I(n2628), .Z(o_data_bus[1660]) );
  BUFFD6BWP30P140LVT U1726 ( .I(n2627), .Z(o_data_bus[1661]) );
  BUFFD6BWP30P140LVT U1727 ( .I(n2626), .Z(o_data_bus[1662]) );
  BUFFD6BWP30P140LVT U1728 ( .I(n2625), .Z(o_data_bus[1663]) );
  BUFFD6BWP30P140LVT U1729 ( .I(n2624), .Z(o_data_bus[1664]) );
  BUFFD6BWP30P140LVT U1730 ( .I(n2623), .Z(o_data_bus[1665]) );
  BUFFD6BWP30P140LVT U1731 ( .I(n2622), .Z(o_data_bus[1666]) );
  BUFFD6BWP30P140LVT U1732 ( .I(n2621), .Z(o_data_bus[1667]) );
  BUFFD6BWP30P140LVT U1733 ( .I(n2620), .Z(o_data_bus[1668]) );
  BUFFD6BWP30P140LVT U1734 ( .I(n2619), .Z(o_data_bus[1669]) );
  BUFFD6BWP30P140LVT U1735 ( .I(n2618), .Z(o_data_bus[1670]) );
  BUFFD6BWP30P140LVT U1736 ( .I(n2617), .Z(o_data_bus[1671]) );
  BUFFD6BWP30P140LVT U1737 ( .I(n2616), .Z(o_data_bus[1672]) );
  BUFFD6BWP30P140LVT U1738 ( .I(n2615), .Z(o_data_bus[1673]) );
  BUFFD6BWP30P140LVT U1739 ( .I(n2614), .Z(o_data_bus[1674]) );
  BUFFD6BWP30P140LVT U1740 ( .I(n2613), .Z(o_data_bus[1675]) );
  BUFFD6BWP30P140LVT U1741 ( .I(n2612), .Z(o_data_bus[1676]) );
  BUFFD6BWP30P140LVT U1742 ( .I(n2611), .Z(o_data_bus[1677]) );
  BUFFD6BWP30P140LVT U1743 ( .I(n2610), .Z(o_data_bus[1678]) );
  BUFFD6BWP30P140LVT U1744 ( .I(n2609), .Z(o_data_bus[1679]) );
  BUFFD6BWP30P140LVT U1745 ( .I(n2608), .Z(o_data_bus[1680]) );
  BUFFD6BWP30P140LVT U1746 ( .I(n2607), .Z(o_data_bus[1681]) );
  BUFFD6BWP30P140LVT U1747 ( .I(n2606), .Z(o_data_bus[1682]) );
  BUFFD6BWP30P140LVT U1748 ( .I(n2605), .Z(o_data_bus[1683]) );
  BUFFD6BWP30P140LVT U1749 ( .I(n2604), .Z(o_data_bus[1684]) );
  BUFFD6BWP30P140LVT U1750 ( .I(n2603), .Z(o_data_bus[1685]) );
  BUFFD6BWP30P140LVT U1751 ( .I(n2602), .Z(o_data_bus[1686]) );
  BUFFD6BWP30P140LVT U1752 ( .I(n2601), .Z(o_data_bus[1687]) );
  BUFFD6BWP30P140LVT U1753 ( .I(n2600), .Z(o_data_bus[1688]) );
  BUFFD6BWP30P140LVT U1754 ( .I(n2599), .Z(o_data_bus[1689]) );
  BUFFD6BWP30P140LVT U1755 ( .I(n2598), .Z(o_data_bus[1690]) );
  BUFFD6BWP30P140LVT U1756 ( .I(n2597), .Z(o_data_bus[1691]) );
  BUFFD6BWP30P140LVT U1757 ( .I(n2596), .Z(o_data_bus[1692]) );
  BUFFD6BWP30P140LVT U1758 ( .I(n2595), .Z(o_data_bus[1693]) );
  BUFFD6BWP30P140LVT U1759 ( .I(n2594), .Z(o_data_bus[1694]) );
  BUFFD6BWP30P140LVT U1760 ( .I(n2593), .Z(o_data_bus[1695]) );
  BUFFD6BWP30P140LVT U1761 ( .I(n2592), .Z(o_data_bus[1696]) );
  BUFFD6BWP30P140LVT U1762 ( .I(n2591), .Z(o_data_bus[1697]) );
  BUFFD6BWP30P140LVT U1763 ( .I(n2590), .Z(o_data_bus[1698]) );
  BUFFD6BWP30P140LVT U1764 ( .I(n2589), .Z(o_data_bus[1699]) );
  BUFFD6BWP30P140LVT U1765 ( .I(n2588), .Z(o_data_bus[1700]) );
  BUFFD6BWP30P140LVT U1766 ( .I(n2587), .Z(o_data_bus[1701]) );
  BUFFD6BWP30P140LVT U1767 ( .I(n2586), .Z(o_data_bus[1702]) );
  BUFFD6BWP30P140LVT U1768 ( .I(n2585), .Z(o_data_bus[1703]) );
  BUFFD6BWP30P140LVT U1769 ( .I(n2584), .Z(o_data_bus[1704]) );
  BUFFD6BWP30P140LVT U1770 ( .I(n2583), .Z(o_data_bus[1705]) );
  BUFFD6BWP30P140LVT U1771 ( .I(n2582), .Z(o_data_bus[1706]) );
  BUFFD6BWP30P140LVT U1772 ( .I(n2581), .Z(o_data_bus[1707]) );
  BUFFD6BWP30P140LVT U1773 ( .I(n2580), .Z(o_data_bus[1708]) );
  BUFFD6BWP30P140LVT U1774 ( .I(n2579), .Z(o_data_bus[1709]) );
  BUFFD6BWP30P140LVT U1775 ( .I(n2578), .Z(o_data_bus[1710]) );
  BUFFD6BWP30P140LVT U1776 ( .I(n2577), .Z(o_data_bus[1711]) );
  BUFFD6BWP30P140LVT U1777 ( .I(n2576), .Z(o_data_bus[1712]) );
  BUFFD6BWP30P140LVT U1778 ( .I(n2575), .Z(o_data_bus[1713]) );
  BUFFD6BWP30P140LVT U1779 ( .I(n2574), .Z(o_data_bus[1714]) );
  BUFFD6BWP30P140LVT U1780 ( .I(n2573), .Z(o_data_bus[1715]) );
  BUFFD6BWP30P140LVT U1781 ( .I(n2572), .Z(o_data_bus[1716]) );
  BUFFD6BWP30P140LVT U1782 ( .I(n2571), .Z(o_data_bus[1717]) );
  BUFFD6BWP30P140LVT U1783 ( .I(n2570), .Z(o_data_bus[1718]) );
  BUFFD6BWP30P140LVT U1784 ( .I(n2569), .Z(o_data_bus[1719]) );
  BUFFD6BWP30P140LVT U1785 ( .I(n2568), .Z(o_data_bus[1720]) );
  BUFFD6BWP30P140LVT U1786 ( .I(n2567), .Z(o_data_bus[1721]) );
  BUFFD6BWP30P140LVT U1787 ( .I(n2566), .Z(o_data_bus[1722]) );
  BUFFD6BWP30P140LVT U1788 ( .I(n2565), .Z(o_data_bus[1723]) );
  BUFFD6BWP30P140LVT U1789 ( .I(n2564), .Z(o_data_bus[1724]) );
  BUFFD6BWP30P140LVT U1790 ( .I(n2563), .Z(o_data_bus[1725]) );
  BUFFD6BWP30P140LVT U1791 ( .I(n2562), .Z(o_data_bus[1726]) );
  BUFFD6BWP30P140LVT U1792 ( .I(n2561), .Z(o_data_bus[1727]) );
  BUFFD6BWP30P140LVT U1793 ( .I(n2560), .Z(o_data_bus[1728]) );
  BUFFD6BWP30P140LVT U1794 ( .I(n2559), .Z(o_data_bus[1729]) );
  BUFFD6BWP30P140LVT U1795 ( .I(n2558), .Z(o_data_bus[1730]) );
  BUFFD6BWP30P140LVT U1796 ( .I(n2557), .Z(o_data_bus[1731]) );
  BUFFD6BWP30P140LVT U1797 ( .I(n2556), .Z(o_data_bus[1732]) );
  BUFFD6BWP30P140LVT U1798 ( .I(n2555), .Z(o_data_bus[1733]) );
  BUFFD6BWP30P140LVT U1799 ( .I(n2554), .Z(o_data_bus[1734]) );
  BUFFD6BWP30P140LVT U1800 ( .I(n2553), .Z(o_data_bus[1735]) );
  BUFFD6BWP30P140LVT U1801 ( .I(n2552), .Z(o_data_bus[1736]) );
  BUFFD6BWP30P140LVT U1802 ( .I(n2551), .Z(o_data_bus[1737]) );
  BUFFD6BWP30P140LVT U1803 ( .I(n2550), .Z(o_data_bus[1738]) );
  BUFFD6BWP30P140LVT U1804 ( .I(n2549), .Z(o_data_bus[1739]) );
  BUFFD6BWP30P140LVT U1805 ( .I(n2548), .Z(o_data_bus[1740]) );
  BUFFD6BWP30P140LVT U1806 ( .I(n2547), .Z(o_data_bus[1741]) );
  BUFFD6BWP30P140LVT U1807 ( .I(n2546), .Z(o_data_bus[1742]) );
  BUFFD6BWP30P140LVT U1808 ( .I(n2545), .Z(o_data_bus[1743]) );
  BUFFD6BWP30P140LVT U1809 ( .I(n2544), .Z(o_data_bus[1744]) );
  BUFFD6BWP30P140LVT U1810 ( .I(n2543), .Z(o_data_bus[1745]) );
  BUFFD6BWP30P140LVT U1811 ( .I(n2542), .Z(o_data_bus[1746]) );
  BUFFD6BWP30P140LVT U1812 ( .I(n2541), .Z(o_data_bus[1747]) );
  BUFFD6BWP30P140LVT U1813 ( .I(n2540), .Z(o_data_bus[1748]) );
  BUFFD6BWP30P140LVT U1814 ( .I(n2539), .Z(o_data_bus[1749]) );
  BUFFD6BWP30P140LVT U1815 ( .I(n2538), .Z(o_data_bus[1750]) );
  BUFFD6BWP30P140LVT U1816 ( .I(n2537), .Z(o_data_bus[1751]) );
  BUFFD6BWP30P140LVT U1817 ( .I(n2536), .Z(o_data_bus[1752]) );
  BUFFD6BWP30P140LVT U1818 ( .I(n2535), .Z(o_data_bus[1753]) );
  BUFFD6BWP30P140LVT U1819 ( .I(n2534), .Z(o_data_bus[1754]) );
  BUFFD6BWP30P140LVT U1820 ( .I(n2533), .Z(o_data_bus[1755]) );
  BUFFD6BWP30P140LVT U1821 ( .I(n2532), .Z(o_data_bus[1756]) );
  BUFFD6BWP30P140LVT U1822 ( .I(n2531), .Z(o_data_bus[1757]) );
  BUFFD6BWP30P140LVT U1823 ( .I(n2530), .Z(o_data_bus[1758]) );
  BUFFD6BWP30P140LVT U1824 ( .I(n2529), .Z(o_data_bus[1759]) );
  BUFFD6BWP30P140LVT U1825 ( .I(n2528), .Z(o_data_bus[1760]) );
  BUFFD6BWP30P140LVT U1826 ( .I(n2527), .Z(o_data_bus[1761]) );
  BUFFD6BWP30P140LVT U1827 ( .I(n2526), .Z(o_data_bus[1762]) );
  BUFFD6BWP30P140LVT U1828 ( .I(n2525), .Z(o_data_bus[1763]) );
  BUFFD6BWP30P140LVT U1829 ( .I(n2524), .Z(o_data_bus[1764]) );
  BUFFD6BWP30P140LVT U1830 ( .I(n2523), .Z(o_data_bus[1765]) );
  BUFFD6BWP30P140LVT U1831 ( .I(n2522), .Z(o_data_bus[1766]) );
  BUFFD6BWP30P140LVT U1832 ( .I(n2521), .Z(o_data_bus[1767]) );
  BUFFD6BWP30P140LVT U1833 ( .I(n2520), .Z(o_data_bus[1768]) );
  BUFFD6BWP30P140LVT U1834 ( .I(n2519), .Z(o_data_bus[1769]) );
  BUFFD6BWP30P140LVT U1835 ( .I(n2518), .Z(o_data_bus[1770]) );
  BUFFD6BWP30P140LVT U1836 ( .I(n2517), .Z(o_data_bus[1771]) );
  BUFFD6BWP30P140LVT U1837 ( .I(n2516), .Z(o_data_bus[1772]) );
  BUFFD6BWP30P140LVT U1838 ( .I(n2515), .Z(o_data_bus[1773]) );
  BUFFD6BWP30P140LVT U1839 ( .I(n2514), .Z(o_data_bus[1774]) );
  BUFFD6BWP30P140LVT U1840 ( .I(n2513), .Z(o_data_bus[1775]) );
  BUFFD6BWP30P140LVT U1841 ( .I(n2512), .Z(o_data_bus[1776]) );
  BUFFD6BWP30P140LVT U1842 ( .I(n2511), .Z(o_data_bus[1777]) );
  BUFFD6BWP30P140LVT U1843 ( .I(n2510), .Z(o_data_bus[1778]) );
  BUFFD6BWP30P140LVT U1844 ( .I(n2509), .Z(o_data_bus[1779]) );
  BUFFD6BWP30P140LVT U1845 ( .I(n2508), .Z(o_data_bus[1780]) );
  BUFFD6BWP30P140LVT U1846 ( .I(n2507), .Z(o_data_bus[1781]) );
  BUFFD6BWP30P140LVT U1847 ( .I(n2506), .Z(o_data_bus[1782]) );
  BUFFD6BWP30P140LVT U1848 ( .I(n2505), .Z(o_data_bus[1783]) );
  BUFFD6BWP30P140LVT U1849 ( .I(n2504), .Z(o_data_bus[1784]) );
  BUFFD6BWP30P140LVT U1850 ( .I(n2503), .Z(o_data_bus[1785]) );
  BUFFD6BWP30P140LVT U1851 ( .I(n2502), .Z(o_data_bus[1786]) );
  BUFFD6BWP30P140LVT U1852 ( .I(n2501), .Z(o_data_bus[1787]) );
  BUFFD6BWP30P140LVT U1853 ( .I(n2500), .Z(o_data_bus[1788]) );
  BUFFD6BWP30P140LVT U1854 ( .I(n2499), .Z(o_data_bus[1789]) );
  BUFFD6BWP30P140LVT U1855 ( .I(n2498), .Z(o_data_bus[1790]) );
  BUFFD6BWP30P140LVT U1856 ( .I(n2497), .Z(o_data_bus[1791]) );
  BUFFD6BWP30P140LVT U1857 ( .I(n2496), .Z(o_data_bus[1792]) );
  BUFFD6BWP30P140LVT U1858 ( .I(n2495), .Z(o_data_bus[1793]) );
  BUFFD6BWP30P140LVT U1859 ( .I(n2494), .Z(o_data_bus[1794]) );
  BUFFD6BWP30P140LVT U1860 ( .I(n2493), .Z(o_data_bus[1795]) );
  BUFFD6BWP30P140LVT U1861 ( .I(n2492), .Z(o_data_bus[1796]) );
  BUFFD6BWP30P140LVT U1862 ( .I(n2491), .Z(o_data_bus[1797]) );
  BUFFD6BWP30P140LVT U1863 ( .I(n2490), .Z(o_data_bus[1798]) );
  BUFFD6BWP30P140LVT U1864 ( .I(n2489), .Z(o_data_bus[1799]) );
  BUFFD6BWP30P140LVT U1865 ( .I(n2488), .Z(o_data_bus[1800]) );
  BUFFD6BWP30P140LVT U1866 ( .I(n2487), .Z(o_data_bus[1801]) );
  BUFFD6BWP30P140LVT U1867 ( .I(n2486), .Z(o_data_bus[1802]) );
  BUFFD6BWP30P140LVT U1868 ( .I(n2485), .Z(o_data_bus[1803]) );
  BUFFD6BWP30P140LVT U1869 ( .I(n2484), .Z(o_data_bus[1804]) );
  BUFFD6BWP30P140LVT U1870 ( .I(n2483), .Z(o_data_bus[1805]) );
  BUFFD6BWP30P140LVT U1871 ( .I(n2482), .Z(o_data_bus[1806]) );
  BUFFD6BWP30P140LVT U1872 ( .I(n2481), .Z(o_data_bus[1807]) );
  BUFFD6BWP30P140LVT U1873 ( .I(n2480), .Z(o_data_bus[1808]) );
  BUFFD6BWP30P140LVT U1874 ( .I(n2479), .Z(o_data_bus[1809]) );
  BUFFD6BWP30P140LVT U1875 ( .I(n2478), .Z(o_data_bus[1810]) );
  BUFFD6BWP30P140LVT U1876 ( .I(n2477), .Z(o_data_bus[1811]) );
  BUFFD6BWP30P140LVT U1877 ( .I(n2476), .Z(o_data_bus[1812]) );
  BUFFD6BWP30P140LVT U1878 ( .I(n2475), .Z(o_data_bus[1813]) );
  BUFFD6BWP30P140LVT U1879 ( .I(n2474), .Z(o_data_bus[1814]) );
  BUFFD6BWP30P140LVT U1880 ( .I(n2473), .Z(o_data_bus[1815]) );
  BUFFD6BWP30P140LVT U1881 ( .I(n2472), .Z(o_data_bus[1816]) );
  BUFFD6BWP30P140LVT U1882 ( .I(n2471), .Z(o_data_bus[1817]) );
  BUFFD6BWP30P140LVT U1883 ( .I(n2470), .Z(o_data_bus[1818]) );
  BUFFD6BWP30P140LVT U1884 ( .I(n2469), .Z(o_data_bus[1819]) );
  BUFFD6BWP30P140LVT U1885 ( .I(n2468), .Z(o_data_bus[1820]) );
  BUFFD6BWP30P140LVT U1886 ( .I(n2467), .Z(o_data_bus[1821]) );
  BUFFD6BWP30P140LVT U1887 ( .I(n2466), .Z(o_data_bus[1822]) );
  BUFFD6BWP30P140LVT U1888 ( .I(n2465), .Z(o_data_bus[1823]) );
  BUFFD6BWP30P140LVT U1889 ( .I(n2464), .Z(o_data_bus[1824]) );
  BUFFD6BWP30P140LVT U1890 ( .I(n2463), .Z(o_data_bus[1825]) );
  BUFFD6BWP30P140LVT U1891 ( .I(n2462), .Z(o_data_bus[1826]) );
  BUFFD6BWP30P140LVT U1892 ( .I(n2461), .Z(o_data_bus[1827]) );
  BUFFD6BWP30P140LVT U1893 ( .I(n2460), .Z(o_data_bus[1828]) );
  BUFFD6BWP30P140LVT U1894 ( .I(n2459), .Z(o_data_bus[1829]) );
  BUFFD6BWP30P140LVT U1895 ( .I(n2458), .Z(o_data_bus[1830]) );
  BUFFD6BWP30P140LVT U1896 ( .I(n2457), .Z(o_data_bus[1831]) );
  BUFFD6BWP30P140LVT U1897 ( .I(n2456), .Z(o_data_bus[1832]) );
  BUFFD6BWP30P140LVT U1898 ( .I(n2455), .Z(o_data_bus[1833]) );
  BUFFD6BWP30P140LVT U1899 ( .I(n2454), .Z(o_data_bus[1834]) );
  BUFFD6BWP30P140LVT U1900 ( .I(n2453), .Z(o_data_bus[1835]) );
  BUFFD6BWP30P140LVT U1901 ( .I(n2452), .Z(o_data_bus[1836]) );
  BUFFD6BWP30P140LVT U1902 ( .I(n2451), .Z(o_data_bus[1837]) );
  BUFFD6BWP30P140LVT U1903 ( .I(n2450), .Z(o_data_bus[1838]) );
  BUFFD6BWP30P140LVT U1904 ( .I(n2449), .Z(o_data_bus[1839]) );
  BUFFD6BWP30P140LVT U1905 ( .I(n2448), .Z(o_data_bus[1840]) );
  BUFFD6BWP30P140LVT U1906 ( .I(n2447), .Z(o_data_bus[1841]) );
  BUFFD6BWP30P140LVT U1907 ( .I(n2446), .Z(o_data_bus[1842]) );
  BUFFD6BWP30P140LVT U1908 ( .I(n2445), .Z(o_data_bus[1843]) );
  BUFFD6BWP30P140LVT U1909 ( .I(n2444), .Z(o_data_bus[1844]) );
  BUFFD6BWP30P140LVT U1910 ( .I(n2443), .Z(o_data_bus[1845]) );
  BUFFD6BWP30P140LVT U1911 ( .I(n2442), .Z(o_data_bus[1846]) );
  BUFFD6BWP30P140LVT U1912 ( .I(n2441), .Z(o_data_bus[1847]) );
  BUFFD6BWP30P140LVT U1913 ( .I(n2440), .Z(o_data_bus[1848]) );
  BUFFD6BWP30P140LVT U1914 ( .I(n2439), .Z(o_data_bus[1849]) );
  BUFFD6BWP30P140LVT U1915 ( .I(n2438), .Z(o_data_bus[1850]) );
  BUFFD6BWP30P140LVT U1916 ( .I(n2437), .Z(o_data_bus[1851]) );
  BUFFD6BWP30P140LVT U1917 ( .I(n2436), .Z(o_data_bus[1852]) );
  BUFFD6BWP30P140LVT U1918 ( .I(n2435), .Z(o_data_bus[1853]) );
  BUFFD6BWP30P140LVT U1919 ( .I(n2434), .Z(o_data_bus[1854]) );
  BUFFD6BWP30P140LVT U1920 ( .I(n2433), .Z(o_data_bus[1855]) );
  BUFFD6BWP30P140LVT U1921 ( .I(n2432), .Z(o_data_bus[1856]) );
  BUFFD6BWP30P140LVT U1922 ( .I(n2431), .Z(o_data_bus[1857]) );
  BUFFD6BWP30P140LVT U1923 ( .I(n2430), .Z(o_data_bus[1858]) );
  BUFFD6BWP30P140LVT U1924 ( .I(n2429), .Z(o_data_bus[1859]) );
  BUFFD6BWP30P140LVT U1925 ( .I(n2428), .Z(o_data_bus[1860]) );
  BUFFD6BWP30P140LVT U1926 ( .I(n2427), .Z(o_data_bus[1861]) );
  BUFFD6BWP30P140LVT U1927 ( .I(n2426), .Z(o_data_bus[1862]) );
  BUFFD6BWP30P140LVT U1928 ( .I(n2425), .Z(o_data_bus[1863]) );
  BUFFD6BWP30P140LVT U1929 ( .I(n2424), .Z(o_data_bus[1864]) );
  BUFFD6BWP30P140LVT U1930 ( .I(n2423), .Z(o_data_bus[1865]) );
  BUFFD6BWP30P140LVT U1931 ( .I(n2422), .Z(o_data_bus[1866]) );
  BUFFD6BWP30P140LVT U1932 ( .I(n2421), .Z(o_data_bus[1867]) );
  BUFFD6BWP30P140LVT U1933 ( .I(n2420), .Z(o_data_bus[1868]) );
  BUFFD6BWP30P140LVT U1934 ( .I(n2419), .Z(o_data_bus[1869]) );
  BUFFD6BWP30P140LVT U1935 ( .I(n2418), .Z(o_data_bus[1870]) );
  BUFFD6BWP30P140LVT U1936 ( .I(n2417), .Z(o_data_bus[1871]) );
  BUFFD6BWP30P140LVT U1937 ( .I(n2416), .Z(o_data_bus[1872]) );
  BUFFD6BWP30P140LVT U1938 ( .I(n2415), .Z(o_data_bus[1873]) );
  BUFFD6BWP30P140LVT U1939 ( .I(n2414), .Z(o_data_bus[1874]) );
  BUFFD6BWP30P140LVT U1940 ( .I(n2413), .Z(o_data_bus[1875]) );
  BUFFD6BWP30P140LVT U1941 ( .I(n2412), .Z(o_data_bus[1876]) );
  BUFFD6BWP30P140LVT U1942 ( .I(n2411), .Z(o_data_bus[1877]) );
  BUFFD6BWP30P140LVT U1943 ( .I(n2410), .Z(o_data_bus[1878]) );
  BUFFD6BWP30P140LVT U1944 ( .I(n2409), .Z(o_data_bus[1879]) );
  BUFFD6BWP30P140LVT U1945 ( .I(n2408), .Z(o_data_bus[1880]) );
  BUFFD6BWP30P140LVT U1946 ( .I(n2407), .Z(o_data_bus[1881]) );
  BUFFD6BWP30P140LVT U1947 ( .I(n2406), .Z(o_data_bus[1882]) );
  BUFFD6BWP30P140LVT U1948 ( .I(n2405), .Z(o_data_bus[1883]) );
  BUFFD6BWP30P140LVT U1949 ( .I(n2404), .Z(o_data_bus[1884]) );
  BUFFD6BWP30P140LVT U1950 ( .I(n2403), .Z(o_data_bus[1885]) );
  BUFFD6BWP30P140LVT U1951 ( .I(n2402), .Z(o_data_bus[1886]) );
  BUFFD6BWP30P140LVT U1952 ( .I(n2401), .Z(o_data_bus[1887]) );
  BUFFD6BWP30P140LVT U1953 ( .I(n2400), .Z(o_data_bus[1888]) );
  BUFFD6BWP30P140LVT U1954 ( .I(n2399), .Z(o_data_bus[1889]) );
  BUFFD6BWP30P140LVT U1955 ( .I(n2398), .Z(o_data_bus[1890]) );
  BUFFD6BWP30P140LVT U1956 ( .I(n2397), .Z(o_data_bus[1891]) );
  BUFFD6BWP30P140LVT U1957 ( .I(n2396), .Z(o_data_bus[1892]) );
  BUFFD6BWP30P140LVT U1958 ( .I(n2395), .Z(o_data_bus[1893]) );
  BUFFD6BWP30P140LVT U1959 ( .I(n2394), .Z(o_data_bus[1894]) );
  BUFFD6BWP30P140LVT U1960 ( .I(n2393), .Z(o_data_bus[1895]) );
  BUFFD6BWP30P140LVT U1961 ( .I(n2392), .Z(o_data_bus[1896]) );
  BUFFD6BWP30P140LVT U1962 ( .I(n2391), .Z(o_data_bus[1897]) );
  BUFFD6BWP30P140LVT U1963 ( .I(n2390), .Z(o_data_bus[1898]) );
  BUFFD6BWP30P140LVT U1964 ( .I(n2389), .Z(o_data_bus[1899]) );
  BUFFD6BWP30P140LVT U1965 ( .I(n2388), .Z(o_data_bus[1900]) );
  BUFFD6BWP30P140LVT U1966 ( .I(n2387), .Z(o_data_bus[1901]) );
  BUFFD6BWP30P140LVT U1967 ( .I(n2386), .Z(o_data_bus[1902]) );
  BUFFD6BWP30P140LVT U1968 ( .I(n2385), .Z(o_data_bus[1903]) );
  BUFFD6BWP30P140LVT U1969 ( .I(n2384), .Z(o_data_bus[1904]) );
  BUFFD6BWP30P140LVT U1970 ( .I(n2383), .Z(o_data_bus[1905]) );
  BUFFD6BWP30P140LVT U1971 ( .I(n2382), .Z(o_data_bus[1906]) );
  BUFFD6BWP30P140LVT U1972 ( .I(n2381), .Z(o_data_bus[1907]) );
  BUFFD6BWP30P140LVT U1973 ( .I(n2380), .Z(o_data_bus[1908]) );
  BUFFD6BWP30P140LVT U1974 ( .I(n2379), .Z(o_data_bus[1909]) );
  BUFFD6BWP30P140LVT U1975 ( .I(n2378), .Z(o_data_bus[1910]) );
  BUFFD6BWP30P140LVT U1976 ( .I(n2377), .Z(o_data_bus[1911]) );
  BUFFD6BWP30P140LVT U1977 ( .I(n2376), .Z(o_data_bus[1912]) );
  BUFFD6BWP30P140LVT U1978 ( .I(n2375), .Z(o_data_bus[1913]) );
  BUFFD6BWP30P140LVT U1979 ( .I(n2374), .Z(o_data_bus[1914]) );
  BUFFD6BWP30P140LVT U1980 ( .I(n2373), .Z(o_data_bus[1915]) );
  BUFFD6BWP30P140LVT U1981 ( .I(n2372), .Z(o_data_bus[1916]) );
  BUFFD6BWP30P140LVT U1982 ( .I(n2371), .Z(o_data_bus[1917]) );
  BUFFD6BWP30P140LVT U1983 ( .I(n2370), .Z(o_data_bus[1918]) );
  BUFFD6BWP30P140LVT U1984 ( .I(n2369), .Z(o_data_bus[1919]) );
  BUFFD6BWP30P140LVT U1985 ( .I(n2368), .Z(o_data_bus[1920]) );
  BUFFD6BWP30P140LVT U1986 ( .I(n2367), .Z(o_data_bus[1921]) );
  BUFFD6BWP30P140LVT U1987 ( .I(n2366), .Z(o_data_bus[1922]) );
  BUFFD6BWP30P140LVT U1988 ( .I(n2365), .Z(o_data_bus[1923]) );
  BUFFD6BWP30P140LVT U1989 ( .I(n2364), .Z(o_data_bus[1924]) );
  BUFFD6BWP30P140LVT U1990 ( .I(n2363), .Z(o_data_bus[1925]) );
  BUFFD6BWP30P140LVT U1991 ( .I(n2362), .Z(o_data_bus[1926]) );
  BUFFD6BWP30P140LVT U1992 ( .I(n2361), .Z(o_data_bus[1927]) );
  BUFFD6BWP30P140LVT U1993 ( .I(n2360), .Z(o_data_bus[1928]) );
  BUFFD6BWP30P140LVT U1994 ( .I(n2359), .Z(o_data_bus[1929]) );
  BUFFD6BWP30P140LVT U1995 ( .I(n2358), .Z(o_data_bus[1930]) );
  BUFFD6BWP30P140LVT U1996 ( .I(n2357), .Z(o_data_bus[1931]) );
  BUFFD6BWP30P140LVT U1997 ( .I(n2356), .Z(o_data_bus[1932]) );
  BUFFD6BWP30P140LVT U1998 ( .I(n2355), .Z(o_data_bus[1933]) );
  BUFFD6BWP30P140LVT U1999 ( .I(n2354), .Z(o_data_bus[1934]) );
  BUFFD6BWP30P140LVT U2000 ( .I(n2353), .Z(o_data_bus[1935]) );
  BUFFD6BWP30P140LVT U2001 ( .I(n2352), .Z(o_data_bus[1936]) );
  BUFFD6BWP30P140LVT U2002 ( .I(n2351), .Z(o_data_bus[1937]) );
  BUFFD6BWP30P140LVT U2003 ( .I(n2350), .Z(o_data_bus[1938]) );
  BUFFD6BWP30P140LVT U2004 ( .I(n2349), .Z(o_data_bus[1939]) );
  BUFFD6BWP30P140LVT U2005 ( .I(n2348), .Z(o_data_bus[1940]) );
  BUFFD6BWP30P140LVT U2006 ( .I(n2347), .Z(o_data_bus[1941]) );
  BUFFD6BWP30P140LVT U2007 ( .I(n2346), .Z(o_data_bus[1942]) );
  BUFFD6BWP30P140LVT U2008 ( .I(n2345), .Z(o_data_bus[1943]) );
  BUFFD6BWP30P140LVT U2009 ( .I(n2344), .Z(o_data_bus[1944]) );
  BUFFD6BWP30P140LVT U2010 ( .I(n2343), .Z(o_data_bus[1945]) );
  BUFFD6BWP30P140LVT U2011 ( .I(n2342), .Z(o_data_bus[1946]) );
  BUFFD6BWP30P140LVT U2012 ( .I(n2341), .Z(o_data_bus[1947]) );
  BUFFD6BWP30P140LVT U2013 ( .I(n2340), .Z(o_data_bus[1948]) );
  BUFFD6BWP30P140LVT U2014 ( .I(n2339), .Z(o_data_bus[1949]) );
  BUFFD6BWP30P140LVT U2015 ( .I(n2338), .Z(o_data_bus[1950]) );
  BUFFD6BWP30P140LVT U2016 ( .I(n2337), .Z(o_data_bus[1951]) );
  BUFFD6BWP30P140LVT U2017 ( .I(n2336), .Z(o_data_bus[1952]) );
  BUFFD6BWP30P140LVT U2018 ( .I(n2335), .Z(o_data_bus[1953]) );
  BUFFD6BWP30P140LVT U2019 ( .I(n2334), .Z(o_data_bus[1954]) );
  BUFFD6BWP30P140LVT U2020 ( .I(n2333), .Z(o_data_bus[1955]) );
  BUFFD6BWP30P140LVT U2021 ( .I(n2332), .Z(o_data_bus[1956]) );
  BUFFD6BWP30P140LVT U2022 ( .I(n2331), .Z(o_data_bus[1957]) );
  BUFFD6BWP30P140LVT U2023 ( .I(n2330), .Z(o_data_bus[1958]) );
  BUFFD6BWP30P140LVT U2024 ( .I(n2329), .Z(o_data_bus[1959]) );
  BUFFD6BWP30P140LVT U2025 ( .I(n2328), .Z(o_data_bus[1960]) );
  BUFFD6BWP30P140LVT U2026 ( .I(n2327), .Z(o_data_bus[1961]) );
  BUFFD6BWP30P140LVT U2027 ( .I(n2326), .Z(o_data_bus[1962]) );
  BUFFD6BWP30P140LVT U2028 ( .I(n2325), .Z(o_data_bus[1963]) );
  BUFFD6BWP30P140LVT U2029 ( .I(n2324), .Z(o_data_bus[1964]) );
  BUFFD6BWP30P140LVT U2030 ( .I(n2323), .Z(o_data_bus[1965]) );
  BUFFD6BWP30P140LVT U2031 ( .I(n2322), .Z(o_data_bus[1966]) );
  BUFFD6BWP30P140LVT U2032 ( .I(n2321), .Z(o_data_bus[1967]) );
  BUFFD6BWP30P140LVT U2033 ( .I(n2320), .Z(o_data_bus[1968]) );
  BUFFD6BWP30P140LVT U2034 ( .I(n2319), .Z(o_data_bus[1969]) );
  BUFFD6BWP30P140LVT U2035 ( .I(n2318), .Z(o_data_bus[1970]) );
  BUFFD6BWP30P140LVT U2036 ( .I(n2317), .Z(o_data_bus[1971]) );
  BUFFD6BWP30P140LVT U2037 ( .I(n2316), .Z(o_data_bus[1972]) );
  BUFFD6BWP30P140LVT U2038 ( .I(n2315), .Z(o_data_bus[1973]) );
  BUFFD6BWP30P140LVT U2039 ( .I(n2314), .Z(o_data_bus[1974]) );
  BUFFD6BWP30P140LVT U2040 ( .I(n2313), .Z(o_data_bus[1975]) );
  BUFFD6BWP30P140LVT U2041 ( .I(n2312), .Z(o_data_bus[1976]) );
  BUFFD6BWP30P140LVT U2042 ( .I(n2311), .Z(o_data_bus[1977]) );
  BUFFD6BWP30P140LVT U2043 ( .I(n2310), .Z(o_data_bus[1978]) );
  BUFFD6BWP30P140LVT U2044 ( .I(n2309), .Z(o_data_bus[1979]) );
  BUFFD6BWP30P140LVT U2045 ( .I(n2308), .Z(o_data_bus[1980]) );
  BUFFD6BWP30P140LVT U2046 ( .I(n2307), .Z(o_data_bus[1981]) );
  BUFFD6BWP30P140LVT U2047 ( .I(n2306), .Z(o_data_bus[1982]) );
  BUFFD6BWP30P140LVT U2048 ( .I(n2305), .Z(o_data_bus[1983]) );
  BUFFD6BWP30P140LVT U2049 ( .I(n2304), .Z(o_data_bus[1984]) );
  BUFFD6BWP30P140LVT U2050 ( .I(n2303), .Z(o_data_bus[1985]) );
  BUFFD6BWP30P140LVT U2051 ( .I(n2302), .Z(o_data_bus[1986]) );
  BUFFD6BWP30P140LVT U2052 ( .I(n2301), .Z(o_data_bus[1987]) );
  BUFFD6BWP30P140LVT U2053 ( .I(n2300), .Z(o_data_bus[1988]) );
  BUFFD6BWP30P140LVT U2054 ( .I(n2299), .Z(o_data_bus[1989]) );
  BUFFD6BWP30P140LVT U2055 ( .I(n2298), .Z(o_data_bus[1990]) );
  BUFFD6BWP30P140LVT U2056 ( .I(n2297), .Z(o_data_bus[1991]) );
  BUFFD6BWP30P140LVT U2057 ( .I(n2296), .Z(o_data_bus[1992]) );
  BUFFD6BWP30P140LVT U2058 ( .I(n2295), .Z(o_data_bus[1993]) );
  BUFFD6BWP30P140LVT U2059 ( .I(n2294), .Z(o_data_bus[1994]) );
  BUFFD6BWP30P140LVT U2060 ( .I(n2293), .Z(o_data_bus[1995]) );
  BUFFD6BWP30P140LVT U2061 ( .I(n2292), .Z(o_data_bus[1996]) );
  BUFFD6BWP30P140LVT U2062 ( .I(n2291), .Z(o_data_bus[1997]) );
  BUFFD6BWP30P140LVT U2063 ( .I(n2290), .Z(o_data_bus[1998]) );
  BUFFD6BWP30P140LVT U2064 ( .I(n2289), .Z(o_data_bus[1999]) );
  BUFFD6BWP30P140LVT U2065 ( .I(n2288), .Z(o_data_bus[2000]) );
  BUFFD6BWP30P140LVT U2066 ( .I(n2287), .Z(o_data_bus[2001]) );
  BUFFD6BWP30P140LVT U2067 ( .I(n2286), .Z(o_data_bus[2002]) );
  BUFFD6BWP30P140LVT U2068 ( .I(n2285), .Z(o_data_bus[2003]) );
  BUFFD6BWP30P140LVT U2069 ( .I(n2284), .Z(o_data_bus[2004]) );
  BUFFD6BWP30P140LVT U2070 ( .I(n2283), .Z(o_data_bus[2005]) );
  BUFFD6BWP30P140LVT U2071 ( .I(n2282), .Z(o_data_bus[2006]) );
  BUFFD6BWP30P140LVT U2072 ( .I(n2281), .Z(o_data_bus[2007]) );
  BUFFD6BWP30P140LVT U2073 ( .I(n2280), .Z(o_data_bus[2008]) );
  BUFFD6BWP30P140LVT U2074 ( .I(n2279), .Z(o_data_bus[2009]) );
  BUFFD6BWP30P140LVT U2075 ( .I(n2278), .Z(o_data_bus[2010]) );
  BUFFD6BWP30P140LVT U2076 ( .I(n2277), .Z(o_data_bus[2011]) );
  BUFFD6BWP30P140LVT U2077 ( .I(n2276), .Z(o_data_bus[2012]) );
  BUFFD6BWP30P140LVT U2078 ( .I(n2275), .Z(o_data_bus[2013]) );
  BUFFD6BWP30P140LVT U2079 ( .I(n2274), .Z(o_data_bus[2014]) );
  BUFFD6BWP30P140LVT U2080 ( .I(n2273), .Z(o_data_bus[2015]) );
  BUFFD6BWP30P140LVT U2081 ( .I(n2272), .Z(o_data_bus[2016]) );
  BUFFD6BWP30P140LVT U2082 ( .I(n2271), .Z(o_data_bus[2017]) );
  BUFFD6BWP30P140LVT U2083 ( .I(n2270), .Z(o_data_bus[2018]) );
  BUFFD6BWP30P140LVT U2084 ( .I(n2269), .Z(o_data_bus[2019]) );
  BUFFD6BWP30P140LVT U2085 ( .I(n2268), .Z(o_data_bus[2020]) );
  BUFFD6BWP30P140LVT U2086 ( .I(n2267), .Z(o_data_bus[2021]) );
  BUFFD6BWP30P140LVT U2087 ( .I(n2266), .Z(o_data_bus[2022]) );
  BUFFD6BWP30P140LVT U2088 ( .I(n2265), .Z(o_data_bus[2023]) );
  BUFFD6BWP30P140LVT U2089 ( .I(n2264), .Z(o_data_bus[2024]) );
  BUFFD6BWP30P140LVT U2090 ( .I(n2263), .Z(o_data_bus[2025]) );
  BUFFD6BWP30P140LVT U2091 ( .I(n2262), .Z(o_data_bus[2026]) );
  BUFFD6BWP30P140LVT U2092 ( .I(n2261), .Z(o_data_bus[2027]) );
  BUFFD6BWP30P140LVT U2093 ( .I(n2260), .Z(o_data_bus[2028]) );
  BUFFD6BWP30P140LVT U2094 ( .I(n2259), .Z(o_data_bus[2029]) );
  BUFFD6BWP30P140LVT U2095 ( .I(n2258), .Z(o_data_bus[2030]) );
  BUFFD6BWP30P140LVT U2096 ( .I(n2257), .Z(o_data_bus[2031]) );
  BUFFD6BWP30P140LVT U2097 ( .I(n2256), .Z(o_data_bus[2032]) );
  BUFFD6BWP30P140LVT U2098 ( .I(n2255), .Z(o_data_bus[2033]) );
  BUFFD6BWP30P140LVT U2099 ( .I(n2254), .Z(o_data_bus[2034]) );
  BUFFD6BWP30P140LVT U2100 ( .I(n2253), .Z(o_data_bus[2035]) );
  BUFFD6BWP30P140LVT U2101 ( .I(n2252), .Z(o_data_bus[2036]) );
  BUFFD6BWP30P140LVT U2102 ( .I(n2251), .Z(o_data_bus[2037]) );
  BUFFD6BWP30P140LVT U2103 ( .I(n2250), .Z(o_data_bus[2038]) );
  BUFFD6BWP30P140LVT U2104 ( .I(n2249), .Z(o_data_bus[2039]) );
  BUFFD6BWP30P140LVT U2105 ( .I(n2248), .Z(o_data_bus[2040]) );
  BUFFD6BWP30P140LVT U2106 ( .I(n2247), .Z(o_data_bus[2041]) );
  BUFFD6BWP30P140LVT U2107 ( .I(n2246), .Z(o_data_bus[2042]) );
  BUFFD6BWP30P140LVT U2108 ( .I(n2245), .Z(o_data_bus[2043]) );
  BUFFD6BWP30P140LVT U2109 ( .I(n2244), .Z(o_data_bus[2044]) );
  BUFFD6BWP30P140LVT U2110 ( .I(n2243), .Z(o_data_bus[2045]) );
  BUFFD6BWP30P140LVT U2111 ( .I(n2242), .Z(o_data_bus[2046]) );
  BUFFD6BWP30P140LVT U2112 ( .I(n2241), .Z(o_data_bus[2047]) );
  BUFFD6BWP30P140LVT U2113 ( .I(n2240), .Z(o_valid[0]) );
  BUFFD6BWP30P140LVT U2114 ( .I(n2239), .Z(o_valid[1]) );
  BUFFD6BWP30P140LVT U2115 ( .I(n2238), .Z(o_valid[2]) );
  BUFFD6BWP30P140LVT U2116 ( .I(n2237), .Z(o_valid[3]) );
  BUFFD6BWP30P140LVT U2117 ( .I(n2236), .Z(o_valid[4]) );
  BUFFD6BWP30P140LVT U2118 ( .I(n2235), .Z(o_valid[5]) );
  BUFFD6BWP30P140LVT U2119 ( .I(n2234), .Z(o_valid[6]) );
  BUFFD6BWP30P140LVT U2120 ( .I(n2233), .Z(o_valid[7]) );
  BUFFD6BWP30P140LVT U2121 ( .I(n2232), .Z(o_valid[8]) );
  BUFFD6BWP30P140LVT U2122 ( .I(n2231), .Z(o_valid[9]) );
  BUFFD6BWP30P140LVT U2123 ( .I(n2230), .Z(o_valid[10]) );
  BUFFD6BWP30P140LVT U2124 ( .I(n2229), .Z(o_valid[11]) );
  BUFFD6BWP30P140LVT U2125 ( .I(n2228), .Z(o_valid[12]) );
  BUFFD6BWP30P140LVT U2126 ( .I(n2227), .Z(o_valid[13]) );
  BUFFD6BWP30P140LVT U2127 ( .I(n2226), .Z(o_valid[14]) );
  BUFFD6BWP30P140LVT U2128 ( .I(n2225), .Z(o_valid[15]) );
  BUFFD6BWP30P140LVT U2129 ( .I(n2224), .Z(o_valid[16]) );
  BUFFD6BWP30P140LVT U2130 ( .I(n2223), .Z(o_valid[17]) );
  BUFFD6BWP30P140LVT U2131 ( .I(n2222), .Z(o_valid[18]) );
  BUFFD6BWP30P140LVT U2132 ( .I(n2221), .Z(o_valid[19]) );
  BUFFD6BWP30P140LVT U2133 ( .I(n2220), .Z(o_valid[20]) );
  BUFFD6BWP30P140LVT U2134 ( .I(n2219), .Z(o_valid[21]) );
  BUFFD6BWP30P140LVT U2135 ( .I(n2218), .Z(o_valid[22]) );
  BUFFD6BWP30P140LVT U2136 ( .I(n2217), .Z(o_valid[23]) );
  BUFFD6BWP30P140LVT U2137 ( .I(n2216), .Z(o_valid[24]) );
  BUFFD6BWP30P140LVT U2138 ( .I(n2215), .Z(o_valid[25]) );
  BUFFD6BWP30P140LVT U2139 ( .I(n2214), .Z(o_valid[26]) );
  BUFFD6BWP30P140LVT U2140 ( .I(n2213), .Z(o_valid[27]) );
  BUFFD6BWP30P140LVT U2141 ( .I(n2212), .Z(o_valid[28]) );
  BUFFD6BWP30P140LVT U2142 ( .I(n2211), .Z(o_valid[29]) );
  BUFFD6BWP30P140LVT U2143 ( .I(n2210), .Z(o_valid[30]) );
  BUFFD6BWP30P140LVT U2144 ( .I(n2209), .Z(o_valid[31]) );
  BUFFD6BWP30P140LVT U2145 ( .I(n2208), .Z(o_valid[32]) );
  BUFFD6BWP30P140LVT U2146 ( .I(n2207), .Z(o_valid[33]) );
  BUFFD6BWP30P140LVT U2147 ( .I(n2206), .Z(o_valid[34]) );
  BUFFD6BWP30P140LVT U2148 ( .I(n2205), .Z(o_valid[35]) );
  BUFFD6BWP30P140LVT U2149 ( .I(n2204), .Z(o_valid[36]) );
  BUFFD6BWP30P140LVT U2150 ( .I(n2203), .Z(o_valid[37]) );
  BUFFD6BWP30P140LVT U2151 ( .I(n2202), .Z(o_valid[38]) );
  BUFFD6BWP30P140LVT U2152 ( .I(n2201), .Z(o_valid[39]) );
  BUFFD6BWP30P140LVT U2153 ( .I(n2200), .Z(o_valid[40]) );
  BUFFD6BWP30P140LVT U2154 ( .I(n2199), .Z(o_valid[41]) );
  BUFFD6BWP30P140LVT U2155 ( .I(n2198), .Z(o_valid[42]) );
  BUFFD6BWP30P140LVT U2156 ( .I(n2197), .Z(o_valid[43]) );
  BUFFD6BWP30P140LVT U2157 ( .I(n2196), .Z(o_valid[44]) );
  BUFFD6BWP30P140LVT U2158 ( .I(n2195), .Z(o_valid[45]) );
  BUFFD6BWP30P140LVT U2159 ( .I(n2194), .Z(o_valid[46]) );
  BUFFD6BWP30P140LVT U2160 ( .I(n2193), .Z(o_valid[47]) );
  BUFFD6BWP30P140LVT U2161 ( .I(n2192), .Z(o_valid[48]) );
  BUFFD6BWP30P140LVT U2162 ( .I(n2191), .Z(o_valid[49]) );
  BUFFD6BWP30P140LVT U2163 ( .I(n2190), .Z(o_valid[50]) );
  BUFFD6BWP30P140LVT U2164 ( .I(n2189), .Z(o_valid[51]) );
  BUFFD6BWP30P140LVT U2165 ( .I(n2188), .Z(o_valid[52]) );
  BUFFD6BWP30P140LVT U2166 ( .I(n2187), .Z(o_valid[53]) );
  BUFFD6BWP30P140LVT U2167 ( .I(n2186), .Z(o_valid[54]) );
  BUFFD6BWP30P140LVT U2168 ( .I(n2185), .Z(o_valid[55]) );
  BUFFD6BWP30P140LVT U2169 ( .I(n2184), .Z(o_valid[56]) );
  BUFFD6BWP30P140LVT U2170 ( .I(n2183), .Z(o_valid[57]) );
  BUFFD6BWP30P140LVT U2171 ( .I(n2182), .Z(o_valid[58]) );
  BUFFD6BWP30P140LVT U2172 ( .I(n2181), .Z(o_valid[59]) );
  BUFFD6BWP30P140LVT U2173 ( .I(n2180), .Z(o_valid[60]) );
  BUFFD6BWP30P140LVT U2174 ( .I(n2179), .Z(o_valid[61]) );
  BUFFD6BWP30P140LVT U2175 ( .I(n2178), .Z(o_valid[62]) );
  BUFFD6BWP30P140LVT U2176 ( .I(n2177), .Z(o_valid[63]) );
endmodule

