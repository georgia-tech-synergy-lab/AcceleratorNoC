

    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        CLK, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input CLK, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;
  wire   [127:0] buf_in_last_level_0__i_data_o_buf;
  wire   [127:0] buf_in_last_level_1__i_data_o_buf;
  wire   [127:0] buf_in_last_level_2__i_data_o_buf;
  wire   [127:0] buf_in_last_level_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[0]), .Z(
        buf_in_last_level_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[0]), .Z(
        buf_in_last_level_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[0]), .Z(
        buf_in_last_level_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[0]), .Z(
        buf_in_last_level_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[1]), .Z(
        buf_in_last_level_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[1]), .Z(
        buf_in_last_level_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[1]), .Z(
        buf_in_last_level_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[1]), .Z(
        buf_in_last_level_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[2]), .Z(
        buf_in_last_level_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[2]), .Z(
        buf_in_last_level_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[2]), .Z(
        buf_in_last_level_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[2]), .Z(
        buf_in_last_level_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[3]), .Z(
        buf_in_last_level_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[3]), .Z(
        buf_in_last_level_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[3]), .Z(
        buf_in_last_level_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[3]), .Z(
        buf_in_last_level_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[4]), .Z(
        buf_in_last_level_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[4]), .Z(
        buf_in_last_level_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[4]), .Z(
        buf_in_last_level_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[4]), .Z(
        buf_in_last_level_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[5]), .Z(
        buf_in_last_level_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[5]), .Z(
        buf_in_last_level_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[5]), .Z(
        buf_in_last_level_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[5]), .Z(
        buf_in_last_level_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[6]), .Z(
        buf_in_last_level_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[6]), .Z(
        buf_in_last_level_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[6]), .Z(
        buf_in_last_level_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[6]), .Z(
        buf_in_last_level_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[7]), .Z(
        buf_in_last_level_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[7]), .Z(
        buf_in_last_level_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[7]), .Z(
        buf_in_last_level_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[7]), .Z(
        buf_in_last_level_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[8]), .Z(
        buf_in_last_level_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[8]), .Z(
        buf_in_last_level_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[8]), .Z(
        buf_in_last_level_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[8]), .Z(
        buf_in_last_level_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[9]), .Z(
        buf_in_last_level_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[9]), .Z(
        buf_in_last_level_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[9]), .Z(
        buf_in_last_level_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[9]), .Z(
        buf_in_last_level_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[10]), .Z(
        buf_in_last_level_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[10]), .Z(
        buf_in_last_level_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[10]), .Z(
        buf_in_last_level_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[10]), .Z(
        buf_in_last_level_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[11]), .Z(
        buf_in_last_level_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[11]), .Z(
        buf_in_last_level_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[11]), .Z(
        buf_in_last_level_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[11]), .Z(
        buf_in_last_level_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[12]), .Z(
        buf_in_last_level_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[12]), .Z(
        buf_in_last_level_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[12]), .Z(
        buf_in_last_level_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[12]), .Z(
        buf_in_last_level_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[13]), .Z(
        buf_in_last_level_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[13]), .Z(
        buf_in_last_level_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[13]), .Z(
        buf_in_last_level_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[13]), .Z(
        buf_in_last_level_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[14]), .Z(
        buf_in_last_level_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[14]), .Z(
        buf_in_last_level_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[14]), .Z(
        buf_in_last_level_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[14]), .Z(
        buf_in_last_level_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[15]), .Z(
        buf_in_last_level_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[15]), .Z(
        buf_in_last_level_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[15]), .Z(
        buf_in_last_level_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[15]), .Z(
        buf_in_last_level_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[16]), .Z(
        buf_in_last_level_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[16]), .Z(
        buf_in_last_level_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[16]), .Z(
        buf_in_last_level_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[16]), .Z(
        buf_in_last_level_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[17]), .Z(
        buf_in_last_level_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[17]), .Z(
        buf_in_last_level_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[17]), .Z(
        buf_in_last_level_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[17]), .Z(
        buf_in_last_level_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[18]), .Z(
        buf_in_last_level_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[18]), .Z(
        buf_in_last_level_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[18]), .Z(
        buf_in_last_level_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[18]), .Z(
        buf_in_last_level_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[19]), .Z(
        buf_in_last_level_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[19]), .Z(
        buf_in_last_level_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[19]), .Z(
        buf_in_last_level_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[19]), .Z(
        buf_in_last_level_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[20]), .Z(
        buf_in_last_level_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[20]), .Z(
        buf_in_last_level_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[20]), .Z(
        buf_in_last_level_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[20]), .Z(
        buf_in_last_level_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[21]), .Z(
        buf_in_last_level_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[21]), .Z(
        buf_in_last_level_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[21]), .Z(
        buf_in_last_level_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[21]), .Z(
        buf_in_last_level_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[22]), .Z(
        buf_in_last_level_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[22]), .Z(
        buf_in_last_level_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[22]), .Z(
        buf_in_last_level_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[22]), .Z(
        buf_in_last_level_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[23]), .Z(
        buf_in_last_level_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[23]), .Z(
        buf_in_last_level_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[23]), .Z(
        buf_in_last_level_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[23]), .Z(
        buf_in_last_level_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[24]), .Z(
        buf_in_last_level_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[24]), .Z(
        buf_in_last_level_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[24]), .Z(
        buf_in_last_level_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[24]), .Z(
        buf_in_last_level_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[25]), .Z(
        buf_in_last_level_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[25]), .Z(
        buf_in_last_level_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[25]), .Z(
        buf_in_last_level_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[25]), .Z(
        buf_in_last_level_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[26]), .Z(
        buf_in_last_level_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[26]), .Z(
        buf_in_last_level_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[26]), .Z(
        buf_in_last_level_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[26]), .Z(
        buf_in_last_level_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[27]), .Z(
        buf_in_last_level_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[27]), .Z(
        buf_in_last_level_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[27]), .Z(
        buf_in_last_level_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[27]), .Z(
        buf_in_last_level_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[28]), .Z(
        buf_in_last_level_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[28]), .Z(
        buf_in_last_level_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[28]), .Z(
        buf_in_last_level_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[28]), .Z(
        buf_in_last_level_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[29]), .Z(
        buf_in_last_level_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[29]), .Z(
        buf_in_last_level_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[29]), .Z(
        buf_in_last_level_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[29]), .Z(
        buf_in_last_level_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[30]), .Z(
        buf_in_last_level_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[30]), .Z(
        buf_in_last_level_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[30]), .Z(
        buf_in_last_level_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[30]), .Z(
        buf_in_last_level_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[31]), .Z(
        buf_in_last_level_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[31]), .Z(
        buf_in_last_level_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[31]), .Z(
        buf_in_last_level_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[31]), .Z(
        buf_in_last_level_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[32]), .Z(
        buf_in_last_level_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[32]), .Z(
        buf_in_last_level_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[32]), .Z(
        buf_in_last_level_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[32]), .Z(
        buf_in_last_level_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[33]), .Z(
        buf_in_last_level_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[33]), .Z(
        buf_in_last_level_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[33]), .Z(
        buf_in_last_level_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[33]), .Z(
        buf_in_last_level_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[34]), .Z(
        buf_in_last_level_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[34]), .Z(
        buf_in_last_level_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[34]), .Z(
        buf_in_last_level_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[34]), .Z(
        buf_in_last_level_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[35]), .Z(
        buf_in_last_level_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[35]), .Z(
        buf_in_last_level_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[35]), .Z(
        buf_in_last_level_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[35]), .Z(
        buf_in_last_level_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[36]), .Z(
        buf_in_last_level_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[36]), .Z(
        buf_in_last_level_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[36]), .Z(
        buf_in_last_level_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[36]), .Z(
        buf_in_last_level_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[37]), .Z(
        buf_in_last_level_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[37]), .Z(
        buf_in_last_level_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[37]), .Z(
        buf_in_last_level_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[37]), .Z(
        buf_in_last_level_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[38]), .Z(
        buf_in_last_level_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[38]), .Z(
        buf_in_last_level_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[38]), .Z(
        buf_in_last_level_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[38]), .Z(
        buf_in_last_level_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[39]), .Z(
        buf_in_last_level_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[39]), .Z(
        buf_in_last_level_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[39]), .Z(
        buf_in_last_level_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[39]), .Z(
        buf_in_last_level_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[40]), .Z(
        buf_in_last_level_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[40]), .Z(
        buf_in_last_level_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[40]), .Z(
        buf_in_last_level_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[40]), .Z(
        buf_in_last_level_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[41]), .Z(
        buf_in_last_level_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[41]), .Z(
        buf_in_last_level_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[41]), .Z(
        buf_in_last_level_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[41]), .Z(
        buf_in_last_level_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[42]), .Z(
        buf_in_last_level_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[42]), .Z(
        buf_in_last_level_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[42]), .Z(
        buf_in_last_level_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[42]), .Z(
        buf_in_last_level_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[43]), .Z(
        buf_in_last_level_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[43]), .Z(
        buf_in_last_level_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[43]), .Z(
        buf_in_last_level_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[43]), .Z(
        buf_in_last_level_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[44]), .Z(
        buf_in_last_level_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[44]), .Z(
        buf_in_last_level_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[44]), .Z(
        buf_in_last_level_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[44]), .Z(
        buf_in_last_level_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[45]), .Z(
        buf_in_last_level_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[45]), .Z(
        buf_in_last_level_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[45]), .Z(
        buf_in_last_level_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[45]), .Z(
        buf_in_last_level_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[46]), .Z(
        buf_in_last_level_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[46]), .Z(
        buf_in_last_level_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[46]), .Z(
        buf_in_last_level_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[46]), .Z(
        buf_in_last_level_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[47]), .Z(
        buf_in_last_level_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[47]), .Z(
        buf_in_last_level_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[47]), .Z(
        buf_in_last_level_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[47]), .Z(
        buf_in_last_level_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[48]), .Z(
        buf_in_last_level_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[48]), .Z(
        buf_in_last_level_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[48]), .Z(
        buf_in_last_level_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[48]), .Z(
        buf_in_last_level_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[49]), .Z(
        buf_in_last_level_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[49]), .Z(
        buf_in_last_level_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[49]), .Z(
        buf_in_last_level_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[49]), .Z(
        buf_in_last_level_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[50]), .Z(
        buf_in_last_level_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[50]), .Z(
        buf_in_last_level_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[50]), .Z(
        buf_in_last_level_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[50]), .Z(
        buf_in_last_level_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[51]), .Z(
        buf_in_last_level_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[51]), .Z(
        buf_in_last_level_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[51]), .Z(
        buf_in_last_level_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[51]), .Z(
        buf_in_last_level_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[52]), .Z(
        buf_in_last_level_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[52]), .Z(
        buf_in_last_level_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[52]), .Z(
        buf_in_last_level_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[52]), .Z(
        buf_in_last_level_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[53]), .Z(
        buf_in_last_level_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[53]), .Z(
        buf_in_last_level_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[53]), .Z(
        buf_in_last_level_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[53]), .Z(
        buf_in_last_level_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[54]), .Z(
        buf_in_last_level_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[54]), .Z(
        buf_in_last_level_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[54]), .Z(
        buf_in_last_level_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[54]), .Z(
        buf_in_last_level_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[55]), .Z(
        buf_in_last_level_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[55]), .Z(
        buf_in_last_level_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[55]), .Z(
        buf_in_last_level_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[55]), .Z(
        buf_in_last_level_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[56]), .Z(
        buf_in_last_level_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[56]), .Z(
        buf_in_last_level_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[56]), .Z(
        buf_in_last_level_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[56]), .Z(
        buf_in_last_level_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[57]), .Z(
        buf_in_last_level_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[57]), .Z(
        buf_in_last_level_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[57]), .Z(
        buf_in_last_level_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[57]), .Z(
        buf_in_last_level_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[58]), .Z(
        buf_in_last_level_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[58]), .Z(
        buf_in_last_level_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[58]), .Z(
        buf_in_last_level_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[58]), .Z(
        buf_in_last_level_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[59]), .Z(
        buf_in_last_level_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[59]), .Z(
        buf_in_last_level_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[59]), .Z(
        buf_in_last_level_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[59]), .Z(
        buf_in_last_level_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[60]), .Z(
        buf_in_last_level_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[60]), .Z(
        buf_in_last_level_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[60]), .Z(
        buf_in_last_level_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[60]), .Z(
        buf_in_last_level_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[61]), .Z(
        buf_in_last_level_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[61]), .Z(
        buf_in_last_level_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[61]), .Z(
        buf_in_last_level_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[61]), .Z(
        buf_in_last_level_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[62]), .Z(
        buf_in_last_level_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[62]), .Z(
        buf_in_last_level_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[62]), .Z(
        buf_in_last_level_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[62]), .Z(
        buf_in_last_level_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[63]), .Z(
        buf_in_last_level_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[63]), .Z(
        buf_in_last_level_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[63]), .Z(
        buf_in_last_level_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[63]), .Z(
        buf_in_last_level_3__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[64]), .Z(
        buf_in_last_level_0__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[64]), .Z(
        buf_in_last_level_1__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[64]), .Z(
        buf_in_last_level_2__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[64]), .Z(
        buf_in_last_level_3__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[65]), .Z(
        buf_in_last_level_0__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[65]), .Z(
        buf_in_last_level_1__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[65]), .Z(
        buf_in_last_level_2__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[65]), .Z(
        buf_in_last_level_3__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[66]), .Z(
        buf_in_last_level_0__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[66]), .Z(
        buf_in_last_level_1__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[66]), .Z(
        buf_in_last_level_2__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[66]), .Z(
        buf_in_last_level_3__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[67]), .Z(
        buf_in_last_level_0__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[67]), .Z(
        buf_in_last_level_1__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[67]), .Z(
        buf_in_last_level_2__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[67]), .Z(
        buf_in_last_level_3__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[68]), .Z(
        buf_in_last_level_0__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[68]), .Z(
        buf_in_last_level_1__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[68]), .Z(
        buf_in_last_level_2__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[68]), .Z(
        buf_in_last_level_3__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[69]), .Z(
        buf_in_last_level_0__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[69]), .Z(
        buf_in_last_level_1__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[69]), .Z(
        buf_in_last_level_2__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[69]), .Z(
        buf_in_last_level_3__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[70]), .Z(
        buf_in_last_level_0__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[70]), .Z(
        buf_in_last_level_1__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[70]), .Z(
        buf_in_last_level_2__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[70]), .Z(
        buf_in_last_level_3__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[71]), .Z(
        buf_in_last_level_0__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[71]), .Z(
        buf_in_last_level_1__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[71]), .Z(
        buf_in_last_level_2__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[71]), .Z(
        buf_in_last_level_3__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[72]), .Z(
        buf_in_last_level_0__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[72]), .Z(
        buf_in_last_level_1__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[72]), .Z(
        buf_in_last_level_2__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[72]), .Z(
        buf_in_last_level_3__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[73]), .Z(
        buf_in_last_level_0__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[73]), .Z(
        buf_in_last_level_1__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[73]), .Z(
        buf_in_last_level_2__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[73]), .Z(
        buf_in_last_level_3__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[74]), .Z(
        buf_in_last_level_0__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[74]), .Z(
        buf_in_last_level_1__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[74]), .Z(
        buf_in_last_level_2__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[74]), .Z(
        buf_in_last_level_3__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[75]), .Z(
        buf_in_last_level_0__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[75]), .Z(
        buf_in_last_level_1__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[75]), .Z(
        buf_in_last_level_2__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[75]), .Z(
        buf_in_last_level_3__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[76]), .Z(
        buf_in_last_level_0__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[76]), .Z(
        buf_in_last_level_1__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[76]), .Z(
        buf_in_last_level_2__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[76]), .Z(
        buf_in_last_level_3__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[77]), .Z(
        buf_in_last_level_0__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[77]), .Z(
        buf_in_last_level_1__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[77]), .Z(
        buf_in_last_level_2__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[77]), .Z(
        buf_in_last_level_3__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[78]), .Z(
        buf_in_last_level_0__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[78]), .Z(
        buf_in_last_level_1__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[78]), .Z(
        buf_in_last_level_2__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[78]), .Z(
        buf_in_last_level_3__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[79]), .Z(
        buf_in_last_level_0__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[79]), .Z(
        buf_in_last_level_1__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[79]), .Z(
        buf_in_last_level_2__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[79]), .Z(
        buf_in_last_level_3__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[80]), .Z(
        buf_in_last_level_0__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[80]), .Z(
        buf_in_last_level_1__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[80]), .Z(
        buf_in_last_level_2__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[80]), .Z(
        buf_in_last_level_3__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[81]), .Z(
        buf_in_last_level_0__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[81]), .Z(
        buf_in_last_level_1__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[81]), .Z(
        buf_in_last_level_2__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[81]), .Z(
        buf_in_last_level_3__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[82]), .Z(
        buf_in_last_level_0__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[82]), .Z(
        buf_in_last_level_1__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[82]), .Z(
        buf_in_last_level_2__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[82]), .Z(
        buf_in_last_level_3__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[83]), .Z(
        buf_in_last_level_0__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[83]), .Z(
        buf_in_last_level_1__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[83]), .Z(
        buf_in_last_level_2__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[83]), .Z(
        buf_in_last_level_3__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[84]), .Z(
        buf_in_last_level_0__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[84]), .Z(
        buf_in_last_level_1__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[84]), .Z(
        buf_in_last_level_2__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[84]), .Z(
        buf_in_last_level_3__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[85]), .Z(
        buf_in_last_level_0__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[85]), .Z(
        buf_in_last_level_1__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[85]), .Z(
        buf_in_last_level_2__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[85]), .Z(
        buf_in_last_level_3__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[86]), .Z(
        buf_in_last_level_0__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[86]), .Z(
        buf_in_last_level_1__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[86]), .Z(
        buf_in_last_level_2__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[86]), .Z(
        buf_in_last_level_3__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[87]), .Z(
        buf_in_last_level_0__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[87]), .Z(
        buf_in_last_level_1__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[87]), .Z(
        buf_in_last_level_2__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[87]), .Z(
        buf_in_last_level_3__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[88]), .Z(
        buf_in_last_level_0__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[88]), .Z(
        buf_in_last_level_1__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[88]), .Z(
        buf_in_last_level_2__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[88]), .Z(
        buf_in_last_level_3__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[89]), .Z(
        buf_in_last_level_0__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[89]), .Z(
        buf_in_last_level_1__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[89]), .Z(
        buf_in_last_level_2__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[89]), .Z(
        buf_in_last_level_3__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[90]), .Z(
        buf_in_last_level_0__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[90]), .Z(
        buf_in_last_level_1__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[90]), .Z(
        buf_in_last_level_2__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[90]), .Z(
        buf_in_last_level_3__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[91]), .Z(
        buf_in_last_level_0__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[91]), .Z(
        buf_in_last_level_1__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[91]), .Z(
        buf_in_last_level_2__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[91]), .Z(
        buf_in_last_level_3__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[92]), .Z(
        buf_in_last_level_0__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[92]), .Z(
        buf_in_last_level_1__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[92]), .Z(
        buf_in_last_level_2__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[92]), .Z(
        buf_in_last_level_3__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[93]), .Z(
        buf_in_last_level_0__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[93]), .Z(
        buf_in_last_level_1__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[93]), .Z(
        buf_in_last_level_2__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[93]), .Z(
        buf_in_last_level_3__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[94]), .Z(
        buf_in_last_level_0__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[94]), .Z(
        buf_in_last_level_1__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[94]), .Z(
        buf_in_last_level_2__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[94]), .Z(
        buf_in_last_level_3__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[95]), .Z(
        buf_in_last_level_0__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[95]), .Z(
        buf_in_last_level_1__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[95]), .Z(
        buf_in_last_level_2__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[95]), .Z(
        buf_in_last_level_3__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[96]), .Z(
        buf_in_last_level_0__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[96]), .Z(
        buf_in_last_level_1__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[96]), .Z(
        buf_in_last_level_2__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[96]), .Z(
        buf_in_last_level_3__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[97]), .Z(
        buf_in_last_level_0__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[97]), .Z(
        buf_in_last_level_1__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[97]), .Z(
        buf_in_last_level_2__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[97]), .Z(
        buf_in_last_level_3__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[98]), .Z(
        buf_in_last_level_0__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[98]), .Z(
        buf_in_last_level_1__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[98]), .Z(
        buf_in_last_level_2__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[98]), .Z(
        buf_in_last_level_3__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[99]), .Z(
        buf_in_last_level_0__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[99]), .Z(
        buf_in_last_level_1__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[99]), .Z(
        buf_in_last_level_2__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[99]), .Z(
        buf_in_last_level_3__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[100]), .Z(
        buf_in_last_level_0__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[100]), .Z(
        buf_in_last_level_1__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[100]), .Z(
        buf_in_last_level_2__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[100]), .Z(
        buf_in_last_level_3__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[101]), .Z(
        buf_in_last_level_0__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[101]), .Z(
        buf_in_last_level_1__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[101]), .Z(
        buf_in_last_level_2__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[101]), .Z(
        buf_in_last_level_3__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[102]), .Z(
        buf_in_last_level_0__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[102]), .Z(
        buf_in_last_level_1__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[102]), .Z(
        buf_in_last_level_2__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[102]), .Z(
        buf_in_last_level_3__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[103]), .Z(
        buf_in_last_level_0__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[103]), .Z(
        buf_in_last_level_1__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[103]), .Z(
        buf_in_last_level_2__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[103]), .Z(
        buf_in_last_level_3__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[104]), .Z(
        buf_in_last_level_0__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[104]), .Z(
        buf_in_last_level_1__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[104]), .Z(
        buf_in_last_level_2__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[104]), .Z(
        buf_in_last_level_3__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[105]), .Z(
        buf_in_last_level_0__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[105]), .Z(
        buf_in_last_level_1__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[105]), .Z(
        buf_in_last_level_2__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[105]), .Z(
        buf_in_last_level_3__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[106]), .Z(
        buf_in_last_level_0__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[106]), .Z(
        buf_in_last_level_1__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[106]), .Z(
        buf_in_last_level_2__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[106]), .Z(
        buf_in_last_level_3__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[107]), .Z(
        buf_in_last_level_0__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[107]), .Z(
        buf_in_last_level_1__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[107]), .Z(
        buf_in_last_level_2__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[107]), .Z(
        buf_in_last_level_3__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[108]), .Z(
        buf_in_last_level_0__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[108]), .Z(
        buf_in_last_level_1__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[108]), .Z(
        buf_in_last_level_2__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[108]), .Z(
        buf_in_last_level_3__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[109]), .Z(
        buf_in_last_level_0__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[109]), .Z(
        buf_in_last_level_1__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[109]), .Z(
        buf_in_last_level_2__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[109]), .Z(
        buf_in_last_level_3__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[110]), .Z(
        buf_in_last_level_0__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[110]), .Z(
        buf_in_last_level_1__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[110]), .Z(
        buf_in_last_level_2__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[110]), .Z(
        buf_in_last_level_3__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[111]), .Z(
        buf_in_last_level_0__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[111]), .Z(
        buf_in_last_level_1__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[111]), .Z(
        buf_in_last_level_2__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[111]), .Z(
        buf_in_last_level_3__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[112]), .Z(
        buf_in_last_level_0__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[112]), .Z(
        buf_in_last_level_1__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[112]), .Z(
        buf_in_last_level_2__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[112]), .Z(
        buf_in_last_level_3__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[113]), .Z(
        buf_in_last_level_0__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[113]), .Z(
        buf_in_last_level_1__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[113]), .Z(
        buf_in_last_level_2__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[113]), .Z(
        buf_in_last_level_3__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[114]), .Z(
        buf_in_last_level_0__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[114]), .Z(
        buf_in_last_level_1__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[114]), .Z(
        buf_in_last_level_2__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[114]), .Z(
        buf_in_last_level_3__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[115]), .Z(
        buf_in_last_level_0__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[115]), .Z(
        buf_in_last_level_1__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[115]), .Z(
        buf_in_last_level_2__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[115]), .Z(
        buf_in_last_level_3__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[116]), .Z(
        buf_in_last_level_0__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[116]), .Z(
        buf_in_last_level_1__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[116]), .Z(
        buf_in_last_level_2__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[116]), .Z(
        buf_in_last_level_3__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[117]), .Z(
        buf_in_last_level_0__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[117]), .Z(
        buf_in_last_level_1__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[117]), .Z(
        buf_in_last_level_2__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[117]), .Z(
        buf_in_last_level_3__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[118]), .Z(
        buf_in_last_level_0__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[118]), .Z(
        buf_in_last_level_1__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[118]), .Z(
        buf_in_last_level_2__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[118]), .Z(
        buf_in_last_level_3__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[119]), .Z(
        buf_in_last_level_0__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[119]), .Z(
        buf_in_last_level_1__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[119]), .Z(
        buf_in_last_level_2__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[119]), .Z(
        buf_in_last_level_3__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[120]), .Z(
        buf_in_last_level_0__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[120]), .Z(
        buf_in_last_level_1__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[120]), .Z(
        buf_in_last_level_2__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[120]), .Z(
        buf_in_last_level_3__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[121]), .Z(
        buf_in_last_level_0__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[121]), .Z(
        buf_in_last_level_1__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[121]), .Z(
        buf_in_last_level_2__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[121]), .Z(
        buf_in_last_level_3__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[122]), .Z(
        buf_in_last_level_0__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[122]), .Z(
        buf_in_last_level_1__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[122]), .Z(
        buf_in_last_level_2__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[122]), .Z(
        buf_in_last_level_3__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[123]), .Z(
        buf_in_last_level_0__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[123]), .Z(
        buf_in_last_level_1__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[123]), .Z(
        buf_in_last_level_2__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[123]), .Z(
        buf_in_last_level_3__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[124]), .Z(
        buf_in_last_level_0__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[124]), .Z(
        buf_in_last_level_1__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[124]), .Z(
        buf_in_last_level_2__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[124]), .Z(
        buf_in_last_level_3__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[125]), .Z(
        buf_in_last_level_0__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[125]), .Z(
        buf_in_last_level_1__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[125]), .Z(
        buf_in_last_level_2__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[125]), .Z(
        buf_in_last_level_3__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[126]), .Z(
        buf_in_last_level_0__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[126]), .Z(
        buf_in_last_level_1__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[126]), .Z(
        buf_in_last_level_2__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[126]), .Z(
        buf_in_last_level_3__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[127]), .Z(
        buf_in_last_level_0__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[127]), .Z(
        buf_in_last_level_1__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[127]), .Z(
        buf_in_last_level_2__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[127]), .Z(
        buf_in_last_level_3__i_data_o_buf[127]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(CLK), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(CLK), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(CLK), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(CLK), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(CLK), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(CLK), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(CLK), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(CLK), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[101]), .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[102]), .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[105]), .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[107]), .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[109]), .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[110]), .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[111]), .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[112]), .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[115]), .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[82]), .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[86]), .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[61]), .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[63]), .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[26]), .Z(N292) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[22]), .Z(N288) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[23]), .Z(N289) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[24]), .Z(N290) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[25]), .Z(N291) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[27]), .Z(N293) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[28]), .Z(N294) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[21]), .Z(N287) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[20]), .Z(N286) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[31]), .Z(N297) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[30]), .Z(N296) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[29]), .Z(N295) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[62]), .Z(N362) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[60]), .Z(N360) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[59]), .Z(N359) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[58]), .Z(N358) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[57]), .Z(N357) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[56]), .Z(N356) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[55]), .Z(N355) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[54]), .Z(N354) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[53]), .Z(N353) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[52]), .Z(N352) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[51]), .Z(N351) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[50]), .Z(N350) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[49]), .Z(N349) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[48]), .Z(N348) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[47]), .Z(N347) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[46]), .Z(N346) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[45]), .Z(N345) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[44]), .Z(N344) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[43]), .Z(N343) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[42]), .Z(N342) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[41]), .Z(N341) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[40]), .Z(N340) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[39]), .Z(N339) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[38]), .Z(N338) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[37]), .Z(N337) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[0]), .Z(N266) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[1]), .Z(N267) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[3]), .Z(N269) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[4]), .Z(N270) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[5]), .Z(N271) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[7]), .Z(N273) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[8]), .Z(N274) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[9]), .Z(N275) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[10]), .Z(N276) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[11]), .Z(N277) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[12]), .Z(N278) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[13]), .Z(N279) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[14]), .Z(N280) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[15]), .Z(N281) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[16]), .Z(N282) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[17]), .Z(N283) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[18]), .Z(N284) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[19]), .Z(N285) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[36]), .Z(N336) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[35]), .Z(N335) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[34]), .Z(N334) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[33]), .Z(N333) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[32]), .Z(N332) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[90]), .Z(N424) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[89]), .Z(N423) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[88]), .Z(N422) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[87]), .Z(N421) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[85]), .Z(N419) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[84]), .Z(N418) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[83]), .Z(N417) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[81]), .Z(N415) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[80]), .Z(N414) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[79]), .Z(N413) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[78]), .Z(N412) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[77]), .Z(N411) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[76]), .Z(N410) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[75]), .Z(N409) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[74]), .Z(N408) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[73]), .Z(N407) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[72]), .Z(N406) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[71]), .Z(N405) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[70]), .Z(N404) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[69]), .Z(N403) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[68]), .Z(N402) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[67]), .Z(N401) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[66]), .Z(N400) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[65]), .Z(N399) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[64]), .Z(N398) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[95]), .Z(N429) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[94]), .Z(N428) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[93]), .Z(N427) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[92]), .Z(N426) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[91]), .Z(N425) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_0 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD2BWP30P140LVT U3 ( .I(n147), .ZN(n3) );
  INVD2BWP30P140LVT U4 ( .I(n145), .ZN(n222) );
  NR3D0P7BWP30P140LVT U5 ( .A1(n40), .A2(n39), .A3(n38), .ZN(n41) );
  NR2D1BWP30P140LVT U6 ( .A1(i_cmd[5]), .A2(i_cmd[6]), .ZN(n8) );
  AN3D1BWP30P140LVT U7 ( .A1(n35), .A2(i_cmd[3]), .A3(i_valid[3]), .Z(n1) );
  CKAN2D4BWP30P140LVT U8 ( .A1(n11), .A2(n42), .Z(n2) );
  ND2D1BWP30P140LVT U9 ( .A1(i_data_bus[0]), .A2(n2), .ZN(n53) );
  ND2OPTIBD2BWP30P140LVT U10 ( .A1(n8), .A2(n7), .ZN(n40) );
  INVD2BWP30P140LVT U11 ( .I(n48), .ZN(n220) );
  ND2OPTIBD1BWP30P140LVT U12 ( .A1(n36), .A2(n33), .ZN(n48) );
  NR2D1BWP30P140LVT U13 ( .A1(n4), .A2(n32), .ZN(n33) );
  ND2D1BWP30P140LVT U14 ( .A1(i_valid[1]), .A2(i_cmd[1]), .ZN(n32) );
  NR2D1BWP30P140LVT U15 ( .A1(n4), .A2(i_cmd[1]), .ZN(n42) );
  INVD1BWP30P140LVT U16 ( .I(n34), .ZN(n35) );
  INVD1BWP30P140LVT U17 ( .I(n5), .ZN(n6) );
  ND2D1BWP30P140LVT U18 ( .A1(n27), .A2(n14), .ZN(n15) );
  MAOI22D1BWP30P140LVT U19 ( .A1(n157), .A2(i_data_bus[205]), .B1(n130), .B2(
        n129), .ZN(n131) );
  AOI21D1BWP30P140LVT U20 ( .A1(n2), .A2(i_data_bus[1]), .B(n26), .ZN(n45) );
  ND3D1BWP30P140LVT U21 ( .A1(n51), .A2(n50), .A3(n49), .ZN(N395) );
  AOI21D1BWP30P140LVT U22 ( .A1(n2), .A2(i_data_bus[26]), .B(n47), .ZN(n51) );
  AOI22D1BWP30P140LVT U23 ( .A1(n3), .A2(i_data_bus[122]), .B1(n162), .B2(
        i_data_bus[154]), .ZN(n49) );
  AOI21D1BWP30P140LVT U24 ( .A1(n2), .A2(i_data_bus[28]), .B(n159), .ZN(n165)
         );
  AOI21D1BWP30P140LVT U25 ( .A1(n2), .A2(i_data_bus[30]), .B(n152), .ZN(n155)
         );
  AOI21D1BWP30P140LVT U26 ( .A1(n2), .A2(i_data_bus[31]), .B(n143), .ZN(n150)
         );
  NR2D1BWP30P140LVT U27 ( .A1(n3), .A2(n162), .ZN(n60) );
  NR2D3BWP30P140LVT U28 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n27) );
  INR2D4BWP30P140LVT U29 ( .A1(n16), .B1(n22), .ZN(n17) );
  OR2D1BWP30P140LVT U30 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .Z(n4) );
  INR2D1BWP30P140LVT U31 ( .A1(i_en), .B1(rst), .ZN(n5) );
  NR2OPTPAD1BWP30P140LVT U32 ( .A1(i_cmd[7]), .A2(n6), .ZN(n7) );
  INR2D1BWP30P140LVT U33 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n9) );
  ND2D1BWP30P140LVT U34 ( .A1(n9), .A2(i_cmd[0]), .ZN(n10) );
  NR2D1BWP30P140LVT U35 ( .A1(n40), .A2(n10), .ZN(n11) );
  ND2OPTIBD1BWP30P140LVT U36 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n12) );
  NR3D0P7BWP30P140LVT U37 ( .A1(n12), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n16)
         );
  OR2D2BWP30P140LVT U38 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .Z(n34) );
  INR2D1BWP30P140LVT U39 ( .A1(i_en), .B1(rst), .ZN(n13) );
  INR2D1BWP30P140LVT U40 ( .A1(n13), .B1(i_cmd[3]), .ZN(n14) );
  OR2D4BWP30P140LVT U41 ( .A1(n34), .A2(n15), .Z(n22) );
  INVD1BWP30P140LVT U42 ( .I(i_cmd[6]), .ZN(n18) );
  INR4D1BWP30P140LVT U43 ( .A1(i_valid[6]), .B1(i_cmd[5]), .B2(i_cmd[7]), .B3(
        n18), .ZN(n19) );
  INR2D1BWP30P140LVT U44 ( .A1(n19), .B1(n22), .ZN(n20) );
  INVD2BWP30P140LVT U45 ( .I(n20), .ZN(n52) );
  INVD3BWP30P140LVT U46 ( .I(n52), .ZN(n157) );
  INVD1BWP30P140LVT U47 ( .I(i_cmd[5]), .ZN(n21) );
  INR4D1BWP30P140LVT U48 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n21), .ZN(n23) );
  INR2D2BWP30P140LVT U49 ( .A1(n23), .B1(n22), .ZN(n24) );
  INVD2BWP30P140LVT U50 ( .I(n24), .ZN(n130) );
  INVD3BWP30P140LVT U51 ( .I(n130), .ZN(n216) );
  AOI22D1BWP30P140LVT U52 ( .A1(n157), .A2(i_data_bus[193]), .B1(n216), .B2(
        i_data_bus[161]), .ZN(n25) );
  IOA21D1BWP30P140LVT U53 ( .A1(n17), .A2(i_data_bus[225]), .B(n25), .ZN(n26)
         );
  INR2D2BWP30P140LVT U54 ( .A1(n27), .B1(n40), .ZN(n36) );
  INVD1BWP30P140LVT U55 ( .I(i_cmd[1]), .ZN(n29) );
  INVD1BWP30P140LVT U56 ( .I(i_cmd[3]), .ZN(n28) );
  ND4D1BWP30P140LVT U57 ( .A1(n29), .A2(n28), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n30) );
  INR2D1BWP30P140LVT U58 ( .A1(n36), .B1(n30), .ZN(n31) );
  INVD2BWP30P140LVT U59 ( .I(n31), .ZN(n65) );
  INVD2BWP30P140LVT U60 ( .I(n65), .ZN(n221) );
  AOI22D1BWP30P140LVT U61 ( .A1(n221), .A2(i_data_bus[65]), .B1(n220), .B2(
        i_data_bus[33]), .ZN(n44) );
  CKND2D2BWP30P140LVT U62 ( .A1(n1), .A2(n36), .ZN(n147) );
  INVD2BWP30P140LVT U63 ( .I(n147), .ZN(n223) );
  INVD1BWP30P140LVT U64 ( .I(i_cmd[0]), .ZN(n37) );
  ND2D1BWP30P140LVT U65 ( .A1(n37), .A2(i_cmd[4]), .ZN(n39) );
  INVD1BWP30P140LVT U66 ( .I(i_valid[4]), .ZN(n38) );
  ND2OPTIBD2BWP30P140LVT U67 ( .A1(n42), .A2(n41), .ZN(n145) );
  AOI22D1BWP30P140LVT U68 ( .A1(n223), .A2(i_data_bus[97]), .B1(n222), .B2(
        i_data_bus[129]), .ZN(n43) );
  ND3D1BWP30P140LVT U69 ( .A1(n45), .A2(n44), .A3(n43), .ZN(N370) );
  INVD4BWP30P140LVT U70 ( .I(n130), .ZN(n156) );
  AOI22D1BWP30P140LVT U71 ( .A1(n157), .A2(i_data_bus[218]), .B1(n156), .B2(
        i_data_bus[186]), .ZN(n46) );
  IOA21D1BWP30P140LVT U72 ( .A1(n17), .A2(i_data_bus[250]), .B(n46), .ZN(n47)
         );
  INVD1BWP30P140LVT U73 ( .I(n65), .ZN(n161) );
  INVD2BWP30P140LVT U74 ( .I(n48), .ZN(n160) );
  AOI22D1BWP30P140LVT U75 ( .A1(n161), .A2(i_data_bus[90]), .B1(n160), .B2(
        i_data_bus[58]), .ZN(n50) );
  INVD3BWP30P140LVT U76 ( .I(n145), .ZN(n162) );
  INVD1BWP30P140LVT U77 ( .I(n17), .ZN(n56) );
  INVD1BWP30P140LVT U78 ( .I(i_data_bus[224]), .ZN(n55) );
  INVD3BWP30P140LVT U79 ( .I(n52), .ZN(n217) );
  AOI22D2BWP30P140LVT U80 ( .A1(n217), .A2(i_data_bus[192]), .B1(n216), .B2(
        i_data_bus[160]), .ZN(n54) );
  OA211D1BWP30P140LVT U81 ( .A1(n56), .A2(n55), .B(n54), .C(n53), .Z(n59) );
  AOI22D1BWP30P140LVT U82 ( .A1(n221), .A2(i_data_bus[64]), .B1(n220), .B2(
        i_data_bus[32]), .ZN(n58) );
  AOI22D1BWP30P140LVT U83 ( .A1(n223), .A2(i_data_bus[96]), .B1(n222), .B2(
        i_data_bus[128]), .ZN(n57) );
  ND3D1BWP30P140LVT U84 ( .A1(n59), .A2(n58), .A3(n57), .ZN(N369) );
  NR4D0BWP30P140LVT U85 ( .A1(n2), .A2(n17), .A3(n157), .A4(n156), .ZN(n62) );
  NR2D1BWP30P140LVT U86 ( .A1(n161), .A2(n160), .ZN(n61) );
  ND3D1BWP30P140LVT U87 ( .A1(n62), .A2(n61), .A3(n60), .ZN(N402) );
  AOI22D1BWP30P140LVT U88 ( .A1(n217), .A2(i_data_bus[214]), .B1(n156), .B2(
        i_data_bus[182]), .ZN(n63) );
  IOA21D1BWP30P140LVT U89 ( .A1(n17), .A2(i_data_bus[246]), .B(n63), .ZN(n64)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n2), .A2(i_data_bus[22]), .B(n64), .ZN(n68) );
  INVD2BWP30P140LVT U91 ( .I(n65), .ZN(n138) );
  AOI22D1BWP30P140LVT U92 ( .A1(n138), .A2(i_data_bus[86]), .B1(n160), .B2(
        i_data_bus[54]), .ZN(n67) );
  AOI22D1BWP30P140LVT U93 ( .A1(n3), .A2(i_data_bus[118]), .B1(n162), .B2(
        i_data_bus[150]), .ZN(n66) );
  ND3D1BWP30P140LVT U94 ( .A1(n68), .A2(n67), .A3(n66), .ZN(N391) );
  AOI22D1BWP30P140LVT U95 ( .A1(n217), .A2(i_data_bus[219]), .B1(n156), .B2(
        i_data_bus[187]), .ZN(n69) );
  IOA21D1BWP30P140LVT U96 ( .A1(n17), .A2(i_data_bus[251]), .B(n69), .ZN(n70)
         );
  AOI21D1BWP30P140LVT U97 ( .A1(n2), .A2(i_data_bus[27]), .B(n70), .ZN(n73) );
  AOI22D1BWP30P140LVT U98 ( .A1(n161), .A2(i_data_bus[91]), .B1(n160), .B2(
        i_data_bus[59]), .ZN(n72) );
  AOI22D1BWP30P140LVT U99 ( .A1(n3), .A2(i_data_bus[123]), .B1(n162), .B2(
        i_data_bus[155]), .ZN(n71) );
  ND3D1BWP30P140LVT U100 ( .A1(n73), .A2(n72), .A3(n71), .ZN(N396) );
  AOI22D1BWP30P140LVT U101 ( .A1(n157), .A2(i_data_bus[221]), .B1(n156), .B2(
        i_data_bus[189]), .ZN(n74) );
  IOA21D1BWP30P140LVT U102 ( .A1(n17), .A2(i_data_bus[253]), .B(n74), .ZN(n75)
         );
  AOI21D1BWP30P140LVT U103 ( .A1(n2), .A2(i_data_bus[29]), .B(n75), .ZN(n78)
         );
  AOI22D1BWP30P140LVT U104 ( .A1(n161), .A2(i_data_bus[93]), .B1(n160), .B2(
        i_data_bus[61]), .ZN(n77) );
  AOI22D1BWP30P140LVT U105 ( .A1(n3), .A2(i_data_bus[125]), .B1(n162), .B2(
        i_data_bus[157]), .ZN(n76) );
  ND3D1BWP30P140LVT U106 ( .A1(n78), .A2(n77), .A3(n76), .ZN(N398) );
  AOI22D1BWP30P140LVT U107 ( .A1(n157), .A2(i_data_bus[215]), .B1(n156), .B2(
        i_data_bus[183]), .ZN(n79) );
  IOA21D1BWP30P140LVT U108 ( .A1(n17), .A2(i_data_bus[247]), .B(n79), .ZN(n80)
         );
  AOI21D1BWP30P140LVT U109 ( .A1(n2), .A2(i_data_bus[23]), .B(n80), .ZN(n83)
         );
  AOI22D1BWP30P140LVT U110 ( .A1(n138), .A2(i_data_bus[87]), .B1(n160), .B2(
        i_data_bus[55]), .ZN(n82) );
  AOI22D1BWP30P140LVT U111 ( .A1(n3), .A2(i_data_bus[119]), .B1(n162), .B2(
        i_data_bus[151]), .ZN(n81) );
  ND3D1BWP30P140LVT U112 ( .A1(n83), .A2(n82), .A3(n81), .ZN(N392) );
  AOI22D1BWP30P140LVT U113 ( .A1(n157), .A2(i_data_bus[216]), .B1(n156), .B2(
        i_data_bus[184]), .ZN(n84) );
  IOA21D1BWP30P140LVT U114 ( .A1(n17), .A2(i_data_bus[248]), .B(n84), .ZN(n85)
         );
  AOI21D1BWP30P140LVT U115 ( .A1(n2), .A2(i_data_bus[24]), .B(n85), .ZN(n88)
         );
  AOI22D1BWP30P140LVT U116 ( .A1(n138), .A2(i_data_bus[88]), .B1(n160), .B2(
        i_data_bus[56]), .ZN(n87) );
  AOI22D1BWP30P140LVT U117 ( .A1(n3), .A2(i_data_bus[120]), .B1(n162), .B2(
        i_data_bus[152]), .ZN(n86) );
  ND3D1BWP30P140LVT U118 ( .A1(n88), .A2(n87), .A3(n86), .ZN(N393) );
  AOI22D1BWP30P140LVT U119 ( .A1(n157), .A2(i_data_bus[210]), .B1(n156), .B2(
        i_data_bus[178]), .ZN(n89) );
  IOA21D1BWP30P140LVT U120 ( .A1(n17), .A2(i_data_bus[242]), .B(n89), .ZN(n90)
         );
  AOI21D1BWP30P140LVT U121 ( .A1(n2), .A2(i_data_bus[18]), .B(n90), .ZN(n93)
         );
  AOI22D1BWP30P140LVT U122 ( .A1(n138), .A2(i_data_bus[82]), .B1(n160), .B2(
        i_data_bus[50]), .ZN(n92) );
  AOI22D1BWP30P140LVT U123 ( .A1(n3), .A2(i_data_bus[114]), .B1(n162), .B2(
        i_data_bus[146]), .ZN(n91) );
  ND3D1BWP30P140LVT U124 ( .A1(n93), .A2(n92), .A3(n91), .ZN(N387) );
  AOI22D1BWP30P140LVT U125 ( .A1(n157), .A2(i_data_bus[211]), .B1(n156), .B2(
        i_data_bus[179]), .ZN(n94) );
  IOA21D1BWP30P140LVT U126 ( .A1(n17), .A2(i_data_bus[243]), .B(n94), .ZN(n95)
         );
  AOI21D1BWP30P140LVT U127 ( .A1(n2), .A2(i_data_bus[19]), .B(n95), .ZN(n98)
         );
  AOI22D1BWP30P140LVT U128 ( .A1(n138), .A2(i_data_bus[83]), .B1(n160), .B2(
        i_data_bus[51]), .ZN(n97) );
  AOI22D1BWP30P140LVT U129 ( .A1(n3), .A2(i_data_bus[115]), .B1(n162), .B2(
        i_data_bus[147]), .ZN(n96) );
  ND3D1BWP30P140LVT U130 ( .A1(n98), .A2(n97), .A3(n96), .ZN(N388) );
  AOI22D1BWP30P140LVT U131 ( .A1(n157), .A2(i_data_bus[212]), .B1(n156), .B2(
        i_data_bus[180]), .ZN(n99) );
  IOA21D1BWP30P140LVT U132 ( .A1(n17), .A2(i_data_bus[244]), .B(n99), .ZN(n100) );
  AOI21D1BWP30P140LVT U133 ( .A1(n2), .A2(i_data_bus[20]), .B(n100), .ZN(n103)
         );
  AOI22D1BWP30P140LVT U134 ( .A1(n138), .A2(i_data_bus[84]), .B1(n160), .B2(
        i_data_bus[52]), .ZN(n102) );
  AOI22D1BWP30P140LVT U135 ( .A1(n3), .A2(i_data_bus[116]), .B1(n162), .B2(
        i_data_bus[148]), .ZN(n101) );
  ND3D1BWP30P140LVT U136 ( .A1(n103), .A2(n102), .A3(n101), .ZN(N389) );
  AOI22D1BWP30P140LVT U137 ( .A1(n157), .A2(i_data_bus[213]), .B1(n156), .B2(
        i_data_bus[181]), .ZN(n104) );
  IOA21D1BWP30P140LVT U138 ( .A1(n17), .A2(i_data_bus[245]), .B(n104), .ZN(
        n105) );
  AOI21D1BWP30P140LVT U139 ( .A1(n2), .A2(i_data_bus[21]), .B(n105), .ZN(n108)
         );
  AOI22D1BWP30P140LVT U140 ( .A1(n138), .A2(i_data_bus[85]), .B1(n160), .B2(
        i_data_bus[53]), .ZN(n107) );
  AOI22D1BWP30P140LVT U141 ( .A1(n3), .A2(i_data_bus[117]), .B1(n162), .B2(
        i_data_bus[149]), .ZN(n106) );
  ND3D1BWP30P140LVT U142 ( .A1(n108), .A2(n107), .A3(n106), .ZN(N390) );
  AOI22D1BWP30P140LVT U143 ( .A1(n157), .A2(i_data_bus[208]), .B1(n156), .B2(
        i_data_bus[176]), .ZN(n109) );
  IOA21D1BWP30P140LVT U144 ( .A1(n17), .A2(i_data_bus[240]), .B(n109), .ZN(
        n110) );
  AOI21D1BWP30P140LVT U145 ( .A1(n2), .A2(i_data_bus[16]), .B(n110), .ZN(n113)
         );
  AOI22D1BWP30P140LVT U146 ( .A1(n138), .A2(i_data_bus[80]), .B1(n160), .B2(
        i_data_bus[48]), .ZN(n112) );
  AOI22D1BWP30P140LVT U147 ( .A1(n3), .A2(i_data_bus[112]), .B1(n162), .B2(
        i_data_bus[144]), .ZN(n111) );
  ND3D1BWP30P140LVT U148 ( .A1(n113), .A2(n112), .A3(n111), .ZN(N385) );
  AOI22D1BWP30P140LVT U149 ( .A1(n217), .A2(i_data_bus[207]), .B1(n156), .B2(
        i_data_bus[175]), .ZN(n114) );
  IOA21D1BWP30P140LVT U150 ( .A1(n17), .A2(i_data_bus[239]), .B(n114), .ZN(
        n115) );
  AOI21D1BWP30P140LVT U151 ( .A1(n2), .A2(i_data_bus[15]), .B(n115), .ZN(n118)
         );
  AOI22D1BWP30P140LVT U152 ( .A1(n138), .A2(i_data_bus[79]), .B1(n160), .B2(
        i_data_bus[47]), .ZN(n117) );
  AOI22D1BWP30P140LVT U153 ( .A1(n3), .A2(i_data_bus[111]), .B1(n162), .B2(
        i_data_bus[143]), .ZN(n116) );
  ND3D1BWP30P140LVT U154 ( .A1(n118), .A2(n117), .A3(n116), .ZN(N384) );
  AOI22D1BWP30P140LVT U155 ( .A1(n217), .A2(i_data_bus[206]), .B1(n156), .B2(
        i_data_bus[174]), .ZN(n119) );
  IOA21D1BWP30P140LVT U156 ( .A1(n17), .A2(i_data_bus[238]), .B(n119), .ZN(
        n120) );
  AOI21D1BWP30P140LVT U157 ( .A1(n2), .A2(i_data_bus[14]), .B(n120), .ZN(n123)
         );
  AOI22D1BWP30P140LVT U158 ( .A1(n138), .A2(i_data_bus[78]), .B1(n160), .B2(
        i_data_bus[46]), .ZN(n122) );
  AOI22D1BWP30P140LVT U159 ( .A1(n3), .A2(i_data_bus[110]), .B1(n162), .B2(
        i_data_bus[142]), .ZN(n121) );
  ND3D1BWP30P140LVT U160 ( .A1(n123), .A2(n122), .A3(n121), .ZN(N383) );
  AOI22D1BWP30P140LVT U161 ( .A1(n157), .A2(i_data_bus[217]), .B1(n156), .B2(
        i_data_bus[185]), .ZN(n124) );
  IOA21D1BWP30P140LVT U162 ( .A1(n17), .A2(i_data_bus[249]), .B(n124), .ZN(
        n125) );
  AOI21D1BWP30P140LVT U163 ( .A1(n2), .A2(i_data_bus[25]), .B(n125), .ZN(n128)
         );
  AOI22D1BWP30P140LVT U164 ( .A1(n138), .A2(i_data_bus[89]), .B1(n160), .B2(
        i_data_bus[57]), .ZN(n127) );
  AOI22D1BWP30P140LVT U165 ( .A1(n3), .A2(i_data_bus[121]), .B1(n162), .B2(
        i_data_bus[153]), .ZN(n126) );
  ND3D1BWP30P140LVT U166 ( .A1(n128), .A2(n127), .A3(n126), .ZN(N394) );
  INVD1BWP30P140LVT U167 ( .I(i_data_bus[173]), .ZN(n129) );
  IOA21D1BWP30P140LVT U168 ( .A1(n17), .A2(i_data_bus[237]), .B(n131), .ZN(
        n132) );
  AOI21D1BWP30P140LVT U169 ( .A1(n2), .A2(i_data_bus[13]), .B(n132), .ZN(n135)
         );
  AOI22D1BWP30P140LVT U170 ( .A1(n138), .A2(i_data_bus[77]), .B1(n160), .B2(
        i_data_bus[45]), .ZN(n134) );
  AOI22D1BWP30P140LVT U171 ( .A1(n3), .A2(i_data_bus[109]), .B1(n162), .B2(
        i_data_bus[141]), .ZN(n133) );
  ND3D1BWP30P140LVT U172 ( .A1(n135), .A2(n134), .A3(n133), .ZN(N382) );
  AOI22D1BWP30P140LVT U173 ( .A1(n157), .A2(i_data_bus[209]), .B1(n156), .B2(
        i_data_bus[177]), .ZN(n136) );
  IOA21D1BWP30P140LVT U174 ( .A1(n17), .A2(i_data_bus[241]), .B(n136), .ZN(
        n137) );
  AOI21D1BWP30P140LVT U175 ( .A1(n2), .A2(i_data_bus[17]), .B(n137), .ZN(n141)
         );
  AOI22D1BWP30P140LVT U176 ( .A1(n138), .A2(i_data_bus[81]), .B1(n160), .B2(
        i_data_bus[49]), .ZN(n140) );
  AOI22D1BWP30P140LVT U177 ( .A1(n3), .A2(i_data_bus[113]), .B1(n162), .B2(
        i_data_bus[145]), .ZN(n139) );
  ND3D1BWP30P140LVT U178 ( .A1(n141), .A2(n140), .A3(n139), .ZN(N386) );
  AOI22D1BWP30P140LVT U179 ( .A1(n157), .A2(i_data_bus[223]), .B1(n156), .B2(
        i_data_bus[191]), .ZN(n142) );
  IOA21D1BWP30P140LVT U180 ( .A1(n17), .A2(i_data_bus[255]), .B(n142), .ZN(
        n143) );
  AOI22D1BWP30P140LVT U181 ( .A1(n161), .A2(i_data_bus[95]), .B1(n160), .B2(
        i_data_bus[63]), .ZN(n149) );
  INVD1BWP30P140LVT U182 ( .I(i_data_bus[127]), .ZN(n146) );
  INVD1BWP30P140LVT U183 ( .I(i_data_bus[159]), .ZN(n144) );
  OA22D1BWP30P140LVT U184 ( .A1(n147), .A2(n146), .B1(n145), .B2(n144), .Z(
        n148) );
  ND3D1BWP30P140LVT U185 ( .A1(n150), .A2(n149), .A3(n148), .ZN(N400) );
  AOI22D1BWP30P140LVT U186 ( .A1(n157), .A2(i_data_bus[222]), .B1(n156), .B2(
        i_data_bus[190]), .ZN(n151) );
  IOA21D1BWP30P140LVT U187 ( .A1(n17), .A2(i_data_bus[254]), .B(n151), .ZN(
        n152) );
  AOI22D1BWP30P140LVT U188 ( .A1(n161), .A2(i_data_bus[94]), .B1(n160), .B2(
        i_data_bus[62]), .ZN(n154) );
  AOI22D1BWP30P140LVT U189 ( .A1(n3), .A2(i_data_bus[126]), .B1(n162), .B2(
        i_data_bus[158]), .ZN(n153) );
  ND3D1BWP30P140LVT U190 ( .A1(n155), .A2(n154), .A3(n153), .ZN(N399) );
  AOI22D1BWP30P140LVT U191 ( .A1(n157), .A2(i_data_bus[220]), .B1(n156), .B2(
        i_data_bus[188]), .ZN(n158) );
  IOA21D1BWP30P140LVT U192 ( .A1(n17), .A2(i_data_bus[252]), .B(n158), .ZN(
        n159) );
  AOI22D1BWP30P140LVT U193 ( .A1(n161), .A2(i_data_bus[92]), .B1(n160), .B2(
        i_data_bus[60]), .ZN(n164) );
  AOI22D1BWP30P140LVT U194 ( .A1(n3), .A2(i_data_bus[124]), .B1(n162), .B2(
        i_data_bus[156]), .ZN(n163) );
  ND3D1BWP30P140LVT U195 ( .A1(n165), .A2(n164), .A3(n163), .ZN(N397) );
  AOI22D1BWP30P140LVT U196 ( .A1(n217), .A2(i_data_bus[204]), .B1(n216), .B2(
        i_data_bus[172]), .ZN(n166) );
  IOA21D1BWP30P140LVT U197 ( .A1(n17), .A2(i_data_bus[236]), .B(n166), .ZN(
        n167) );
  AOI21D1BWP30P140LVT U198 ( .A1(n2), .A2(i_data_bus[12]), .B(n167), .ZN(n170)
         );
  AOI22D1BWP30P140LVT U199 ( .A1(n221), .A2(i_data_bus[76]), .B1(n220), .B2(
        i_data_bus[44]), .ZN(n169) );
  AOI22D1BWP30P140LVT U200 ( .A1(n223), .A2(i_data_bus[108]), .B1(n222), .B2(
        i_data_bus[140]), .ZN(n168) );
  ND3D1BWP30P140LVT U201 ( .A1(n170), .A2(n169), .A3(n168), .ZN(N381) );
  AOI22D1BWP30P140LVT U202 ( .A1(n217), .A2(i_data_bus[203]), .B1(n216), .B2(
        i_data_bus[171]), .ZN(n171) );
  IOA21D1BWP30P140LVT U203 ( .A1(n17), .A2(i_data_bus[235]), .B(n171), .ZN(
        n172) );
  AOI21D1BWP30P140LVT U204 ( .A1(n2), .A2(i_data_bus[11]), .B(n172), .ZN(n175)
         );
  AOI22D1BWP30P140LVT U205 ( .A1(n221), .A2(i_data_bus[75]), .B1(n220), .B2(
        i_data_bus[43]), .ZN(n174) );
  AOI22D1BWP30P140LVT U206 ( .A1(n223), .A2(i_data_bus[107]), .B1(n222), .B2(
        i_data_bus[139]), .ZN(n173) );
  ND3D1BWP30P140LVT U207 ( .A1(n175), .A2(n174), .A3(n173), .ZN(N380) );
  AOI22D1BWP30P140LVT U208 ( .A1(n217), .A2(i_data_bus[202]), .B1(n216), .B2(
        i_data_bus[170]), .ZN(n176) );
  IOA21D1BWP30P140LVT U209 ( .A1(n17), .A2(i_data_bus[234]), .B(n176), .ZN(
        n177) );
  AOI21D1BWP30P140LVT U210 ( .A1(n2), .A2(i_data_bus[10]), .B(n177), .ZN(n180)
         );
  AOI22D1BWP30P140LVT U211 ( .A1(n221), .A2(i_data_bus[74]), .B1(n220), .B2(
        i_data_bus[42]), .ZN(n179) );
  AOI22D1BWP30P140LVT U212 ( .A1(n223), .A2(i_data_bus[106]), .B1(n222), .B2(
        i_data_bus[138]), .ZN(n178) );
  ND3D1BWP30P140LVT U213 ( .A1(n180), .A2(n179), .A3(n178), .ZN(N379) );
  AOI22D1BWP30P140LVT U214 ( .A1(n217), .A2(i_data_bus[201]), .B1(n216), .B2(
        i_data_bus[169]), .ZN(n181) );
  IOA21D1BWP30P140LVT U215 ( .A1(n17), .A2(i_data_bus[233]), .B(n181), .ZN(
        n182) );
  AOI21D1BWP30P140LVT U216 ( .A1(n2), .A2(i_data_bus[9]), .B(n182), .ZN(n185)
         );
  AOI22D1BWP30P140LVT U217 ( .A1(n221), .A2(i_data_bus[73]), .B1(n220), .B2(
        i_data_bus[41]), .ZN(n184) );
  AOI22D1BWP30P140LVT U218 ( .A1(n223), .A2(i_data_bus[105]), .B1(n222), .B2(
        i_data_bus[137]), .ZN(n183) );
  ND3D1BWP30P140LVT U219 ( .A1(n185), .A2(n184), .A3(n183), .ZN(N378) );
  AOI22D1BWP30P140LVT U220 ( .A1(n217), .A2(i_data_bus[200]), .B1(n216), .B2(
        i_data_bus[168]), .ZN(n186) );
  IOA21D1BWP30P140LVT U221 ( .A1(n17), .A2(i_data_bus[232]), .B(n186), .ZN(
        n187) );
  AOI21D1BWP30P140LVT U222 ( .A1(n2), .A2(i_data_bus[8]), .B(n187), .ZN(n190)
         );
  AOI22D1BWP30P140LVT U223 ( .A1(n221), .A2(i_data_bus[72]), .B1(n220), .B2(
        i_data_bus[40]), .ZN(n189) );
  AOI22D1BWP30P140LVT U224 ( .A1(n223), .A2(i_data_bus[104]), .B1(n222), .B2(
        i_data_bus[136]), .ZN(n188) );
  ND3D1BWP30P140LVT U225 ( .A1(n190), .A2(n189), .A3(n188), .ZN(N377) );
  AOI22D1BWP30P140LVT U226 ( .A1(n217), .A2(i_data_bus[198]), .B1(n216), .B2(
        i_data_bus[166]), .ZN(n191) );
  IOA21D1BWP30P140LVT U227 ( .A1(n17), .A2(i_data_bus[230]), .B(n191), .ZN(
        n192) );
  AOI21D1BWP30P140LVT U228 ( .A1(n2), .A2(i_data_bus[6]), .B(n192), .ZN(n195)
         );
  AOI22D1BWP30P140LVT U229 ( .A1(n221), .A2(i_data_bus[70]), .B1(n220), .B2(
        i_data_bus[38]), .ZN(n194) );
  AOI22D1BWP30P140LVT U230 ( .A1(n223), .A2(i_data_bus[102]), .B1(n222), .B2(
        i_data_bus[134]), .ZN(n193) );
  ND3D1BWP30P140LVT U231 ( .A1(n195), .A2(n194), .A3(n193), .ZN(N375) );
  AOI22D1BWP30P140LVT U232 ( .A1(n217), .A2(i_data_bus[197]), .B1(n216), .B2(
        i_data_bus[165]), .ZN(n196) );
  IOA21D1BWP30P140LVT U233 ( .A1(n17), .A2(i_data_bus[229]), .B(n196), .ZN(
        n197) );
  AOI21D1BWP30P140LVT U234 ( .A1(n2), .A2(i_data_bus[5]), .B(n197), .ZN(n200)
         );
  AOI22D1BWP30P140LVT U235 ( .A1(n221), .A2(i_data_bus[69]), .B1(n220), .B2(
        i_data_bus[37]), .ZN(n199) );
  AOI22D1BWP30P140LVT U236 ( .A1(n223), .A2(i_data_bus[101]), .B1(n222), .B2(
        i_data_bus[133]), .ZN(n198) );
  ND3D1BWP30P140LVT U237 ( .A1(n200), .A2(n199), .A3(n198), .ZN(N374) );
  AOI22D1BWP30P140LVT U238 ( .A1(n217), .A2(i_data_bus[196]), .B1(n216), .B2(
        i_data_bus[164]), .ZN(n201) );
  IOA21D1BWP30P140LVT U239 ( .A1(n17), .A2(i_data_bus[228]), .B(n201), .ZN(
        n202) );
  AOI21D1BWP30P140LVT U240 ( .A1(n2), .A2(i_data_bus[4]), .B(n202), .ZN(n205)
         );
  AOI22D1BWP30P140LVT U241 ( .A1(n221), .A2(i_data_bus[68]), .B1(n220), .B2(
        i_data_bus[36]), .ZN(n204) );
  AOI22D1BWP30P140LVT U242 ( .A1(n223), .A2(i_data_bus[100]), .B1(n222), .B2(
        i_data_bus[132]), .ZN(n203) );
  ND3D1BWP30P140LVT U243 ( .A1(n205), .A2(n204), .A3(n203), .ZN(N373) );
  AOI22D1BWP30P140LVT U244 ( .A1(n217), .A2(i_data_bus[195]), .B1(n216), .B2(
        i_data_bus[163]), .ZN(n206) );
  IOA21D1BWP30P140LVT U245 ( .A1(n17), .A2(i_data_bus[227]), .B(n206), .ZN(
        n207) );
  AOI21D1BWP30P140LVT U246 ( .A1(n2), .A2(i_data_bus[3]), .B(n207), .ZN(n210)
         );
  AOI22D1BWP30P140LVT U247 ( .A1(n221), .A2(i_data_bus[67]), .B1(n220), .B2(
        i_data_bus[35]), .ZN(n209) );
  AOI22D1BWP30P140LVT U248 ( .A1(n223), .A2(i_data_bus[99]), .B1(n222), .B2(
        i_data_bus[131]), .ZN(n208) );
  ND3D1BWP30P140LVT U249 ( .A1(n210), .A2(n209), .A3(n208), .ZN(N372) );
  AOI22D1BWP30P140LVT U250 ( .A1(n217), .A2(i_data_bus[194]), .B1(n216), .B2(
        i_data_bus[162]), .ZN(n211) );
  IOA21D1BWP30P140LVT U251 ( .A1(n17), .A2(i_data_bus[226]), .B(n211), .ZN(
        n212) );
  AOI21D1BWP30P140LVT U252 ( .A1(n2), .A2(i_data_bus[2]), .B(n212), .ZN(n215)
         );
  AOI22D1BWP30P140LVT U253 ( .A1(n221), .A2(i_data_bus[66]), .B1(n220), .B2(
        i_data_bus[34]), .ZN(n214) );
  AOI22D1BWP30P140LVT U254 ( .A1(n223), .A2(i_data_bus[98]), .B1(n222), .B2(
        i_data_bus[130]), .ZN(n213) );
  ND3D1BWP30P140LVT U255 ( .A1(n215), .A2(n214), .A3(n213), .ZN(N371) );
  AOI22D1BWP30P140LVT U256 ( .A1(n217), .A2(i_data_bus[199]), .B1(n216), .B2(
        i_data_bus[167]), .ZN(n218) );
  IOA21D1BWP30P140LVT U257 ( .A1(n17), .A2(i_data_bus[231]), .B(n218), .ZN(
        n219) );
  AOI21D1BWP30P140LVT U258 ( .A1(n2), .A2(i_data_bus[7]), .B(n219), .ZN(n226)
         );
  AOI22D1BWP30P140LVT U259 ( .A1(n221), .A2(i_data_bus[71]), .B1(n220), .B2(
        i_data_bus[39]), .ZN(n225) );
  AOI22D1BWP30P140LVT U260 ( .A1(n223), .A2(i_data_bus[103]), .B1(n222), .B2(
        i_data_bus[135]), .ZN(n224) );
  ND3D1BWP30P140LVT U261 ( .A1(n226), .A2(n225), .A3(n224), .ZN(N376) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_1 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD3BWP30P140LVT U3 ( .I(n146), .ZN(n2) );
  INVD1BWP30P140LVT U4 ( .I(n145), .ZN(n114) );
  OR2D1BWP30P140LVT U5 ( .A1(n20), .A2(n19), .Z(n21) );
  INVD4BWP30P140LVT U6 ( .I(n40), .ZN(n216) );
  INVD4BWP30P140LVT U7 ( .I(n54), .ZN(n3) );
  OR2D1BWP30P140LVT U8 ( .A1(n39), .A2(n38), .Z(n40) );
  NR3D1P5BWP30P140LVT U9 ( .A1(i_cmd[6]), .A2(i_cmd[5]), .A3(i_cmd[7]), .ZN(n9) );
  INR2D1BWP30P140LVT U10 ( .A1(n11), .B1(n10), .ZN(n23) );
  CKAN2D4BWP30P140LVT U11 ( .A1(n23), .A2(n13), .Z(n1) );
  INVD6BWP30P140LVT U12 ( .I(n21), .ZN(n219) );
  NR3D0P7BWP30P140LVT U13 ( .A1(n24), .A2(i_cmd[5]), .A3(i_cmd[7]), .ZN(n30)
         );
  ND2D1BWP30P140LVT U14 ( .A1(i_valid[6]), .A2(i_cmd[6]), .ZN(n24) );
  INVD1BWP30P140LVT U15 ( .I(n49), .ZN(n50) );
  OAI21D1BWP30P140LVT U16 ( .A1(n183), .A2(n42), .B(n41), .ZN(n43) );
  INVD1BWP30P140LVT U17 ( .I(i_data_bus[160]), .ZN(n42) );
  ND2D1BWP30P140LVT U18 ( .A1(n216), .A2(i_data_bus[224]), .ZN(n41) );
  INVD1BWP30P140LVT U19 ( .I(i_data_bus[192]), .ZN(n32) );
  INVD1BWP30P140LVT U20 ( .I(i_valid[5]), .ZN(n33) );
  OR2D2BWP30P140LVT U21 ( .A1(n29), .A2(n28), .Z(n38) );
  ND3D1BWP30P140LVT U22 ( .A1(n48), .A2(n47), .A3(n46), .ZN(N369) );
  NR3D0P7BWP30P140LVT U23 ( .A1(n45), .A2(n44), .A3(n43), .ZN(n46) );
  NR2D1BWP30P140LVT U24 ( .A1(n2), .A2(n1), .ZN(n51) );
  OR2D1BWP30P140LVT U25 ( .A1(n20), .A2(n6), .Z(n146) );
  OR2D1BWP30P140LVT U26 ( .A1(n20), .A2(n16), .Z(n145) );
  IND2D1BWP30P140LVT U27 ( .A1(rst), .B1(i_en), .ZN(n7) );
  NR2OPTPAD1BWP30P140LVT U28 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n27) );
  IND3D1BWP30P140LVT U29 ( .A1(n7), .B1(n27), .B2(n9), .ZN(n20) );
  INVD1BWP30P140LVT U30 ( .I(i_cmd[2]), .ZN(n4) );
  INVD1BWP30P140LVT U31 ( .I(i_cmd[1]), .ZN(n15) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n4), .A2(n15), .ZN(n29) );
  INVD1BWP30P140LVT U33 ( .I(n29), .ZN(n5) );
  ND3D1BWP30P140LVT U34 ( .A1(n5), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n6) );
  OR2D4BWP30P140LVT U35 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n17) );
  NR2D1BWP30P140LVT U36 ( .A1(n17), .A2(i_cmd[1]), .ZN(n11) );
  INVD1BWP30P140LVT U37 ( .I(n7), .ZN(n8) );
  ND2OPTIBD1BWP30P140LVT U38 ( .A1(n9), .A2(n8), .ZN(n10) );
  IND3D1BWP30P140LVT U39 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n12) );
  INVD1BWP30P140LVT U40 ( .I(n12), .ZN(n13) );
  AOI22D1BWP30P140LVT U41 ( .A1(n2), .A2(i_data_bus[96]), .B1(n1), .B2(
        i_data_bus[128]), .ZN(n48) );
  INVD1BWP30P140LVT U42 ( .I(i_cmd[3]), .ZN(n14) );
  ND4D1BWP30P140LVT U43 ( .A1(n15), .A2(n14), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n16) );
  INVD1BWP30P140LVT U44 ( .I(n17), .ZN(n18) );
  ND3D1BWP30P140LVT U45 ( .A1(n18), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n19)
         );
  AOI22D1BWP30P140LVT U46 ( .A1(n114), .A2(i_data_bus[64]), .B1(n219), .B2(
        i_data_bus[32]), .ZN(n47) );
  INR2D1BWP30P140LVT U47 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n22) );
  ND3D1BWP30P140LVT U48 ( .A1(n23), .A2(i_cmd[0]), .A3(n22), .ZN(n49) );
  INR2D1BWP30P140LVT U49 ( .A1(i_data_bus[0]), .B1(n49), .ZN(n45) );
  INR2D1BWP30P140LVT U50 ( .A1(i_en), .B1(rst), .ZN(n25) );
  INR2D1BWP30P140LVT U51 ( .A1(n25), .B1(i_cmd[3]), .ZN(n26) );
  ND2OPTIBD1BWP30P140LVT U52 ( .A1(n27), .A2(n26), .ZN(n28) );
  INR2D1BWP30P140LVT U53 ( .A1(n30), .B1(n38), .ZN(n31) );
  INVD2BWP30P140LVT U54 ( .I(n31), .ZN(n54) );
  NR2D1BWP30P140LVT U55 ( .A1(n54), .A2(n32), .ZN(n44) );
  INVD1BWP30P140LVT U56 ( .I(i_cmd[5]), .ZN(n34) );
  NR4D1BWP30P140LVT U57 ( .A1(n34), .A2(n33), .A3(i_cmd[6]), .A4(i_cmd[7]), 
        .ZN(n35) );
  INR2D2BWP30P140LVT U58 ( .A1(n35), .B1(n38), .ZN(n36) );
  INVD2BWP30P140LVT U59 ( .I(n36), .ZN(n183) );
  ND2D1BWP30P140LVT U60 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n37) );
  OR3D1BWP30P140LVT U61 ( .A1(n37), .A2(i_cmd[5]), .A3(i_cmd[6]), .Z(n39) );
  INVD2BWP30P140LVT U62 ( .I(n50), .ZN(n156) );
  INVD2BWP30P140LVT U63 ( .I(n156), .ZN(n152) );
  INVD3BWP30P140LVT U64 ( .I(n183), .ZN(n214) );
  NR4D0BWP30P140LVT U65 ( .A1(n152), .A2(n216), .A3(n3), .A4(n214), .ZN(n53)
         );
  NR2D1BWP30P140LVT U66 ( .A1(n220), .A2(n219), .ZN(n52) );
  ND3D1BWP30P140LVT U67 ( .A1(n53), .A2(n52), .A3(n51), .ZN(N402) );
  INVD2BWP30P140LVT U68 ( .I(n156), .ZN(n113) );
  INVD2BWP30P140LVT U69 ( .I(n183), .ZN(n110) );
  AOI22D1BWP30P140LVT U70 ( .A1(n3), .A2(i_data_bus[204]), .B1(n110), .B2(
        i_data_bus[172]), .ZN(n55) );
  IOA21D1BWP30P140LVT U71 ( .A1(n216), .A2(i_data_bus[236]), .B(n55), .ZN(n56)
         );
  AOI21D1BWP30P140LVT U72 ( .A1(n113), .A2(i_data_bus[12]), .B(n56), .ZN(n59)
         );
  AOI22D1BWP30P140LVT U73 ( .A1(n114), .A2(i_data_bus[76]), .B1(n219), .B2(
        i_data_bus[44]), .ZN(n58) );
  AOI22D1BWP30P140LVT U74 ( .A1(n2), .A2(i_data_bus[108]), .B1(n1), .B2(
        i_data_bus[140]), .ZN(n57) );
  ND3D1BWP30P140LVT U75 ( .A1(n59), .A2(n58), .A3(n57), .ZN(N381) );
  AOI22D1BWP30P140LVT U76 ( .A1(n3), .A2(i_data_bus[194]), .B1(n110), .B2(
        i_data_bus[162]), .ZN(n60) );
  IOA21D1BWP30P140LVT U77 ( .A1(n216), .A2(i_data_bus[226]), .B(n60), .ZN(n61)
         );
  AOI21D1BWP30P140LVT U78 ( .A1(n113), .A2(i_data_bus[2]), .B(n61), .ZN(n64)
         );
  AOI22D1BWP30P140LVT U79 ( .A1(n114), .A2(i_data_bus[66]), .B1(n219), .B2(
        i_data_bus[34]), .ZN(n63) );
  AOI22D1BWP30P140LVT U80 ( .A1(n2), .A2(i_data_bus[98]), .B1(n1), .B2(
        i_data_bus[130]), .ZN(n62) );
  ND3D1BWP30P140LVT U81 ( .A1(n64), .A2(n63), .A3(n62), .ZN(N371) );
  AOI22D1BWP30P140LVT U82 ( .A1(n3), .A2(i_data_bus[196]), .B1(n110), .B2(
        i_data_bus[164]), .ZN(n65) );
  IOA21D1BWP30P140LVT U83 ( .A1(n216), .A2(i_data_bus[228]), .B(n65), .ZN(n66)
         );
  AOI21D1BWP30P140LVT U84 ( .A1(n113), .A2(i_data_bus[4]), .B(n66), .ZN(n69)
         );
  AOI22D1BWP30P140LVT U85 ( .A1(n114), .A2(i_data_bus[68]), .B1(n219), .B2(
        i_data_bus[36]), .ZN(n68) );
  AOI22D1BWP30P140LVT U86 ( .A1(n2), .A2(i_data_bus[100]), .B1(n1), .B2(
        i_data_bus[132]), .ZN(n67) );
  ND3D1BWP30P140LVT U87 ( .A1(n69), .A2(n68), .A3(n67), .ZN(N373) );
  AOI22D1BWP30P140LVT U88 ( .A1(n3), .A2(i_data_bus[197]), .B1(n110), .B2(
        i_data_bus[165]), .ZN(n70) );
  IOA21D1BWP30P140LVT U89 ( .A1(n216), .A2(i_data_bus[229]), .B(n70), .ZN(n71)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n113), .A2(i_data_bus[5]), .B(n71), .ZN(n74)
         );
  AOI22D1BWP30P140LVT U91 ( .A1(n114), .A2(i_data_bus[69]), .B1(n219), .B2(
        i_data_bus[37]), .ZN(n73) );
  AOI22D1BWP30P140LVT U92 ( .A1(n2), .A2(i_data_bus[101]), .B1(n1), .B2(
        i_data_bus[133]), .ZN(n72) );
  ND3D1BWP30P140LVT U93 ( .A1(n74), .A2(n73), .A3(n72), .ZN(N374) );
  AOI22D1BWP30P140LVT U94 ( .A1(n3), .A2(i_data_bus[198]), .B1(n110), .B2(
        i_data_bus[166]), .ZN(n75) );
  IOA21D1BWP30P140LVT U95 ( .A1(n216), .A2(i_data_bus[230]), .B(n75), .ZN(n76)
         );
  AOI21D1BWP30P140LVT U96 ( .A1(n113), .A2(i_data_bus[6]), .B(n76), .ZN(n79)
         );
  AOI22D1BWP30P140LVT U97 ( .A1(n114), .A2(i_data_bus[70]), .B1(n219), .B2(
        i_data_bus[38]), .ZN(n78) );
  AOI22D1BWP30P140LVT U98 ( .A1(n2), .A2(i_data_bus[102]), .B1(n1), .B2(
        i_data_bus[134]), .ZN(n77) );
  ND3D1BWP30P140LVT U99 ( .A1(n79), .A2(n78), .A3(n77), .ZN(N375) );
  AOI22D1BWP30P140LVT U100 ( .A1(n3), .A2(i_data_bus[195]), .B1(n110), .B2(
        i_data_bus[163]), .ZN(n80) );
  IOA21D1BWP30P140LVT U101 ( .A1(n216), .A2(i_data_bus[227]), .B(n80), .ZN(n81) );
  AOI21D1BWP30P140LVT U102 ( .A1(n113), .A2(i_data_bus[3]), .B(n81), .ZN(n84)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n114), .A2(i_data_bus[67]), .B1(n219), .B2(
        i_data_bus[35]), .ZN(n83) );
  AOI22D1BWP30P140LVT U104 ( .A1(n2), .A2(i_data_bus[99]), .B1(n1), .B2(
        i_data_bus[131]), .ZN(n82) );
  ND3D1BWP30P140LVT U105 ( .A1(n84), .A2(n83), .A3(n82), .ZN(N372) );
  AOI22D1BWP30P140LVT U106 ( .A1(n3), .A2(i_data_bus[193]), .B1(n110), .B2(
        i_data_bus[161]), .ZN(n85) );
  IOA21D1BWP30P140LVT U107 ( .A1(n216), .A2(i_data_bus[225]), .B(n85), .ZN(n86) );
  AOI21D1BWP30P140LVT U108 ( .A1(n113), .A2(i_data_bus[1]), .B(n86), .ZN(n89)
         );
  AOI22D1BWP30P140LVT U109 ( .A1(n114), .A2(i_data_bus[65]), .B1(n219), .B2(
        i_data_bus[33]), .ZN(n88) );
  AOI22D1BWP30P140LVT U110 ( .A1(n2), .A2(i_data_bus[97]), .B1(n1), .B2(
        i_data_bus[129]), .ZN(n87) );
  ND3D1BWP30P140LVT U111 ( .A1(n89), .A2(n88), .A3(n87), .ZN(N370) );
  AOI22D1BWP30P140LVT U112 ( .A1(n3), .A2(i_data_bus[200]), .B1(n110), .B2(
        i_data_bus[168]), .ZN(n90) );
  IOA21D1BWP30P140LVT U113 ( .A1(n216), .A2(i_data_bus[232]), .B(n90), .ZN(n91) );
  AOI21D1BWP30P140LVT U114 ( .A1(n113), .A2(i_data_bus[8]), .B(n91), .ZN(n94)
         );
  AOI22D1BWP30P140LVT U115 ( .A1(n114), .A2(i_data_bus[72]), .B1(n219), .B2(
        i_data_bus[40]), .ZN(n93) );
  AOI22D1BWP30P140LVT U116 ( .A1(n2), .A2(i_data_bus[104]), .B1(n1), .B2(
        i_data_bus[136]), .ZN(n92) );
  ND3D1BWP30P140LVT U117 ( .A1(n94), .A2(n93), .A3(n92), .ZN(N377) );
  AOI22D1BWP30P140LVT U118 ( .A1(n3), .A2(i_data_bus[199]), .B1(n110), .B2(
        i_data_bus[167]), .ZN(n95) );
  IOA21D1BWP30P140LVT U119 ( .A1(n216), .A2(i_data_bus[231]), .B(n95), .ZN(n96) );
  AOI21D1BWP30P140LVT U120 ( .A1(n113), .A2(i_data_bus[7]), .B(n96), .ZN(n99)
         );
  AOI22D1BWP30P140LVT U121 ( .A1(n114), .A2(i_data_bus[71]), .B1(n219), .B2(
        i_data_bus[39]), .ZN(n98) );
  AOI22D1BWP30P140LVT U122 ( .A1(n2), .A2(i_data_bus[103]), .B1(n1), .B2(
        i_data_bus[135]), .ZN(n97) );
  ND3D1BWP30P140LVT U123 ( .A1(n99), .A2(n98), .A3(n97), .ZN(N376) );
  AOI22D1BWP30P140LVT U124 ( .A1(n3), .A2(i_data_bus[203]), .B1(n110), .B2(
        i_data_bus[171]), .ZN(n100) );
  IOA21D1BWP30P140LVT U125 ( .A1(n216), .A2(i_data_bus[235]), .B(n100), .ZN(
        n101) );
  AOI21D1BWP30P140LVT U126 ( .A1(n113), .A2(i_data_bus[11]), .B(n101), .ZN(
        n104) );
  AOI22D1BWP30P140LVT U127 ( .A1(n114), .A2(i_data_bus[75]), .B1(n219), .B2(
        i_data_bus[43]), .ZN(n103) );
  AOI22D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[107]), .B1(n1), .B2(
        i_data_bus[139]), .ZN(n102) );
  ND3D1BWP30P140LVT U129 ( .A1(n104), .A2(n103), .A3(n102), .ZN(N380) );
  AOI22D1BWP30P140LVT U130 ( .A1(n3), .A2(i_data_bus[202]), .B1(n110), .B2(
        i_data_bus[170]), .ZN(n105) );
  IOA21D1BWP30P140LVT U131 ( .A1(n216), .A2(i_data_bus[234]), .B(n105), .ZN(
        n106) );
  AOI21D1BWP30P140LVT U132 ( .A1(n113), .A2(i_data_bus[10]), .B(n106), .ZN(
        n109) );
  AOI22D1BWP30P140LVT U133 ( .A1(n114), .A2(i_data_bus[74]), .B1(n219), .B2(
        i_data_bus[42]), .ZN(n108) );
  AOI22D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[106]), .B1(n1), .B2(
        i_data_bus[138]), .ZN(n107) );
  ND3D1BWP30P140LVT U135 ( .A1(n109), .A2(n108), .A3(n107), .ZN(N379) );
  AOI22D1BWP30P140LVT U136 ( .A1(n3), .A2(i_data_bus[201]), .B1(n110), .B2(
        i_data_bus[169]), .ZN(n111) );
  IOA21D1BWP30P140LVT U137 ( .A1(n216), .A2(i_data_bus[233]), .B(n111), .ZN(
        n112) );
  AOI21D1BWP30P140LVT U138 ( .A1(n113), .A2(i_data_bus[9]), .B(n112), .ZN(n117) );
  AOI22D1BWP30P140LVT U139 ( .A1(n114), .A2(i_data_bus[73]), .B1(n219), .B2(
        i_data_bus[41]), .ZN(n116) );
  AOI22D1BWP30P140LVT U140 ( .A1(n2), .A2(i_data_bus[105]), .B1(n1), .B2(
        i_data_bus[137]), .ZN(n115) );
  ND3D1BWP30P140LVT U141 ( .A1(n117), .A2(n116), .A3(n115), .ZN(N378) );
  AOI22D1BWP30P140LVT U142 ( .A1(n3), .A2(i_data_bus[222]), .B1(n214), .B2(
        i_data_bus[190]), .ZN(n118) );
  IOA21D1BWP30P140LVT U143 ( .A1(n216), .A2(i_data_bus[254]), .B(n118), .ZN(
        n119) );
  AOI21D1BWP30P140LVT U144 ( .A1(n152), .A2(i_data_bus[30]), .B(n119), .ZN(
        n122) );
  AOI22D1BWP30P140LVT U145 ( .A1(n220), .A2(i_data_bus[94]), .B1(n219), .B2(
        i_data_bus[62]), .ZN(n121) );
  AOI22D1BWP30P140LVT U146 ( .A1(n2), .A2(i_data_bus[126]), .B1(n1), .B2(
        i_data_bus[158]), .ZN(n120) );
  ND3D1BWP30P140LVT U147 ( .A1(n122), .A2(n121), .A3(n120), .ZN(N399) );
  AOI22D1BWP30P140LVT U148 ( .A1(n3), .A2(i_data_bus[221]), .B1(n214), .B2(
        i_data_bus[189]), .ZN(n123) );
  IOA21D1BWP30P140LVT U149 ( .A1(n216), .A2(i_data_bus[253]), .B(n123), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U150 ( .A1(n152), .A2(i_data_bus[29]), .B(n124), .ZN(
        n127) );
  AOI22D1BWP30P140LVT U151 ( .A1(n220), .A2(i_data_bus[93]), .B1(n219), .B2(
        i_data_bus[61]), .ZN(n126) );
  AOI22D1BWP30P140LVT U152 ( .A1(n2), .A2(i_data_bus[125]), .B1(n1), .B2(
        i_data_bus[157]), .ZN(n125) );
  ND3D1BWP30P140LVT U153 ( .A1(n127), .A2(n126), .A3(n125), .ZN(N398) );
  AOI22D1BWP30P140LVT U154 ( .A1(n3), .A2(i_data_bus[220]), .B1(n214), .B2(
        i_data_bus[188]), .ZN(n128) );
  IOA21D1BWP30P140LVT U155 ( .A1(n216), .A2(i_data_bus[252]), .B(n128), .ZN(
        n129) );
  AOI21D1BWP30P140LVT U156 ( .A1(n152), .A2(i_data_bus[28]), .B(n129), .ZN(
        n132) );
  AOI22D1BWP30P140LVT U157 ( .A1(n220), .A2(i_data_bus[92]), .B1(n219), .B2(
        i_data_bus[60]), .ZN(n131) );
  AOI22D1BWP30P140LVT U158 ( .A1(n2), .A2(i_data_bus[124]), .B1(n1), .B2(
        i_data_bus[156]), .ZN(n130) );
  ND3D1BWP30P140LVT U159 ( .A1(n132), .A2(n131), .A3(n130), .ZN(N397) );
  AOI22D1BWP30P140LVT U160 ( .A1(n3), .A2(i_data_bus[219]), .B1(n214), .B2(
        i_data_bus[187]), .ZN(n133) );
  IOA21D1BWP30P140LVT U161 ( .A1(n216), .A2(i_data_bus[251]), .B(n133), .ZN(
        n134) );
  AOI21D1BWP30P140LVT U162 ( .A1(n152), .A2(i_data_bus[27]), .B(n134), .ZN(
        n137) );
  AOI22D1BWP30P140LVT U163 ( .A1(n220), .A2(i_data_bus[91]), .B1(n219), .B2(
        i_data_bus[59]), .ZN(n136) );
  AOI22D1BWP30P140LVT U164 ( .A1(n2), .A2(i_data_bus[123]), .B1(n1), .B2(
        i_data_bus[155]), .ZN(n135) );
  ND3D1BWP30P140LVT U165 ( .A1(n137), .A2(n136), .A3(n135), .ZN(N396) );
  AOI22D1BWP30P140LVT U166 ( .A1(n3), .A2(i_data_bus[218]), .B1(n214), .B2(
        i_data_bus[186]), .ZN(n138) );
  IOA21D1BWP30P140LVT U167 ( .A1(n216), .A2(i_data_bus[250]), .B(n138), .ZN(
        n139) );
  AOI21D1BWP30P140LVT U168 ( .A1(n152), .A2(i_data_bus[26]), .B(n139), .ZN(
        n142) );
  AOI22D1BWP30P140LVT U169 ( .A1(n220), .A2(i_data_bus[90]), .B1(n219), .B2(
        i_data_bus[58]), .ZN(n141) );
  AOI22D1BWP30P140LVT U170 ( .A1(n2), .A2(i_data_bus[122]), .B1(n1), .B2(
        i_data_bus[154]), .ZN(n140) );
  ND3D1BWP30P140LVT U171 ( .A1(n142), .A2(n141), .A3(n140), .ZN(N395) );
  AOI22D1BWP30P140LVT U172 ( .A1(n3), .A2(i_data_bus[217]), .B1(n214), .B2(
        i_data_bus[185]), .ZN(n143) );
  IOA21D1BWP30P140LVT U173 ( .A1(n216), .A2(i_data_bus[249]), .B(n143), .ZN(
        n144) );
  AOI21D1BWP30P140LVT U174 ( .A1(n152), .A2(i_data_bus[25]), .B(n144), .ZN(
        n149) );
  INVD2BWP30P140LVT U175 ( .I(n145), .ZN(n220) );
  AOI22D1BWP30P140LVT U176 ( .A1(n220), .A2(i_data_bus[89]), .B1(n219), .B2(
        i_data_bus[57]), .ZN(n148) );
  AOI22D1BWP30P140LVT U177 ( .A1(n2), .A2(i_data_bus[121]), .B1(n1), .B2(
        i_data_bus[153]), .ZN(n147) );
  ND3D1BWP30P140LVT U178 ( .A1(n149), .A2(n148), .A3(n147), .ZN(N394) );
  AOI22D1BWP30P140LVT U179 ( .A1(n3), .A2(i_data_bus[223]), .B1(n214), .B2(
        i_data_bus[191]), .ZN(n150) );
  IOA21D1BWP30P140LVT U180 ( .A1(n216), .A2(i_data_bus[255]), .B(n150), .ZN(
        n151) );
  AOI21D1BWP30P140LVT U181 ( .A1(n152), .A2(i_data_bus[31]), .B(n151), .ZN(
        n155) );
  AOI22D1BWP30P140LVT U182 ( .A1(n220), .A2(i_data_bus[95]), .B1(n219), .B2(
        i_data_bus[63]), .ZN(n154) );
  AOI22D1BWP30P140LVT U183 ( .A1(n2), .A2(i_data_bus[127]), .B1(n1), .B2(
        i_data_bus[159]), .ZN(n153) );
  ND3D1BWP30P140LVT U184 ( .A1(n155), .A2(n154), .A3(n153), .ZN(N400) );
  INVD2BWP30P140LVT U185 ( .I(n156), .ZN(n218) );
  AOI22D1BWP30P140LVT U186 ( .A1(n3), .A2(i_data_bus[210]), .B1(n214), .B2(
        i_data_bus[178]), .ZN(n157) );
  IOA21D1BWP30P140LVT U187 ( .A1(n216), .A2(i_data_bus[242]), .B(n157), .ZN(
        n158) );
  AOI21D1BWP30P140LVT U188 ( .A1(n218), .A2(i_data_bus[18]), .B(n158), .ZN(
        n161) );
  AOI22D1BWP30P140LVT U189 ( .A1(n220), .A2(i_data_bus[82]), .B1(n219), .B2(
        i_data_bus[50]), .ZN(n160) );
  AOI22D1BWP30P140LVT U190 ( .A1(n2), .A2(i_data_bus[114]), .B1(n1), .B2(
        i_data_bus[146]), .ZN(n159) );
  ND3D1BWP30P140LVT U191 ( .A1(n161), .A2(n160), .A3(n159), .ZN(N387) );
  AOI22D1BWP30P140LVT U192 ( .A1(n3), .A2(i_data_bus[209]), .B1(n214), .B2(
        i_data_bus[177]), .ZN(n162) );
  IOA21D1BWP30P140LVT U193 ( .A1(n216), .A2(i_data_bus[241]), .B(n162), .ZN(
        n163) );
  AOI21D1BWP30P140LVT U194 ( .A1(n218), .A2(i_data_bus[17]), .B(n163), .ZN(
        n166) );
  AOI22D1BWP30P140LVT U195 ( .A1(n220), .A2(i_data_bus[81]), .B1(n219), .B2(
        i_data_bus[49]), .ZN(n165) );
  AOI22D1BWP30P140LVT U196 ( .A1(n2), .A2(i_data_bus[113]), .B1(n1), .B2(
        i_data_bus[145]), .ZN(n164) );
  ND3D1BWP30P140LVT U197 ( .A1(n166), .A2(n165), .A3(n164), .ZN(N386) );
  AOI22D1BWP30P140LVT U198 ( .A1(n3), .A2(i_data_bus[208]), .B1(n214), .B2(
        i_data_bus[176]), .ZN(n167) );
  IOA21D1BWP30P140LVT U199 ( .A1(n216), .A2(i_data_bus[240]), .B(n167), .ZN(
        n168) );
  AOI21D1BWP30P140LVT U200 ( .A1(n218), .A2(i_data_bus[16]), .B(n168), .ZN(
        n171) );
  AOI22D1BWP30P140LVT U201 ( .A1(n220), .A2(i_data_bus[80]), .B1(n219), .B2(
        i_data_bus[48]), .ZN(n170) );
  AOI22D1BWP30P140LVT U202 ( .A1(n2), .A2(i_data_bus[112]), .B1(n1), .B2(
        i_data_bus[144]), .ZN(n169) );
  ND3D1BWP30P140LVT U203 ( .A1(n171), .A2(n170), .A3(n169), .ZN(N385) );
  AOI22D1BWP30P140LVT U204 ( .A1(n3), .A2(i_data_bus[207]), .B1(n214), .B2(
        i_data_bus[175]), .ZN(n172) );
  IOA21D1BWP30P140LVT U205 ( .A1(n216), .A2(i_data_bus[239]), .B(n172), .ZN(
        n173) );
  AOI21D1BWP30P140LVT U206 ( .A1(n218), .A2(i_data_bus[15]), .B(n173), .ZN(
        n176) );
  AOI22D1BWP30P140LVT U207 ( .A1(n220), .A2(i_data_bus[79]), .B1(n219), .B2(
        i_data_bus[47]), .ZN(n175) );
  AOI22D1BWP30P140LVT U208 ( .A1(n2), .A2(i_data_bus[111]), .B1(n1), .B2(
        i_data_bus[143]), .ZN(n174) );
  ND3D1BWP30P140LVT U209 ( .A1(n176), .A2(n175), .A3(n174), .ZN(N384) );
  AOI22D1BWP30P140LVT U210 ( .A1(n3), .A2(i_data_bus[206]), .B1(n214), .B2(
        i_data_bus[174]), .ZN(n177) );
  IOA21D1BWP30P140LVT U211 ( .A1(n216), .A2(i_data_bus[238]), .B(n177), .ZN(
        n178) );
  AOI21D1BWP30P140LVT U212 ( .A1(n218), .A2(i_data_bus[14]), .B(n178), .ZN(
        n181) );
  AOI22D1BWP30P140LVT U213 ( .A1(n220), .A2(i_data_bus[78]), .B1(n219), .B2(
        i_data_bus[46]), .ZN(n180) );
  AOI22D1BWP30P140LVT U214 ( .A1(n2), .A2(i_data_bus[110]), .B1(n1), .B2(
        i_data_bus[142]), .ZN(n179) );
  ND3D1BWP30P140LVT U215 ( .A1(n181), .A2(n180), .A3(n179), .ZN(N383) );
  INVD1BWP30P140LVT U216 ( .I(i_data_bus[173]), .ZN(n182) );
  MAOI22D1BWP30P140LVT U217 ( .A1(n3), .A2(i_data_bus[205]), .B1(n183), .B2(
        n182), .ZN(n184) );
  IOA21D1BWP30P140LVT U218 ( .A1(n216), .A2(i_data_bus[237]), .B(n184), .ZN(
        n185) );
  AOI21D1BWP30P140LVT U219 ( .A1(n218), .A2(i_data_bus[13]), .B(n185), .ZN(
        n188) );
  AOI22D1BWP30P140LVT U220 ( .A1(n220), .A2(i_data_bus[77]), .B1(n219), .B2(
        i_data_bus[45]), .ZN(n187) );
  AOI22D1BWP30P140LVT U221 ( .A1(n2), .A2(i_data_bus[109]), .B1(n1), .B2(
        i_data_bus[141]), .ZN(n186) );
  ND3D1BWP30P140LVT U222 ( .A1(n188), .A2(n187), .A3(n186), .ZN(N382) );
  AOI22D1BWP30P140LVT U223 ( .A1(n3), .A2(i_data_bus[216]), .B1(n214), .B2(
        i_data_bus[184]), .ZN(n189) );
  IOA21D1BWP30P140LVT U224 ( .A1(n216), .A2(i_data_bus[248]), .B(n189), .ZN(
        n190) );
  AOI21D1BWP30P140LVT U225 ( .A1(n218), .A2(i_data_bus[24]), .B(n190), .ZN(
        n193) );
  AOI22D1BWP30P140LVT U226 ( .A1(n220), .A2(i_data_bus[88]), .B1(n219), .B2(
        i_data_bus[56]), .ZN(n192) );
  AOI22D1BWP30P140LVT U227 ( .A1(n2), .A2(i_data_bus[120]), .B1(n1), .B2(
        i_data_bus[152]), .ZN(n191) );
  ND3D1BWP30P140LVT U228 ( .A1(n193), .A2(n192), .A3(n191), .ZN(N393) );
  AOI22D1BWP30P140LVT U229 ( .A1(n3), .A2(i_data_bus[215]), .B1(n214), .B2(
        i_data_bus[183]), .ZN(n194) );
  IOA21D1BWP30P140LVT U230 ( .A1(n216), .A2(i_data_bus[247]), .B(n194), .ZN(
        n195) );
  AOI21D1BWP30P140LVT U231 ( .A1(n218), .A2(i_data_bus[23]), .B(n195), .ZN(
        n198) );
  AOI22D1BWP30P140LVT U232 ( .A1(n220), .A2(i_data_bus[87]), .B1(n219), .B2(
        i_data_bus[55]), .ZN(n197) );
  AOI22D1BWP30P140LVT U233 ( .A1(n2), .A2(i_data_bus[119]), .B1(n1), .B2(
        i_data_bus[151]), .ZN(n196) );
  ND3D1BWP30P140LVT U234 ( .A1(n198), .A2(n197), .A3(n196), .ZN(N392) );
  AOI22D1BWP30P140LVT U235 ( .A1(n3), .A2(i_data_bus[214]), .B1(n214), .B2(
        i_data_bus[182]), .ZN(n199) );
  IOA21D1BWP30P140LVT U236 ( .A1(n216), .A2(i_data_bus[246]), .B(n199), .ZN(
        n200) );
  AOI21D1BWP30P140LVT U237 ( .A1(n218), .A2(i_data_bus[22]), .B(n200), .ZN(
        n203) );
  AOI22D1BWP30P140LVT U238 ( .A1(n220), .A2(i_data_bus[86]), .B1(n219), .B2(
        i_data_bus[54]), .ZN(n202) );
  AOI22D1BWP30P140LVT U239 ( .A1(n2), .A2(i_data_bus[118]), .B1(n1), .B2(
        i_data_bus[150]), .ZN(n201) );
  ND3D1BWP30P140LVT U240 ( .A1(n203), .A2(n202), .A3(n201), .ZN(N391) );
  AOI22D1BWP30P140LVT U241 ( .A1(n3), .A2(i_data_bus[213]), .B1(n214), .B2(
        i_data_bus[181]), .ZN(n204) );
  IOA21D1BWP30P140LVT U242 ( .A1(n216), .A2(i_data_bus[245]), .B(n204), .ZN(
        n205) );
  AOI21D1BWP30P140LVT U243 ( .A1(n218), .A2(i_data_bus[21]), .B(n205), .ZN(
        n208) );
  AOI22D1BWP30P140LVT U244 ( .A1(n220), .A2(i_data_bus[85]), .B1(n219), .B2(
        i_data_bus[53]), .ZN(n207) );
  AOI22D1BWP30P140LVT U245 ( .A1(n2), .A2(i_data_bus[117]), .B1(n1), .B2(
        i_data_bus[149]), .ZN(n206) );
  ND3D1BWP30P140LVT U246 ( .A1(n208), .A2(n207), .A3(n206), .ZN(N390) );
  AOI22D1BWP30P140LVT U247 ( .A1(n3), .A2(i_data_bus[212]), .B1(n214), .B2(
        i_data_bus[180]), .ZN(n209) );
  IOA21D1BWP30P140LVT U248 ( .A1(n216), .A2(i_data_bus[244]), .B(n209), .ZN(
        n210) );
  AOI21D1BWP30P140LVT U249 ( .A1(n218), .A2(i_data_bus[20]), .B(n210), .ZN(
        n213) );
  AOI22D1BWP30P140LVT U250 ( .A1(n220), .A2(i_data_bus[84]), .B1(n219), .B2(
        i_data_bus[52]), .ZN(n212) );
  AOI22D1BWP30P140LVT U251 ( .A1(n2), .A2(i_data_bus[116]), .B1(n1), .B2(
        i_data_bus[148]), .ZN(n211) );
  ND3D1BWP30P140LVT U252 ( .A1(n213), .A2(n212), .A3(n211), .ZN(N389) );
  AOI22D1BWP30P140LVT U253 ( .A1(n3), .A2(i_data_bus[211]), .B1(n214), .B2(
        i_data_bus[179]), .ZN(n215) );
  IOA21D1BWP30P140LVT U254 ( .A1(n216), .A2(i_data_bus[243]), .B(n215), .ZN(
        n217) );
  AOI21D1BWP30P140LVT U255 ( .A1(n218), .A2(i_data_bus[19]), .B(n217), .ZN(
        n223) );
  AOI22D1BWP30P140LVT U256 ( .A1(n220), .A2(i_data_bus[83]), .B1(n219), .B2(
        i_data_bus[51]), .ZN(n222) );
  AOI22D1BWP30P140LVT U257 ( .A1(n2), .A2(i_data_bus[115]), .B1(n1), .B2(
        i_data_bus[147]), .ZN(n221) );
  ND3D1BWP30P140LVT U258 ( .A1(n223), .A2(n222), .A3(n221), .ZN(N388) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_2 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  AOI21D1BWP30P140LVT U3 ( .A1(n220), .A2(i_data_bus[4]), .B(n88), .ZN(n91) );
  INVD3BWP30P140LVT U4 ( .I(n174), .ZN(n3) );
  INVD2BWP30P140LVT U5 ( .I(n172), .ZN(n163) );
  NR2D1BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n26) );
  INR4D2BWP30P140LVT U7 ( .A1(i_valid[6]), .B1(i_cmd[5]), .B2(i_cmd[7]), .B3(
        n18), .ZN(n19) );
  INVD4BWP30P140LVT U8 ( .I(n211), .ZN(n1) );
  INVD8BWP30P140LVT U9 ( .I(n226), .ZN(n2) );
  INVD2BWP30P140LVT U10 ( .I(n53), .ZN(n164) );
  ND2D1BWP30P140LVT U11 ( .A1(n11), .A2(n27), .ZN(n34) );
  ND2D1BWP30P140LVT U12 ( .A1(n42), .A2(n9), .ZN(n47) );
  ND2OPTIBD1BWP30P140LVT U13 ( .A1(n42), .A2(n41), .ZN(n53) );
  INVD1BWP30P140LVT U14 ( .I(n39), .ZN(n104) );
  INVD1BWP30P140LVT U15 ( .I(n104), .ZN(n165) );
  INVD1BWP30P140LVT U16 ( .I(n33), .ZN(n172) );
  INVD1BWP30P140LVT U17 ( .I(n104), .ZN(n231) );
  INVD2BWP30P140LVT U18 ( .I(n53), .ZN(n230) );
  INVD2BWP30P140LVT U19 ( .I(n172), .ZN(n229) );
  INR4D1BWP30P140LVT U20 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n21), .ZN(n23) );
  INVD2BWP30P140LVT U21 ( .I(n47), .ZN(n220) );
  INVD1BWP30P140LVT U22 ( .I(n29), .ZN(n174) );
  OR2D1BWP30P140LVT U23 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n30) );
  NR2OPTPAD1BWP30P140LVT U24 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .ZN(n6) );
  INR2D1BWP30P140LVT U25 ( .A1(i_en), .B1(rst), .ZN(n4) );
  INR2D1BWP30P140LVT U26 ( .A1(n4), .B1(i_cmd[6]), .ZN(n5) );
  ND2OPTIBD2BWP30P140LVT U27 ( .A1(n6), .A2(n5), .ZN(n25) );
  NR3D0P7BWP30P140LVT U28 ( .A1(n30), .A2(n25), .A3(i_cmd[1]), .ZN(n42) );
  INR2D1BWP30P140LVT U29 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n7) );
  INVD1BWP30P140LVT U30 ( .I(n7), .ZN(n8) );
  INR2D1BWP30P140LVT U31 ( .A1(i_cmd[0]), .B1(n8), .ZN(n9) );
  ND2D1BWP30P140LVT U32 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n10) );
  NR3D0P7BWP30P140LVT U33 ( .A1(n10), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n16)
         );
  INVD1BWP30P140LVT U34 ( .I(i_cmd[2]), .ZN(n11) );
  INVD2BWP30P140LVT U35 ( .I(i_cmd[1]), .ZN(n27) );
  NR2OPTPAD1BWP30P140LVT U36 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n14) );
  INR2D1BWP30P140LVT U37 ( .A1(i_en), .B1(rst), .ZN(n12) );
  INR2D1BWP30P140LVT U38 ( .A1(n12), .B1(i_cmd[3]), .ZN(n13) );
  ND2OPTIBD1BWP30P140LVT U39 ( .A1(n14), .A2(n13), .ZN(n15) );
  OR2D4BWP30P140LVT U40 ( .A1(n34), .A2(n15), .Z(n22) );
  INR2D2BWP30P140LVT U41 ( .A1(n16), .B1(n22), .ZN(n17) );
  INVD1BWP30P140LVT U42 ( .I(i_cmd[6]), .ZN(n18) );
  INR2D1BWP30P140LVT U43 ( .A1(n19), .B1(n22), .ZN(n20) );
  INVD3BWP30P140LVT U44 ( .I(n20), .ZN(n226) );
  INVD1BWP30P140LVT U45 ( .I(i_cmd[5]), .ZN(n21) );
  INR2D2BWP30P140LVT U46 ( .A1(n23), .B1(n22), .ZN(n24) );
  INVD2BWP30P140LVT U47 ( .I(n24), .ZN(n211) );
  NR4D0BWP30P140LVT U48 ( .A1(n220), .A2(n17), .A3(n2), .A4(n1), .ZN(n45) );
  INR2D2BWP30P140LVT U49 ( .A1(n26), .B1(n25), .ZN(n38) );
  INVD1BWP30P140LVT U50 ( .I(i_cmd[3]), .ZN(n35) );
  ND4D1BWP30P140LVT U51 ( .A1(n27), .A2(n35), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n28) );
  INR2D1BWP30P140LVT U52 ( .A1(n38), .B1(n28), .ZN(n29) );
  INVD1BWP30P140LVT U53 ( .I(n30), .ZN(n31) );
  ND3D1BWP30P140LVT U54 ( .A1(n31), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n32)
         );
  INR2D1BWP30P140LVT U55 ( .A1(n38), .B1(n32), .ZN(n33) );
  NR2D1BWP30P140LVT U56 ( .A1(n29), .A2(n229), .ZN(n44) );
  INVD1BWP30P140LVT U57 ( .I(n34), .ZN(n36) );
  ND3D1BWP30P140LVT U58 ( .A1(n36), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n37)
         );
  INR2D1BWP30P140LVT U59 ( .A1(n38), .B1(n37), .ZN(n39) );
  INVD1BWP30P140LVT U60 ( .I(n104), .ZN(n221) );
  IND3D1BWP30P140LVT U61 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n40) );
  INVD1BWP30P140LVT U62 ( .I(n40), .ZN(n41) );
  NR2D1BWP30P140LVT U63 ( .A1(n221), .A2(n230), .ZN(n43) );
  ND3D1BWP30P140LVT U64 ( .A1(n45), .A2(n44), .A3(n43), .ZN(N402) );
  INVD1BWP30P140LVT U65 ( .I(n17), .ZN(n52) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[224]), .ZN(n51) );
  INVD1BWP30P140LVT U67 ( .I(i_data_bus[192]), .ZN(n46) );
  MAOI22D1BWP30P140LVT U68 ( .A1(n1), .A2(i_data_bus[160]), .B1(n226), .B2(n46), .ZN(n50) );
  INR2D1BWP30P140LVT U69 ( .A1(i_data_bus[0]), .B1(n47), .ZN(n48) );
  INVD1BWP30P140LVT U70 ( .I(n48), .ZN(n49) );
  OA211D1BWP30P140LVT U71 ( .A1(n52), .A2(n51), .B(n50), .C(n49), .Z(n56) );
  AOI22D1BWP30P140LVT U72 ( .A1(n3), .A2(i_data_bus[64]), .B1(n163), .B2(
        i_data_bus[32]), .ZN(n55) );
  AOI22D1BWP30P140LVT U73 ( .A1(n165), .A2(i_data_bus[96]), .B1(n164), .B2(
        i_data_bus[128]), .ZN(n54) );
  ND3D1BWP30P140LVT U74 ( .A1(n56), .A2(n55), .A3(n54), .ZN(N369) );
  AOI22D1BWP30P140LVT U75 ( .A1(n2), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n57) );
  IOA21D1BWP30P140LVT U76 ( .A1(n17), .A2(i_data_bus[233]), .B(n57), .ZN(n58)
         );
  AOI21D1BWP30P140LVT U77 ( .A1(n220), .A2(i_data_bus[9]), .B(n58), .ZN(n61)
         );
  AOI22D1BWP30P140LVT U78 ( .A1(n3), .A2(i_data_bus[73]), .B1(n163), .B2(
        i_data_bus[41]), .ZN(n60) );
  AOI22D1BWP30P140LVT U79 ( .A1(n165), .A2(i_data_bus[105]), .B1(n164), .B2(
        i_data_bus[137]), .ZN(n59) );
  ND3D1BWP30P140LVT U80 ( .A1(n61), .A2(n60), .A3(n59), .ZN(N378) );
  AOI22D1BWP30P140LVT U81 ( .A1(n2), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n62) );
  IOA21D1BWP30P140LVT U82 ( .A1(n17), .A2(i_data_bus[235]), .B(n62), .ZN(n63)
         );
  AOI21D1BWP30P140LVT U83 ( .A1(n220), .A2(i_data_bus[11]), .B(n63), .ZN(n66)
         );
  AOI22D1BWP30P140LVT U84 ( .A1(n3), .A2(i_data_bus[75]), .B1(n163), .B2(
        i_data_bus[43]), .ZN(n65) );
  AOI22D1BWP30P140LVT U85 ( .A1(n165), .A2(i_data_bus[107]), .B1(n164), .B2(
        i_data_bus[139]), .ZN(n64) );
  ND3D1BWP30P140LVT U86 ( .A1(n66), .A2(n65), .A3(n64), .ZN(N380) );
  AOI22D1BWP30P140LVT U87 ( .A1(n2), .A2(i_data_bus[199]), .B1(n1), .B2(
        i_data_bus[167]), .ZN(n67) );
  IOA21D1BWP30P140LVT U88 ( .A1(n17), .A2(i_data_bus[231]), .B(n67), .ZN(n68)
         );
  AOI21D1BWP30P140LVT U89 ( .A1(n220), .A2(i_data_bus[7]), .B(n68), .ZN(n71)
         );
  AOI22D1BWP30P140LVT U90 ( .A1(n3), .A2(i_data_bus[71]), .B1(n163), .B2(
        i_data_bus[39]), .ZN(n70) );
  AOI22D1BWP30P140LVT U91 ( .A1(n165), .A2(i_data_bus[103]), .B1(n164), .B2(
        i_data_bus[135]), .ZN(n69) );
  ND3D1BWP30P140LVT U92 ( .A1(n71), .A2(n70), .A3(n69), .ZN(N376) );
  AOI22D1BWP30P140LVT U93 ( .A1(n2), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n72) );
  IOA21D1BWP30P140LVT U94 ( .A1(n17), .A2(i_data_bus[229]), .B(n72), .ZN(n73)
         );
  AOI21D1BWP30P140LVT U95 ( .A1(n220), .A2(i_data_bus[5]), .B(n73), .ZN(n76)
         );
  AOI22D1BWP30P140LVT U96 ( .A1(n3), .A2(i_data_bus[69]), .B1(n163), .B2(
        i_data_bus[37]), .ZN(n75) );
  AOI22D1BWP30P140LVT U97 ( .A1(n165), .A2(i_data_bus[101]), .B1(n164), .B2(
        i_data_bus[133]), .ZN(n74) );
  ND3D1BWP30P140LVT U98 ( .A1(n76), .A2(n75), .A3(n74), .ZN(N374) );
  AOI22D1BWP30P140LVT U99 ( .A1(n2), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n77) );
  IOA21D1BWP30P140LVT U100 ( .A1(n17), .A2(i_data_bus[230]), .B(n77), .ZN(n78)
         );
  AOI21D1BWP30P140LVT U101 ( .A1(n220), .A2(i_data_bus[6]), .B(n78), .ZN(n81)
         );
  AOI22D1BWP30P140LVT U102 ( .A1(n3), .A2(i_data_bus[70]), .B1(n163), .B2(
        i_data_bus[38]), .ZN(n80) );
  AOI22D1BWP30P140LVT U103 ( .A1(n165), .A2(i_data_bus[102]), .B1(n164), .B2(
        i_data_bus[134]), .ZN(n79) );
  ND3D1BWP30P140LVT U104 ( .A1(n81), .A2(n80), .A3(n79), .ZN(N375) );
  AOI22D1BWP30P140LVT U105 ( .A1(n2), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n82) );
  IOA21D1BWP30P140LVT U106 ( .A1(n17), .A2(i_data_bus[232]), .B(n82), .ZN(n83)
         );
  AOI21D1BWP30P140LVT U107 ( .A1(n220), .A2(i_data_bus[8]), .B(n83), .ZN(n86)
         );
  AOI22D1BWP30P140LVT U108 ( .A1(n3), .A2(i_data_bus[72]), .B1(n163), .B2(
        i_data_bus[40]), .ZN(n85) );
  AOI22D1BWP30P140LVT U109 ( .A1(n165), .A2(i_data_bus[104]), .B1(n164), .B2(
        i_data_bus[136]), .ZN(n84) );
  ND3D1BWP30P140LVT U110 ( .A1(n86), .A2(n85), .A3(n84), .ZN(N377) );
  AOI22D1BWP30P140LVT U111 ( .A1(n2), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n87) );
  IOA21D1BWP30P140LVT U112 ( .A1(n17), .A2(i_data_bus[228]), .B(n87), .ZN(n88)
         );
  AOI22D1BWP30P140LVT U113 ( .A1(n3), .A2(i_data_bus[68]), .B1(n163), .B2(
        i_data_bus[36]), .ZN(n90) );
  AOI22D1BWP30P140LVT U114 ( .A1(n165), .A2(i_data_bus[100]), .B1(n164), .B2(
        i_data_bus[132]), .ZN(n89) );
  ND3D1BWP30P140LVT U115 ( .A1(n91), .A2(n90), .A3(n89), .ZN(N373) );
  AOI22D1BWP30P140LVT U116 ( .A1(n2), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n92) );
  IOA21D1BWP30P140LVT U117 ( .A1(n17), .A2(i_data_bus[234]), .B(n92), .ZN(n93)
         );
  AOI21D1BWP30P140LVT U118 ( .A1(n220), .A2(i_data_bus[10]), .B(n93), .ZN(n96)
         );
  AOI22D1BWP30P140LVT U119 ( .A1(n3), .A2(i_data_bus[74]), .B1(n163), .B2(
        i_data_bus[42]), .ZN(n95) );
  AOI22D1BWP30P140LVT U120 ( .A1(n165), .A2(i_data_bus[106]), .B1(n164), .B2(
        i_data_bus[138]), .ZN(n94) );
  ND3D1BWP30P140LVT U121 ( .A1(n96), .A2(n95), .A3(n94), .ZN(N379) );
  AOI22D1BWP30P140LVT U122 ( .A1(n2), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n97) );
  IOA21D1BWP30P140LVT U123 ( .A1(n17), .A2(i_data_bus[236]), .B(n97), .ZN(n98)
         );
  AOI21D1BWP30P140LVT U124 ( .A1(n220), .A2(i_data_bus[12]), .B(n98), .ZN(n101) );
  AOI22D1BWP30P140LVT U125 ( .A1(n3), .A2(i_data_bus[76]), .B1(n163), .B2(
        i_data_bus[44]), .ZN(n100) );
  AOI22D1BWP30P140LVT U126 ( .A1(n165), .A2(i_data_bus[108]), .B1(n164), .B2(
        i_data_bus[140]), .ZN(n99) );
  ND3D1BWP30P140LVT U127 ( .A1(n101), .A2(n100), .A3(n99), .ZN(N381) );
  AOI22D1BWP30P140LVT U128 ( .A1(n2), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n102) );
  IOA21D1BWP30P140LVT U129 ( .A1(n17), .A2(i_data_bus[245]), .B(n102), .ZN(
        n103) );
  AOI21D1BWP30P140LVT U130 ( .A1(n220), .A2(i_data_bus[21]), .B(n103), .ZN(
        n107) );
  AOI22D1BWP30P140LVT U131 ( .A1(n3), .A2(i_data_bus[85]), .B1(n229), .B2(
        i_data_bus[53]), .ZN(n106) );
  AOI22D1BWP30P140LVT U132 ( .A1(n231), .A2(i_data_bus[117]), .B1(n230), .B2(
        i_data_bus[149]), .ZN(n105) );
  ND3D1BWP30P140LVT U133 ( .A1(n107), .A2(n106), .A3(n105), .ZN(N390) );
  AOI22D1BWP30P140LVT U134 ( .A1(n2), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n108) );
  IOA21D1BWP30P140LVT U135 ( .A1(n17), .A2(i_data_bus[247]), .B(n108), .ZN(
        n109) );
  AOI21D1BWP30P140LVT U136 ( .A1(n220), .A2(i_data_bus[23]), .B(n109), .ZN(
        n112) );
  AOI22D1BWP30P140LVT U137 ( .A1(n3), .A2(i_data_bus[87]), .B1(n229), .B2(
        i_data_bus[55]), .ZN(n111) );
  AOI22D1BWP30P140LVT U138 ( .A1(n231), .A2(i_data_bus[119]), .B1(n230), .B2(
        i_data_bus[151]), .ZN(n110) );
  ND3D1BWP30P140LVT U139 ( .A1(n112), .A2(n111), .A3(n110), .ZN(N392) );
  AOI22D1BWP30P140LVT U140 ( .A1(n2), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n113) );
  IOA21D1BWP30P140LVT U141 ( .A1(n17), .A2(i_data_bus[242]), .B(n113), .ZN(
        n114) );
  AOI21D1BWP30P140LVT U142 ( .A1(n220), .A2(i_data_bus[18]), .B(n114), .ZN(
        n117) );
  AOI22D1BWP30P140LVT U143 ( .A1(n3), .A2(i_data_bus[82]), .B1(n229), .B2(
        i_data_bus[50]), .ZN(n116) );
  AOI22D1BWP30P140LVT U144 ( .A1(n231), .A2(i_data_bus[114]), .B1(n230), .B2(
        i_data_bus[146]), .ZN(n115) );
  ND3D1BWP30P140LVT U145 ( .A1(n117), .A2(n116), .A3(n115), .ZN(N387) );
  AOI22D1BWP30P140LVT U146 ( .A1(n2), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n118) );
  IOA21D1BWP30P140LVT U147 ( .A1(n17), .A2(i_data_bus[243]), .B(n118), .ZN(
        n119) );
  AOI21D1BWP30P140LVT U148 ( .A1(n220), .A2(i_data_bus[19]), .B(n119), .ZN(
        n122) );
  AOI22D1BWP30P140LVT U149 ( .A1(n3), .A2(i_data_bus[83]), .B1(n229), .B2(
        i_data_bus[51]), .ZN(n121) );
  AOI22D1BWP30P140LVT U150 ( .A1(n231), .A2(i_data_bus[115]), .B1(n230), .B2(
        i_data_bus[147]), .ZN(n120) );
  ND3D1BWP30P140LVT U151 ( .A1(n122), .A2(n121), .A3(n120), .ZN(N388) );
  AOI22D1BWP30P140LVT U152 ( .A1(n2), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n123) );
  IOA21D1BWP30P140LVT U153 ( .A1(n17), .A2(i_data_bus[244]), .B(n123), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U154 ( .A1(n220), .A2(i_data_bus[20]), .B(n124), .ZN(
        n127) );
  AOI22D1BWP30P140LVT U155 ( .A1(n3), .A2(i_data_bus[84]), .B1(n229), .B2(
        i_data_bus[52]), .ZN(n126) );
  AOI22D1BWP30P140LVT U156 ( .A1(n231), .A2(i_data_bus[116]), .B1(n230), .B2(
        i_data_bus[148]), .ZN(n125) );
  ND3D1BWP30P140LVT U157 ( .A1(n127), .A2(n126), .A3(n125), .ZN(N389) );
  AOI22D1BWP30P140LVT U158 ( .A1(n2), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n128) );
  IOA21D1BWP30P140LVT U159 ( .A1(n17), .A2(i_data_bus[241]), .B(n128), .ZN(
        n129) );
  AOI21D1BWP30P140LVT U160 ( .A1(n220), .A2(i_data_bus[17]), .B(n129), .ZN(
        n132) );
  AOI22D1BWP30P140LVT U161 ( .A1(n3), .A2(i_data_bus[81]), .B1(n229), .B2(
        i_data_bus[49]), .ZN(n131) );
  AOI22D1BWP30P140LVT U162 ( .A1(n231), .A2(i_data_bus[113]), .B1(n230), .B2(
        i_data_bus[145]), .ZN(n130) );
  ND3D1BWP30P140LVT U163 ( .A1(n132), .A2(n131), .A3(n130), .ZN(N386) );
  AOI22D1BWP30P140LVT U164 ( .A1(n2), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n133) );
  IOA21D1BWP30P140LVT U165 ( .A1(n17), .A2(i_data_bus[248]), .B(n133), .ZN(
        n134) );
  AOI21D1BWP30P140LVT U166 ( .A1(n220), .A2(i_data_bus[24]), .B(n134), .ZN(
        n137) );
  AOI22D1BWP30P140LVT U167 ( .A1(n3), .A2(i_data_bus[88]), .B1(n229), .B2(
        i_data_bus[56]), .ZN(n136) );
  AOI22D1BWP30P140LVT U168 ( .A1(n231), .A2(i_data_bus[120]), .B1(n230), .B2(
        i_data_bus[152]), .ZN(n135) );
  ND3D1BWP30P140LVT U169 ( .A1(n137), .A2(n136), .A3(n135), .ZN(N393) );
  AOI22D1BWP30P140LVT U170 ( .A1(n2), .A2(i_data_bus[206]), .B1(n1), .B2(
        i_data_bus[174]), .ZN(n138) );
  IOA21D1BWP30P140LVT U171 ( .A1(n17), .A2(i_data_bus[238]), .B(n138), .ZN(
        n139) );
  AOI21D1BWP30P140LVT U172 ( .A1(n220), .A2(i_data_bus[14]), .B(n139), .ZN(
        n142) );
  AOI22D1BWP30P140LVT U173 ( .A1(n3), .A2(i_data_bus[78]), .B1(n229), .B2(
        i_data_bus[46]), .ZN(n141) );
  AOI22D1BWP30P140LVT U174 ( .A1(n231), .A2(i_data_bus[110]), .B1(n230), .B2(
        i_data_bus[142]), .ZN(n140) );
  ND3D1BWP30P140LVT U175 ( .A1(n142), .A2(n141), .A3(n140), .ZN(N383) );
  AOI22D1BWP30P140LVT U176 ( .A1(n2), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n143) );
  IOA21D1BWP30P140LVT U177 ( .A1(n17), .A2(i_data_bus[246]), .B(n143), .ZN(
        n144) );
  AOI21D1BWP30P140LVT U178 ( .A1(n220), .A2(i_data_bus[22]), .B(n144), .ZN(
        n147) );
  AOI22D1BWP30P140LVT U179 ( .A1(n3), .A2(i_data_bus[86]), .B1(n229), .B2(
        i_data_bus[54]), .ZN(n146) );
  AOI22D1BWP30P140LVT U180 ( .A1(n231), .A2(i_data_bus[118]), .B1(n230), .B2(
        i_data_bus[150]), .ZN(n145) );
  ND3D1BWP30P140LVT U181 ( .A1(n147), .A2(n146), .A3(n145), .ZN(N391) );
  INVD1BWP30P140LVT U182 ( .I(i_data_bus[195]), .ZN(n148) );
  MAOI22D1BWP30P140LVT U183 ( .A1(n1), .A2(i_data_bus[163]), .B1(n226), .B2(
        n148), .ZN(n149) );
  IOA21D1BWP30P140LVT U184 ( .A1(n17), .A2(i_data_bus[227]), .B(n149), .ZN(
        n150) );
  AOI21D1BWP30P140LVT U185 ( .A1(n220), .A2(i_data_bus[3]), .B(n150), .ZN(n153) );
  AOI22D1BWP30P140LVT U186 ( .A1(n3), .A2(i_data_bus[67]), .B1(n163), .B2(
        i_data_bus[35]), .ZN(n152) );
  AOI22D1BWP30P140LVT U187 ( .A1(n165), .A2(i_data_bus[99]), .B1(n164), .B2(
        i_data_bus[131]), .ZN(n151) );
  ND3D1BWP30P140LVT U188 ( .A1(n153), .A2(n152), .A3(n151), .ZN(N372) );
  INVD1BWP30P140LVT U189 ( .I(i_data_bus[193]), .ZN(n154) );
  MAOI22D1BWP30P140LVT U190 ( .A1(n1), .A2(i_data_bus[161]), .B1(n226), .B2(
        n154), .ZN(n155) );
  IOA21D1BWP30P140LVT U191 ( .A1(n17), .A2(i_data_bus[225]), .B(n155), .ZN(
        n156) );
  AOI21D1BWP30P140LVT U192 ( .A1(n220), .A2(i_data_bus[1]), .B(n156), .ZN(n159) );
  AOI22D1BWP30P140LVT U193 ( .A1(n3), .A2(i_data_bus[65]), .B1(n163), .B2(
        i_data_bus[33]), .ZN(n158) );
  AOI22D1BWP30P140LVT U194 ( .A1(n165), .A2(i_data_bus[97]), .B1(n164), .B2(
        i_data_bus[129]), .ZN(n157) );
  ND3D1BWP30P140LVT U195 ( .A1(n159), .A2(n158), .A3(n157), .ZN(N370) );
  INVD1BWP30P140LVT U196 ( .I(i_data_bus[194]), .ZN(n160) );
  MAOI22D1BWP30P140LVT U197 ( .A1(n1), .A2(i_data_bus[162]), .B1(n226), .B2(
        n160), .ZN(n161) );
  IOA21D1BWP30P140LVT U198 ( .A1(n17), .A2(i_data_bus[226]), .B(n161), .ZN(
        n162) );
  AOI21D1BWP30P140LVT U199 ( .A1(n220), .A2(i_data_bus[2]), .B(n162), .ZN(n168) );
  AOI22D1BWP30P140LVT U200 ( .A1(n3), .A2(i_data_bus[66]), .B1(n163), .B2(
        i_data_bus[34]), .ZN(n167) );
  AOI22D1BWP30P140LVT U201 ( .A1(n165), .A2(i_data_bus[98]), .B1(n164), .B2(
        i_data_bus[130]), .ZN(n166) );
  ND3D1BWP30P140LVT U202 ( .A1(n168), .A2(n167), .A3(n166), .ZN(N371) );
  AOI22D1BWP30P140LVT U203 ( .A1(n2), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n169) );
  IOA21D1BWP30P140LVT U204 ( .A1(n17), .A2(i_data_bus[239]), .B(n169), .ZN(
        n170) );
  AOI21D1BWP30P140LVT U205 ( .A1(n220), .A2(i_data_bus[15]), .B(n170), .ZN(
        n177) );
  INVD1BWP30P140LVT U206 ( .I(i_data_bus[79]), .ZN(n173) );
  INVD1BWP30P140LVT U207 ( .I(i_data_bus[47]), .ZN(n171) );
  OA22D1BWP30P140LVT U208 ( .A1(n174), .A2(n173), .B1(n172), .B2(n171), .Z(
        n176) );
  AOI22D1BWP30P140LVT U209 ( .A1(n231), .A2(i_data_bus[111]), .B1(n230), .B2(
        i_data_bus[143]), .ZN(n175) );
  ND3D1BWP30P140LVT U210 ( .A1(n177), .A2(n176), .A3(n175), .ZN(N384) );
  AOI22D1BWP30P140LVT U211 ( .A1(n2), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n178) );
  IOA21D1BWP30P140LVT U212 ( .A1(n17), .A2(i_data_bus[249]), .B(n178), .ZN(
        n179) );
  AOI21D1BWP30P140LVT U213 ( .A1(n220), .A2(i_data_bus[25]), .B(n179), .ZN(
        n182) );
  AOI22D1BWP30P140LVT U214 ( .A1(n3), .A2(i_data_bus[89]), .B1(n229), .B2(
        i_data_bus[57]), .ZN(n181) );
  AOI22D1BWP30P140LVT U215 ( .A1(n231), .A2(i_data_bus[121]), .B1(n230), .B2(
        i_data_bus[153]), .ZN(n180) );
  ND3D1BWP30P140LVT U216 ( .A1(n182), .A2(n181), .A3(n180), .ZN(N394) );
  AOI22D1BWP30P140LVT U217 ( .A1(n2), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n183) );
  IOA21D1BWP30P140LVT U218 ( .A1(n17), .A2(i_data_bus[251]), .B(n183), .ZN(
        n184) );
  AOI21D1BWP30P140LVT U219 ( .A1(n220), .A2(i_data_bus[27]), .B(n184), .ZN(
        n187) );
  AOI22D1BWP30P140LVT U220 ( .A1(n3), .A2(i_data_bus[91]), .B1(n229), .B2(
        i_data_bus[59]), .ZN(n186) );
  AOI22D1BWP30P140LVT U221 ( .A1(n221), .A2(i_data_bus[123]), .B1(n230), .B2(
        i_data_bus[155]), .ZN(n185) );
  ND3D1BWP30P140LVT U222 ( .A1(n187), .A2(n186), .A3(n185), .ZN(N396) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[221]), .ZN(n188) );
  MAOI22D1BWP30P140LVT U224 ( .A1(n1), .A2(i_data_bus[189]), .B1(n226), .B2(
        n188), .ZN(n189) );
  IOA21D1BWP30P140LVT U225 ( .A1(n17), .A2(i_data_bus[253]), .B(n189), .ZN(
        n190) );
  AOI21D1BWP30P140LVT U226 ( .A1(n220), .A2(i_data_bus[29]), .B(n190), .ZN(
        n193) );
  AOI22D1BWP30P140LVT U227 ( .A1(n3), .A2(i_data_bus[93]), .B1(n229), .B2(
        i_data_bus[61]), .ZN(n192) );
  AOI22D1BWP30P140LVT U228 ( .A1(n221), .A2(i_data_bus[125]), .B1(n230), .B2(
        i_data_bus[157]), .ZN(n191) );
  ND3D1BWP30P140LVT U229 ( .A1(n193), .A2(n192), .A3(n191), .ZN(N398) );
  AOI22D1BWP30P140LVT U230 ( .A1(n2), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n194) );
  IOA21D1BWP30P140LVT U231 ( .A1(n17), .A2(i_data_bus[250]), .B(n194), .ZN(
        n195) );
  AOI21D1BWP30P140LVT U232 ( .A1(n220), .A2(i_data_bus[26]), .B(n195), .ZN(
        n198) );
  AOI22D1BWP30P140LVT U233 ( .A1(n3), .A2(i_data_bus[90]), .B1(n229), .B2(
        i_data_bus[58]), .ZN(n197) );
  AOI22D1BWP30P140LVT U234 ( .A1(n221), .A2(i_data_bus[122]), .B1(n230), .B2(
        i_data_bus[154]), .ZN(n196) );
  ND3D1BWP30P140LVT U235 ( .A1(n198), .A2(n197), .A3(n196), .ZN(N395) );
  INVD1BWP30P140LVT U236 ( .I(i_data_bus[223]), .ZN(n199) );
  MAOI22D1BWP30P140LVT U237 ( .A1(n1), .A2(i_data_bus[191]), .B1(n226), .B2(
        n199), .ZN(n200) );
  IOA21D1BWP30P140LVT U238 ( .A1(n17), .A2(i_data_bus[255]), .B(n200), .ZN(
        n201) );
  AOI21D1BWP30P140LVT U239 ( .A1(n220), .A2(i_data_bus[31]), .B(n201), .ZN(
        n204) );
  AOI22D1BWP30P140LVT U240 ( .A1(n3), .A2(i_data_bus[95]), .B1(n229), .B2(
        i_data_bus[63]), .ZN(n203) );
  AOI22D1BWP30P140LVT U241 ( .A1(n221), .A2(i_data_bus[127]), .B1(n230), .B2(
        i_data_bus[159]), .ZN(n202) );
  ND3D1BWP30P140LVT U242 ( .A1(n204), .A2(n203), .A3(n202), .ZN(N400) );
  AOI22D1BWP30P140LVT U243 ( .A1(n2), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n205) );
  IOA21D1BWP30P140LVT U244 ( .A1(n17), .A2(i_data_bus[252]), .B(n205), .ZN(
        n206) );
  AOI21D1BWP30P140LVT U245 ( .A1(n220), .A2(i_data_bus[28]), .B(n206), .ZN(
        n209) );
  AOI22D1BWP30P140LVT U246 ( .A1(n3), .A2(i_data_bus[92]), .B1(n229), .B2(
        i_data_bus[60]), .ZN(n208) );
  AOI22D1BWP30P140LVT U247 ( .A1(n221), .A2(i_data_bus[124]), .B1(n230), .B2(
        i_data_bus[156]), .ZN(n207) );
  ND3D1BWP30P140LVT U248 ( .A1(n209), .A2(n208), .A3(n207), .ZN(N397) );
  INVD1BWP30P140LVT U249 ( .I(i_data_bus[173]), .ZN(n210) );
  MAOI22D1BWP30P140LVT U250 ( .A1(n2), .A2(i_data_bus[205]), .B1(n211), .B2(
        n210), .ZN(n212) );
  IOA21D1BWP30P140LVT U251 ( .A1(n17), .A2(i_data_bus[237]), .B(n212), .ZN(
        n213) );
  AOI21D1BWP30P140LVT U252 ( .A1(n220), .A2(i_data_bus[13]), .B(n213), .ZN(
        n216) );
  AOI22D1BWP30P140LVT U253 ( .A1(n3), .A2(i_data_bus[77]), .B1(n229), .B2(
        i_data_bus[45]), .ZN(n215) );
  AOI22D1BWP30P140LVT U254 ( .A1(n231), .A2(i_data_bus[109]), .B1(n230), .B2(
        i_data_bus[141]), .ZN(n214) );
  ND3D1BWP30P140LVT U255 ( .A1(n216), .A2(n215), .A3(n214), .ZN(N382) );
  INVD1BWP30P140LVT U256 ( .I(i_data_bus[222]), .ZN(n217) );
  MAOI22D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[190]), .B1(n226), .B2(
        n217), .ZN(n218) );
  IOA21D1BWP30P140LVT U258 ( .A1(n17), .A2(i_data_bus[254]), .B(n218), .ZN(
        n219) );
  AOI21D1BWP30P140LVT U259 ( .A1(n220), .A2(i_data_bus[30]), .B(n219), .ZN(
        n224) );
  AOI22D1BWP30P140LVT U260 ( .A1(n29), .A2(i_data_bus[94]), .B1(n229), .B2(
        i_data_bus[62]), .ZN(n223) );
  AOI22D1BWP30P140LVT U261 ( .A1(n221), .A2(i_data_bus[126]), .B1(n230), .B2(
        i_data_bus[158]), .ZN(n222) );
  ND3D1BWP30P140LVT U262 ( .A1(n224), .A2(n223), .A3(n222), .ZN(N399) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[208]), .ZN(n225) );
  MAOI22D1BWP30P140LVT U264 ( .A1(n1), .A2(i_data_bus[176]), .B1(n226), .B2(
        n225), .ZN(n227) );
  IOA21D1BWP30P140LVT U265 ( .A1(n17), .A2(i_data_bus[240]), .B(n227), .ZN(
        n228) );
  AOI21D1BWP30P140LVT U266 ( .A1(n220), .A2(i_data_bus[16]), .B(n228), .ZN(
        n234) );
  AOI22D1BWP30P140LVT U267 ( .A1(n3), .A2(i_data_bus[80]), .B1(n229), .B2(
        i_data_bus[48]), .ZN(n233) );
  AOI22D1BWP30P140LVT U268 ( .A1(n231), .A2(i_data_bus[112]), .B1(n230), .B2(
        i_data_bus[144]), .ZN(n232) );
  ND3D1BWP30P140LVT U269 ( .A1(n234), .A2(n233), .A3(n232), .ZN(N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_3 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  AOI21D1BWP30P140LVT U3 ( .A1(n205), .A2(i_data_bus[6]), .B(n94), .ZN(n97) );
  INVD2BWP30P140LVT U4 ( .I(n216), .ZN(n206) );
  INVD6BWP30P140LVT U5 ( .I(n164), .ZN(n2) );
  NR2D1BWP30P140LVT U6 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n22) );
  INVD1BWP30P140LVT U7 ( .I(n29), .ZN(n216) );
  AOI21D1BWP30P140LVT U8 ( .A1(n205), .A2(i_data_bus[5]), .B(n99), .ZN(n102)
         );
  INVD4BWP30P140LVT U9 ( .I(n223), .ZN(n1) );
  IND2D2BWP30P140LVT U10 ( .A1(n30), .B1(n13), .ZN(n20) );
  INR2D2BWP30P140LVT U11 ( .A1(n22), .B1(n21), .ZN(n34) );
  ND2OPTIBD2BWP30P140LVT U12 ( .A1(n6), .A2(n5), .ZN(n21) );
  NR2D1BWP30P140LVT U13 ( .A1(i_cmd[6]), .A2(i_cmd[7]), .ZN(n18) );
  ND2D1BWP30P140LVT U14 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n9) );
  INR4D1BWP30P140LVT U15 ( .A1(i_valid[6]), .B1(i_cmd[5]), .B2(i_cmd[7]), .B3(
        n15), .ZN(n16) );
  INVD2BWP30P140LVT U16 ( .I(n49), .ZN(n208) );
  IND3D2BWP30P140LVT U17 ( .A1(n8), .B1(i_cmd[0]), .B2(n38), .ZN(n43) );
  INVD2BWP30P140LVT U18 ( .I(n218), .ZN(n207) );
  OR2D2BWP30P140LVT U19 ( .A1(n20), .A2(n19), .Z(n164) );
  INR2D2BWP30P140LVT U20 ( .A1(n4), .B1(i_cmd[6]), .ZN(n5) );
  INR2D1BWP30P140LVT U21 ( .A1(i_en), .B1(rst), .ZN(n4) );
  NR2OPTPAD1BWP30P140LVT U22 ( .A1(n7), .A2(n21), .ZN(n38) );
  INVD1BWP30P140LVT U23 ( .I(n11), .ZN(n12) );
  ND3D1BWP30P140LVT U24 ( .A1(i_cmd[5]), .A2(i_valid[5]), .A3(n18), .ZN(n19)
         );
  ND2OPTIBD1BWP30P140LVT U25 ( .A1(n38), .A2(n37), .ZN(n49) );
  INVD1BWP30P140LVT U26 ( .I(n225), .ZN(n48) );
  INVD1BWP30P140LVT U27 ( .I(n43), .ZN(n205) );
  INVD1BWP30P140LVT U28 ( .I(n25), .ZN(n218) );
  INVD1BWP30P140LVT U29 ( .I(n43), .ZN(n227) );
  INVD1BWP30P140LVT U30 ( .I(n218), .ZN(n229) );
  INVD1BWP30P140LVT U31 ( .I(n43), .ZN(n88) );
  INVD2BWP30P140LVT U32 ( .I(n216), .ZN(n228) );
  INVD1BWP30P140LVT U33 ( .I(n35), .ZN(n89) );
  INVD1BWP30P140LVT U34 ( .I(i_cmd[3]), .ZN(n31) );
  INR2D1BWP30P140LVT U35 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n3) );
  INVD1BWP30P140LVT U36 ( .I(n3), .ZN(n8) );
  OR2D1BWP30P140LVT U37 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n26) );
  OR2D1BWP30P140LVT U38 ( .A1(n26), .A2(i_cmd[1]), .Z(n7) );
  NR2OPTPAD1BWP30P140LVT U39 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .ZN(n6) );
  NR3D0P7BWP30P140LVT U40 ( .A1(n9), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n14) );
  INVD1BWP30P140LVT U41 ( .I(i_cmd[1]), .ZN(n23) );
  INVD1BWP30P140LVT U42 ( .I(i_cmd[2]), .ZN(n10) );
  CKND2D2BWP30P140LVT U43 ( .A1(n23), .A2(n10), .ZN(n30) );
  INR2D1BWP30P140LVT U44 ( .A1(i_en), .B1(rst), .ZN(n11) );
  NR4D1BWP30P140LVT U45 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .A3(i_cmd[3]), .A4(n12), .ZN(n13) );
  INR2D2BWP30P140LVT U46 ( .A1(n14), .B1(n20), .ZN(n225) );
  INVD1BWP30P140LVT U47 ( .I(i_cmd[6]), .ZN(n15) );
  INR2D2BWP30P140LVT U48 ( .A1(n16), .B1(n20), .ZN(n17) );
  INVD3BWP30P140LVT U49 ( .I(n17), .ZN(n223) );
  NR4D0BWP30P140LVT U50 ( .A1(n88), .A2(n225), .A3(n1), .A4(n2), .ZN(n41) );
  ND4D1BWP30P140LVT U51 ( .A1(n23), .A2(n31), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n24) );
  INR2D1BWP30P140LVT U52 ( .A1(n34), .B1(n24), .ZN(n25) );
  INVD1BWP30P140LVT U53 ( .I(n26), .ZN(n27) );
  ND3D1BWP30P140LVT U54 ( .A1(n27), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n28)
         );
  INR2D1BWP30P140LVT U55 ( .A1(n34), .B1(n28), .ZN(n29) );
  NR2D1BWP30P140LVT U56 ( .A1(n207), .A2(n228), .ZN(n40) );
  INVD1BWP30P140LVT U57 ( .I(n30), .ZN(n32) );
  ND3D1BWP30P140LVT U58 ( .A1(n32), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n33)
         );
  INR2D1BWP30P140LVT U59 ( .A1(n34), .B1(n33), .ZN(n35) );
  IND3D1BWP30P140LVT U60 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n36) );
  INVD1BWP30P140LVT U61 ( .I(n36), .ZN(n37) );
  INVD2BWP30P140LVT U62 ( .I(n49), .ZN(n230) );
  NR2D1BWP30P140LVT U63 ( .A1(n35), .A2(n230), .ZN(n39) );
  ND3D1BWP30P140LVT U64 ( .A1(n41), .A2(n40), .A3(n39), .ZN(N402) );
  INVD1BWP30P140LVT U65 ( .I(i_data_bus[224]), .ZN(n47) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[192]), .ZN(n42) );
  MAOI22D1BWP30P140LVT U67 ( .A1(n2), .A2(i_data_bus[160]), .B1(n223), .B2(n42), .ZN(n46) );
  INR2D1BWP30P140LVT U68 ( .A1(i_data_bus[0]), .B1(n43), .ZN(n44) );
  INVD1BWP30P140LVT U69 ( .I(n44), .ZN(n45) );
  OA211D1BWP30P140LVT U70 ( .A1(n48), .A2(n47), .B(n46), .C(n45), .Z(n52) );
  AOI22D1BWP30P140LVT U71 ( .A1(n207), .A2(i_data_bus[64]), .B1(n206), .B2(
        i_data_bus[32]), .ZN(n51) );
  INVD2BWP30P140LVT U72 ( .I(n89), .ZN(n209) );
  AOI22D1BWP30P140LVT U73 ( .A1(n209), .A2(i_data_bus[96]), .B1(n208), .B2(
        i_data_bus[128]), .ZN(n50) );
  ND3D1BWP30P140LVT U74 ( .A1(n52), .A2(n51), .A3(n50), .ZN(N369) );
  AOI22D1BWP30P140LVT U75 ( .A1(n1), .A2(i_data_bus[220]), .B1(n2), .B2(
        i_data_bus[188]), .ZN(n53) );
  IOA21D1BWP30P140LVT U76 ( .A1(n225), .A2(i_data_bus[252]), .B(n53), .ZN(n54)
         );
  AOI21D1BWP30P140LVT U77 ( .A1(n88), .A2(i_data_bus[28]), .B(n54), .ZN(n57)
         );
  AOI22D1BWP30P140LVT U78 ( .A1(n207), .A2(i_data_bus[92]), .B1(n228), .B2(
        i_data_bus[60]), .ZN(n56) );
  AOI22D1BWP30P140LVT U79 ( .A1(n231), .A2(i_data_bus[124]), .B1(n230), .B2(
        i_data_bus[156]), .ZN(n55) );
  ND3D1BWP30P140LVT U80 ( .A1(n57), .A2(n56), .A3(n55), .ZN(N397) );
  AOI22D1BWP30P140LVT U81 ( .A1(n1), .A2(i_data_bus[218]), .B1(n2), .B2(
        i_data_bus[186]), .ZN(n58) );
  IOA21D1BWP30P140LVT U82 ( .A1(n225), .A2(i_data_bus[250]), .B(n58), .ZN(n59)
         );
  AOI21D1BWP30P140LVT U83 ( .A1(n88), .A2(i_data_bus[26]), .B(n59), .ZN(n62)
         );
  AOI22D1BWP30P140LVT U84 ( .A1(n207), .A2(i_data_bus[90]), .B1(n228), .B2(
        i_data_bus[58]), .ZN(n61) );
  AOI22D1BWP30P140LVT U85 ( .A1(n209), .A2(i_data_bus[122]), .B1(n230), .B2(
        i_data_bus[154]), .ZN(n60) );
  ND3D1BWP30P140LVT U86 ( .A1(n62), .A2(n61), .A3(n60), .ZN(N395) );
  INVD1BWP30P140LVT U87 ( .I(i_data_bus[221]), .ZN(n63) );
  MAOI22D1BWP30P140LVT U88 ( .A1(n2), .A2(i_data_bus[189]), .B1(n223), .B2(n63), .ZN(n64) );
  IOA21D1BWP30P140LVT U89 ( .A1(n225), .A2(i_data_bus[253]), .B(n64), .ZN(n65)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n88), .A2(i_data_bus[29]), .B(n65), .ZN(n68)
         );
  AOI22D1BWP30P140LVT U91 ( .A1(n207), .A2(i_data_bus[93]), .B1(n228), .B2(
        i_data_bus[61]), .ZN(n67) );
  AOI22D1BWP30P140LVT U92 ( .A1(n231), .A2(i_data_bus[125]), .B1(n230), .B2(
        i_data_bus[157]), .ZN(n66) );
  ND3D1BWP30P140LVT U93 ( .A1(n68), .A2(n67), .A3(n66), .ZN(N398) );
  INVD1BWP30P140LVT U94 ( .I(i_data_bus[222]), .ZN(n69) );
  MAOI22D1BWP30P140LVT U95 ( .A1(n2), .A2(i_data_bus[190]), .B1(n223), .B2(n69), .ZN(n70) );
  IOA21D1BWP30P140LVT U96 ( .A1(n225), .A2(i_data_bus[254]), .B(n70), .ZN(n71)
         );
  AOI21D1BWP30P140LVT U97 ( .A1(n88), .A2(i_data_bus[30]), .B(n71), .ZN(n74)
         );
  AOI22D1BWP30P140LVT U98 ( .A1(n207), .A2(i_data_bus[94]), .B1(n228), .B2(
        i_data_bus[62]), .ZN(n73) );
  AOI22D1BWP30P140LVT U99 ( .A1(n209), .A2(i_data_bus[126]), .B1(n230), .B2(
        i_data_bus[158]), .ZN(n72) );
  ND3D1BWP30P140LVT U100 ( .A1(n74), .A2(n73), .A3(n72), .ZN(N399) );
  INVD1BWP30P140LVT U101 ( .I(i_data_bus[223]), .ZN(n75) );
  MAOI22D1BWP30P140LVT U102 ( .A1(n2), .A2(i_data_bus[191]), .B1(n223), .B2(
        n75), .ZN(n76) );
  IOA21D1BWP30P140LVT U103 ( .A1(n225), .A2(i_data_bus[255]), .B(n76), .ZN(n77) );
  AOI21D1BWP30P140LVT U104 ( .A1(n88), .A2(i_data_bus[31]), .B(n77), .ZN(n80)
         );
  AOI22D1BWP30P140LVT U105 ( .A1(n207), .A2(i_data_bus[95]), .B1(n228), .B2(
        i_data_bus[63]), .ZN(n79) );
  AOI22D1BWP30P140LVT U106 ( .A1(n35), .A2(i_data_bus[127]), .B1(n230), .B2(
        i_data_bus[159]), .ZN(n78) );
  ND3D1BWP30P140LVT U107 ( .A1(n80), .A2(n79), .A3(n78), .ZN(N400) );
  AOI22D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[219]), .B1(n2), .B2(
        i_data_bus[187]), .ZN(n81) );
  IOA21D1BWP30P140LVT U109 ( .A1(n225), .A2(i_data_bus[251]), .B(n81), .ZN(n82) );
  AOI21D1BWP30P140LVT U110 ( .A1(n88), .A2(i_data_bus[27]), .B(n82), .ZN(n85)
         );
  AOI22D1BWP30P140LVT U111 ( .A1(n207), .A2(i_data_bus[91]), .B1(n228), .B2(
        i_data_bus[59]), .ZN(n84) );
  AOI22D1BWP30P140LVT U112 ( .A1(n35), .A2(i_data_bus[123]), .B1(n230), .B2(
        i_data_bus[155]), .ZN(n83) );
  ND3D1BWP30P140LVT U113 ( .A1(n85), .A2(n84), .A3(n83), .ZN(N396) );
  AOI22D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[217]), .B1(n2), .B2(
        i_data_bus[185]), .ZN(n86) );
  IOA21D1BWP30P140LVT U115 ( .A1(n225), .A2(i_data_bus[249]), .B(n86), .ZN(n87) );
  AOI21D1BWP30P140LVT U116 ( .A1(n88), .A2(i_data_bus[25]), .B(n87), .ZN(n92)
         );
  AOI22D1BWP30P140LVT U117 ( .A1(n229), .A2(i_data_bus[89]), .B1(n228), .B2(
        i_data_bus[57]), .ZN(n91) );
  INVD2BWP30P140LVT U118 ( .I(n89), .ZN(n231) );
  AOI22D1BWP30P140LVT U119 ( .A1(n231), .A2(i_data_bus[121]), .B1(n230), .B2(
        i_data_bus[153]), .ZN(n90) );
  ND3D1BWP30P140LVT U120 ( .A1(n92), .A2(n91), .A3(n90), .ZN(N394) );
  AOI22D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[198]), .B1(n2), .B2(
        i_data_bus[166]), .ZN(n93) );
  IOA21D1BWP30P140LVT U122 ( .A1(n225), .A2(i_data_bus[230]), .B(n93), .ZN(n94) );
  AOI22D1BWP30P140LVT U123 ( .A1(n207), .A2(i_data_bus[70]), .B1(n206), .B2(
        i_data_bus[38]), .ZN(n96) );
  AOI22D1BWP30P140LVT U124 ( .A1(n209), .A2(i_data_bus[102]), .B1(n208), .B2(
        i_data_bus[134]), .ZN(n95) );
  ND3D1BWP30P140LVT U125 ( .A1(n97), .A2(n96), .A3(n95), .ZN(N375) );
  AOI22D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[197]), .B1(n2), .B2(
        i_data_bus[165]), .ZN(n98) );
  IOA21D1BWP30P140LVT U127 ( .A1(n225), .A2(i_data_bus[229]), .B(n98), .ZN(n99) );
  AOI22D1BWP30P140LVT U128 ( .A1(n207), .A2(i_data_bus[69]), .B1(n206), .B2(
        i_data_bus[37]), .ZN(n101) );
  AOI22D1BWP30P140LVT U129 ( .A1(n209), .A2(i_data_bus[101]), .B1(n208), .B2(
        i_data_bus[133]), .ZN(n100) );
  ND3D1BWP30P140LVT U130 ( .A1(n102), .A2(n101), .A3(n100), .ZN(N374) );
  AOI22D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[196]), .B1(n2), .B2(
        i_data_bus[164]), .ZN(n103) );
  IOA21D1BWP30P140LVT U132 ( .A1(n225), .A2(i_data_bus[228]), .B(n103), .ZN(
        n104) );
  AOI21D1BWP30P140LVT U133 ( .A1(n205), .A2(i_data_bus[4]), .B(n104), .ZN(n107) );
  AOI22D1BWP30P140LVT U134 ( .A1(n207), .A2(i_data_bus[68]), .B1(n206), .B2(
        i_data_bus[36]), .ZN(n106) );
  AOI22D1BWP30P140LVT U135 ( .A1(n209), .A2(i_data_bus[100]), .B1(n208), .B2(
        i_data_bus[132]), .ZN(n105) );
  ND3D1BWP30P140LVT U136 ( .A1(n107), .A2(n106), .A3(n105), .ZN(N373) );
  AOI22D1BWP30P140LVT U137 ( .A1(n1), .A2(i_data_bus[199]), .B1(n2), .B2(
        i_data_bus[167]), .ZN(n108) );
  IOA21D1BWP30P140LVT U138 ( .A1(n225), .A2(i_data_bus[231]), .B(n108), .ZN(
        n109) );
  AOI21D1BWP30P140LVT U139 ( .A1(n205), .A2(i_data_bus[7]), .B(n109), .ZN(n112) );
  AOI22D1BWP30P140LVT U140 ( .A1(n207), .A2(i_data_bus[71]), .B1(n206), .B2(
        i_data_bus[39]), .ZN(n111) );
  AOI22D1BWP30P140LVT U141 ( .A1(n209), .A2(i_data_bus[103]), .B1(n208), .B2(
        i_data_bus[135]), .ZN(n110) );
  ND3D1BWP30P140LVT U142 ( .A1(n112), .A2(n111), .A3(n110), .ZN(N376) );
  AOI22D1BWP30P140LVT U143 ( .A1(n1), .A2(i_data_bus[201]), .B1(n2), .B2(
        i_data_bus[169]), .ZN(n113) );
  IOA21D1BWP30P140LVT U144 ( .A1(n225), .A2(i_data_bus[233]), .B(n113), .ZN(
        n114) );
  AOI21D1BWP30P140LVT U145 ( .A1(n205), .A2(i_data_bus[9]), .B(n114), .ZN(n117) );
  AOI22D1BWP30P140LVT U146 ( .A1(n207), .A2(i_data_bus[73]), .B1(n206), .B2(
        i_data_bus[41]), .ZN(n116) );
  AOI22D1BWP30P140LVT U147 ( .A1(n209), .A2(i_data_bus[105]), .B1(n208), .B2(
        i_data_bus[137]), .ZN(n115) );
  ND3D1BWP30P140LVT U148 ( .A1(n117), .A2(n116), .A3(n115), .ZN(N378) );
  AOI22D1BWP30P140LVT U149 ( .A1(n1), .A2(i_data_bus[200]), .B1(n2), .B2(
        i_data_bus[168]), .ZN(n118) );
  IOA21D1BWP30P140LVT U150 ( .A1(n225), .A2(i_data_bus[232]), .B(n118), .ZN(
        n119) );
  AOI21D1BWP30P140LVT U151 ( .A1(n205), .A2(i_data_bus[8]), .B(n119), .ZN(n122) );
  AOI22D1BWP30P140LVT U152 ( .A1(n207), .A2(i_data_bus[72]), .B1(n206), .B2(
        i_data_bus[40]), .ZN(n121) );
  AOI22D1BWP30P140LVT U153 ( .A1(n209), .A2(i_data_bus[104]), .B1(n208), .B2(
        i_data_bus[136]), .ZN(n120) );
  ND3D1BWP30P140LVT U154 ( .A1(n122), .A2(n121), .A3(n120), .ZN(N377) );
  AOI22D1BWP30P140LVT U155 ( .A1(n1), .A2(i_data_bus[203]), .B1(n2), .B2(
        i_data_bus[171]), .ZN(n123) );
  IOA21D1BWP30P140LVT U156 ( .A1(n225), .A2(i_data_bus[235]), .B(n123), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U157 ( .A1(n205), .A2(i_data_bus[11]), .B(n124), .ZN(
        n127) );
  AOI22D1BWP30P140LVT U158 ( .A1(n207), .A2(i_data_bus[75]), .B1(n206), .B2(
        i_data_bus[43]), .ZN(n126) );
  AOI22D1BWP30P140LVT U159 ( .A1(n209), .A2(i_data_bus[107]), .B1(n208), .B2(
        i_data_bus[139]), .ZN(n125) );
  ND3D1BWP30P140LVT U160 ( .A1(n127), .A2(n126), .A3(n125), .ZN(N380) );
  AOI22D1BWP30P140LVT U161 ( .A1(n1), .A2(i_data_bus[202]), .B1(n2), .B2(
        i_data_bus[170]), .ZN(n128) );
  IOA21D1BWP30P140LVT U162 ( .A1(n225), .A2(i_data_bus[234]), .B(n128), .ZN(
        n129) );
  AOI21D1BWP30P140LVT U163 ( .A1(n205), .A2(i_data_bus[10]), .B(n129), .ZN(
        n132) );
  AOI22D1BWP30P140LVT U164 ( .A1(n207), .A2(i_data_bus[74]), .B1(n206), .B2(
        i_data_bus[42]), .ZN(n131) );
  AOI22D1BWP30P140LVT U165 ( .A1(n209), .A2(i_data_bus[106]), .B1(n208), .B2(
        i_data_bus[138]), .ZN(n130) );
  ND3D1BWP30P140LVT U166 ( .A1(n132), .A2(n131), .A3(n130), .ZN(N379) );
  AOI22D1BWP30P140LVT U167 ( .A1(n1), .A2(i_data_bus[204]), .B1(n2), .B2(
        i_data_bus[172]), .ZN(n133) );
  IOA21D1BWP30P140LVT U168 ( .A1(n225), .A2(i_data_bus[236]), .B(n133), .ZN(
        n134) );
  AOI21D1BWP30P140LVT U169 ( .A1(n205), .A2(i_data_bus[12]), .B(n134), .ZN(
        n137) );
  AOI22D1BWP30P140LVT U170 ( .A1(n207), .A2(i_data_bus[76]), .B1(n206), .B2(
        i_data_bus[44]), .ZN(n136) );
  AOI22D1BWP30P140LVT U171 ( .A1(n209), .A2(i_data_bus[108]), .B1(n208), .B2(
        i_data_bus[140]), .ZN(n135) );
  ND3D1BWP30P140LVT U172 ( .A1(n137), .A2(n136), .A3(n135), .ZN(N381) );
  AOI22D1BWP30P140LVT U173 ( .A1(n1), .A2(i_data_bus[213]), .B1(n2), .B2(
        i_data_bus[181]), .ZN(n138) );
  IOA21D1BWP30P140LVT U174 ( .A1(n225), .A2(i_data_bus[245]), .B(n138), .ZN(
        n139) );
  AOI21D1BWP30P140LVT U175 ( .A1(n227), .A2(i_data_bus[21]), .B(n139), .ZN(
        n142) );
  AOI22D1BWP30P140LVT U176 ( .A1(n229), .A2(i_data_bus[85]), .B1(n228), .B2(
        i_data_bus[53]), .ZN(n141) );
  AOI22D1BWP30P140LVT U177 ( .A1(n231), .A2(i_data_bus[117]), .B1(n230), .B2(
        i_data_bus[149]), .ZN(n140) );
  ND3D1BWP30P140LVT U178 ( .A1(n142), .A2(n141), .A3(n140), .ZN(N390) );
  AOI22D1BWP30P140LVT U179 ( .A1(n1), .A2(i_data_bus[212]), .B1(n2), .B2(
        i_data_bus[180]), .ZN(n143) );
  IOA21D1BWP30P140LVT U180 ( .A1(n225), .A2(i_data_bus[244]), .B(n143), .ZN(
        n144) );
  AOI21D1BWP30P140LVT U181 ( .A1(n227), .A2(i_data_bus[20]), .B(n144), .ZN(
        n147) );
  AOI22D1BWP30P140LVT U182 ( .A1(n229), .A2(i_data_bus[84]), .B1(n228), .B2(
        i_data_bus[52]), .ZN(n146) );
  AOI22D1BWP30P140LVT U183 ( .A1(n231), .A2(i_data_bus[116]), .B1(n230), .B2(
        i_data_bus[148]), .ZN(n145) );
  ND3D1BWP30P140LVT U184 ( .A1(n147), .A2(n146), .A3(n145), .ZN(N389) );
  AOI22D1BWP30P140LVT U185 ( .A1(n1), .A2(i_data_bus[215]), .B1(n2), .B2(
        i_data_bus[183]), .ZN(n148) );
  IOA21D1BWP30P140LVT U186 ( .A1(n225), .A2(i_data_bus[247]), .B(n148), .ZN(
        n149) );
  AOI21D1BWP30P140LVT U187 ( .A1(n227), .A2(i_data_bus[23]), .B(n149), .ZN(
        n152) );
  AOI22D1BWP30P140LVT U188 ( .A1(n229), .A2(i_data_bus[87]), .B1(n228), .B2(
        i_data_bus[55]), .ZN(n151) );
  AOI22D1BWP30P140LVT U189 ( .A1(n231), .A2(i_data_bus[119]), .B1(n230), .B2(
        i_data_bus[151]), .ZN(n150) );
  ND3D1BWP30P140LVT U190 ( .A1(n152), .A2(n151), .A3(n150), .ZN(N392) );
  AOI22D1BWP30P140LVT U191 ( .A1(n1), .A2(i_data_bus[214]), .B1(n2), .B2(
        i_data_bus[182]), .ZN(n153) );
  IOA21D1BWP30P140LVT U192 ( .A1(n225), .A2(i_data_bus[246]), .B(n153), .ZN(
        n154) );
  AOI21D1BWP30P140LVT U193 ( .A1(n227), .A2(i_data_bus[22]), .B(n154), .ZN(
        n157) );
  AOI22D1BWP30P140LVT U194 ( .A1(n229), .A2(i_data_bus[86]), .B1(n228), .B2(
        i_data_bus[54]), .ZN(n156) );
  AOI22D1BWP30P140LVT U195 ( .A1(n231), .A2(i_data_bus[118]), .B1(n230), .B2(
        i_data_bus[150]), .ZN(n155) );
  ND3D1BWP30P140LVT U196 ( .A1(n157), .A2(n156), .A3(n155), .ZN(N391) );
  AOI22D1BWP30P140LVT U197 ( .A1(n1), .A2(i_data_bus[206]), .B1(n2), .B2(
        i_data_bus[174]), .ZN(n158) );
  IOA21D1BWP30P140LVT U198 ( .A1(n225), .A2(i_data_bus[238]), .B(n158), .ZN(
        n159) );
  AOI21D1BWP30P140LVT U199 ( .A1(n227), .A2(i_data_bus[14]), .B(n159), .ZN(
        n162) );
  AOI22D1BWP30P140LVT U200 ( .A1(n229), .A2(i_data_bus[78]), .B1(n228), .B2(
        i_data_bus[46]), .ZN(n161) );
  AOI22D1BWP30P140LVT U201 ( .A1(n231), .A2(i_data_bus[110]), .B1(n230), .B2(
        i_data_bus[142]), .ZN(n160) );
  ND3D1BWP30P140LVT U202 ( .A1(n162), .A2(n161), .A3(n160), .ZN(N383) );
  INVD1BWP30P140LVT U203 ( .I(i_data_bus[173]), .ZN(n163) );
  MAOI22D1BWP30P140LVT U204 ( .A1(n1), .A2(i_data_bus[205]), .B1(n164), .B2(
        n163), .ZN(n165) );
  IOA21D1BWP30P140LVT U205 ( .A1(n225), .A2(i_data_bus[237]), .B(n165), .ZN(
        n166) );
  AOI21D1BWP30P140LVT U206 ( .A1(n227), .A2(i_data_bus[13]), .B(n166), .ZN(
        n169) );
  AOI22D1BWP30P140LVT U207 ( .A1(n229), .A2(i_data_bus[77]), .B1(n228), .B2(
        i_data_bus[45]), .ZN(n168) );
  AOI22D1BWP30P140LVT U208 ( .A1(n231), .A2(i_data_bus[109]), .B1(n230), .B2(
        i_data_bus[141]), .ZN(n167) );
  ND3D1BWP30P140LVT U209 ( .A1(n169), .A2(n168), .A3(n167), .ZN(N382) );
  AOI22D1BWP30P140LVT U210 ( .A1(n1), .A2(i_data_bus[211]), .B1(n2), .B2(
        i_data_bus[179]), .ZN(n170) );
  IOA21D1BWP30P140LVT U211 ( .A1(n225), .A2(i_data_bus[243]), .B(n170), .ZN(
        n171) );
  AOI21D1BWP30P140LVT U212 ( .A1(n227), .A2(i_data_bus[19]), .B(n171), .ZN(
        n174) );
  AOI22D1BWP30P140LVT U213 ( .A1(n229), .A2(i_data_bus[83]), .B1(n228), .B2(
        i_data_bus[51]), .ZN(n173) );
  AOI22D1BWP30P140LVT U214 ( .A1(n231), .A2(i_data_bus[115]), .B1(n230), .B2(
        i_data_bus[147]), .ZN(n172) );
  ND3D1BWP30P140LVT U215 ( .A1(n174), .A2(n173), .A3(n172), .ZN(N388) );
  AOI22D1BWP30P140LVT U216 ( .A1(n1), .A2(i_data_bus[210]), .B1(n2), .B2(
        i_data_bus[178]), .ZN(n175) );
  IOA21D1BWP30P140LVT U217 ( .A1(n225), .A2(i_data_bus[242]), .B(n175), .ZN(
        n176) );
  AOI21D1BWP30P140LVT U218 ( .A1(n227), .A2(i_data_bus[18]), .B(n176), .ZN(
        n179) );
  AOI22D1BWP30P140LVT U219 ( .A1(n229), .A2(i_data_bus[82]), .B1(n228), .B2(
        i_data_bus[50]), .ZN(n178) );
  AOI22D1BWP30P140LVT U220 ( .A1(n231), .A2(i_data_bus[114]), .B1(n230), .B2(
        i_data_bus[146]), .ZN(n177) );
  ND3D1BWP30P140LVT U221 ( .A1(n179), .A2(n178), .A3(n177), .ZN(N387) );
  AOI22D1BWP30P140LVT U222 ( .A1(n1), .A2(i_data_bus[209]), .B1(n2), .B2(
        i_data_bus[177]), .ZN(n180) );
  IOA21D1BWP30P140LVT U223 ( .A1(n225), .A2(i_data_bus[241]), .B(n180), .ZN(
        n181) );
  AOI21D1BWP30P140LVT U224 ( .A1(n227), .A2(i_data_bus[17]), .B(n181), .ZN(
        n184) );
  AOI22D1BWP30P140LVT U225 ( .A1(n229), .A2(i_data_bus[81]), .B1(n228), .B2(
        i_data_bus[49]), .ZN(n183) );
  AOI22D1BWP30P140LVT U226 ( .A1(n231), .A2(i_data_bus[113]), .B1(n230), .B2(
        i_data_bus[145]), .ZN(n182) );
  ND3D1BWP30P140LVT U227 ( .A1(n184), .A2(n183), .A3(n182), .ZN(N386) );
  AOI22D1BWP30P140LVT U228 ( .A1(n1), .A2(i_data_bus[216]), .B1(n2), .B2(
        i_data_bus[184]), .ZN(n185) );
  IOA21D1BWP30P140LVT U229 ( .A1(n225), .A2(i_data_bus[248]), .B(n185), .ZN(
        n186) );
  AOI21D1BWP30P140LVT U230 ( .A1(n227), .A2(i_data_bus[24]), .B(n186), .ZN(
        n189) );
  AOI22D1BWP30P140LVT U231 ( .A1(n229), .A2(i_data_bus[88]), .B1(n228), .B2(
        i_data_bus[56]), .ZN(n188) );
  AOI22D1BWP30P140LVT U232 ( .A1(n231), .A2(i_data_bus[120]), .B1(n230), .B2(
        i_data_bus[152]), .ZN(n187) );
  ND3D1BWP30P140LVT U233 ( .A1(n189), .A2(n188), .A3(n187), .ZN(N393) );
  INVD1BWP30P140LVT U234 ( .I(i_data_bus[195]), .ZN(n190) );
  MAOI22D1BWP30P140LVT U235 ( .A1(n2), .A2(i_data_bus[163]), .B1(n223), .B2(
        n190), .ZN(n191) );
  IOA21D1BWP30P140LVT U236 ( .A1(n225), .A2(i_data_bus[227]), .B(n191), .ZN(
        n192) );
  AOI21D1BWP30P140LVT U237 ( .A1(n205), .A2(i_data_bus[3]), .B(n192), .ZN(n195) );
  AOI22D1BWP30P140LVT U238 ( .A1(n207), .A2(i_data_bus[67]), .B1(n206), .B2(
        i_data_bus[35]), .ZN(n194) );
  AOI22D1BWP30P140LVT U239 ( .A1(n209), .A2(i_data_bus[99]), .B1(n208), .B2(
        i_data_bus[131]), .ZN(n193) );
  ND3D1BWP30P140LVT U240 ( .A1(n195), .A2(n194), .A3(n193), .ZN(N372) );
  INVD1BWP30P140LVT U241 ( .I(i_data_bus[194]), .ZN(n196) );
  MAOI22D1BWP30P140LVT U242 ( .A1(n2), .A2(i_data_bus[162]), .B1(n223), .B2(
        n196), .ZN(n197) );
  IOA21D1BWP30P140LVT U243 ( .A1(n225), .A2(i_data_bus[226]), .B(n197), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U244 ( .A1(n205), .A2(i_data_bus[2]), .B(n198), .ZN(n201) );
  AOI22D1BWP30P140LVT U245 ( .A1(n207), .A2(i_data_bus[66]), .B1(n206), .B2(
        i_data_bus[34]), .ZN(n200) );
  AOI22D1BWP30P140LVT U246 ( .A1(n209), .A2(i_data_bus[98]), .B1(n208), .B2(
        i_data_bus[130]), .ZN(n199) );
  ND3D1BWP30P140LVT U247 ( .A1(n201), .A2(n200), .A3(n199), .ZN(N371) );
  INVD1BWP30P140LVT U248 ( .I(i_data_bus[193]), .ZN(n202) );
  MAOI22D1BWP30P140LVT U249 ( .A1(n2), .A2(i_data_bus[161]), .B1(n223), .B2(
        n202), .ZN(n203) );
  IOA21D1BWP30P140LVT U250 ( .A1(n225), .A2(i_data_bus[225]), .B(n203), .ZN(
        n204) );
  AOI21D1BWP30P140LVT U251 ( .A1(n205), .A2(i_data_bus[1]), .B(n204), .ZN(n212) );
  AOI22D1BWP30P140LVT U252 ( .A1(n207), .A2(i_data_bus[65]), .B1(n206), .B2(
        i_data_bus[33]), .ZN(n211) );
  AOI22D1BWP30P140LVT U253 ( .A1(n209), .A2(i_data_bus[97]), .B1(n208), .B2(
        i_data_bus[129]), .ZN(n210) );
  ND3D1BWP30P140LVT U254 ( .A1(n212), .A2(n211), .A3(n210), .ZN(N370) );
  AOI22D1BWP30P140LVT U255 ( .A1(n1), .A2(i_data_bus[207]), .B1(n2), .B2(
        i_data_bus[175]), .ZN(n213) );
  IOA21D1BWP30P140LVT U256 ( .A1(n225), .A2(i_data_bus[239]), .B(n213), .ZN(
        n214) );
  AOI21D1BWP30P140LVT U257 ( .A1(n227), .A2(i_data_bus[15]), .B(n214), .ZN(
        n221) );
  INVD1BWP30P140LVT U258 ( .I(i_data_bus[79]), .ZN(n217) );
  INVD1BWP30P140LVT U259 ( .I(i_data_bus[47]), .ZN(n215) );
  OA22D1BWP30P140LVT U260 ( .A1(n218), .A2(n217), .B1(n216), .B2(n215), .Z(
        n220) );
  AOI22D1BWP30P140LVT U261 ( .A1(n231), .A2(i_data_bus[111]), .B1(n230), .B2(
        i_data_bus[143]), .ZN(n219) );
  ND3D1BWP30P140LVT U262 ( .A1(n221), .A2(n220), .A3(n219), .ZN(N384) );
  INVD1BWP30P140LVT U263 ( .I(i_data_bus[208]), .ZN(n222) );
  MAOI22D1BWP30P140LVT U264 ( .A1(n2), .A2(i_data_bus[176]), .B1(n223), .B2(
        n222), .ZN(n224) );
  IOA21D1BWP30P140LVT U265 ( .A1(n225), .A2(i_data_bus[240]), .B(n224), .ZN(
        n226) );
  AOI21D1BWP30P140LVT U266 ( .A1(n227), .A2(i_data_bus[16]), .B(n226), .ZN(
        n234) );
  AOI22D1BWP30P140LVT U267 ( .A1(n229), .A2(i_data_bus[80]), .B1(n228), .B2(
        i_data_bus[48]), .ZN(n233) );
  AOI22D1BWP30P140LVT U268 ( .A1(n231), .A2(i_data_bus[112]), .B1(n230), .B2(
        i_data_bus[144]), .ZN(n232) );
  ND3D1BWP30P140LVT U269 ( .A1(n234), .A2(n233), .A3(n232), .ZN(N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_4 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  BUFFD3BWP30P140LVT U3 ( .I(n227), .Z(n2) );
  INR2D1BWP30P140LVT U4 ( .A1(n18), .B1(n23), .ZN(n227) );
  INR2D1BWP30P140LVT U5 ( .A1(n7), .B1(i_cmd[5]), .ZN(n8) );
  INR4D1BWP30P140LVT U6 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n22), .ZN(n24) );
  INVD1BWP30P140LVT U7 ( .I(n230), .ZN(n205) );
  CKAN2D4BWP30P140LVT U8 ( .A1(n43), .A2(n42), .Z(n1) );
  INVD6BWP30P140LVT U9 ( .I(n174), .ZN(n3) );
  INVD8BWP30P140LVT U10 ( .I(n212), .ZN(n4) );
  INVD2BWP30P140LVT U11 ( .I(n187), .ZN(n5) );
  INR2D2BWP30P140LVT U12 ( .A1(n27), .B1(n26), .ZN(n39) );
  OR2D2BWP30P140LVT U13 ( .A1(n35), .A2(n17), .Z(n23) );
  ND2OPTIBD2BWP30P140LVT U14 ( .A1(n9), .A2(n8), .ZN(n26) );
  INR2D2BWP30P140LVT U15 ( .A1(n24), .B1(n23), .ZN(n25) );
  INVD3BWP30P140LVT U16 ( .I(n21), .ZN(n212) );
  INR2D1BWP30P140LVT U17 ( .A1(i_en), .B1(rst), .ZN(n7) );
  INVD1BWP30P140LVT U18 ( .I(n40), .ZN(n129) );
  INVD1BWP30P140LVT U19 ( .I(n30), .ZN(n232) );
  INVD2BWP30P140LVT U20 ( .I(n34), .ZN(n230) );
  INVD1BWP30P140LVT U21 ( .I(n129), .ZN(n233) );
  INVD1BWP30P140LVT U22 ( .I(n232), .ZN(n222) );
  INVD2BWP30P140LVT U23 ( .I(n230), .ZN(n221) );
  NR2D1BWP30P140LVT U24 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n27) );
  NR3D0P7BWP30P140LVT U25 ( .A1(n19), .A2(i_cmd[5]), .A3(i_cmd[7]), .ZN(n20)
         );
  ND2D1BWP30P140LVT U26 ( .A1(i_valid[6]), .A2(i_cmd[6]), .ZN(n19) );
  NR2D1BWP30P140LVT U27 ( .A1(n10), .A2(n26), .ZN(n43) );
  INVD1BWP30P140LVT U28 ( .I(n129), .ZN(n207) );
  INVD1BWP30P140LVT U29 ( .I(n232), .ZN(n206) );
  INVD1BWP30P140LVT U30 ( .I(n187), .ZN(n220) );
  AOI21D1BWP30P140LVT U31 ( .A1(n220), .A2(i_data_bus[14]), .B(n169), .ZN(n172) );
  INR2D1BWP30P140LVT U32 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n6) );
  INVD1BWP30P140LVT U33 ( .I(n6), .ZN(n11) );
  OR2D1BWP30P140LVT U34 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n31) );
  OR2D1BWP30P140LVT U35 ( .A1(n31), .A2(i_cmd[1]), .Z(n10) );
  NR2OPTPAD1BWP30P140LVT U36 ( .A1(i_cmd[7]), .A2(i_cmd[6]), .ZN(n9) );
  IND3D2BWP30P140LVT U37 ( .A1(n11), .B1(i_cmd[0]), .B2(n43), .ZN(n187) );
  ND2D1BWP30P140LVT U38 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n12) );
  NR3D0P7BWP30P140LVT U39 ( .A1(n12), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n18)
         );
  INVD1BWP30P140LVT U40 ( .I(i_cmd[2]), .ZN(n13) );
  INVD1BWP30P140LVT U41 ( .I(i_cmd[1]), .ZN(n28) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n13), .A2(n28), .ZN(n35) );
  NR2OPTPAD1BWP30P140LVT U43 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n16) );
  INR2D1BWP30P140LVT U44 ( .A1(i_en), .B1(rst), .ZN(n14) );
  INR2D1BWP30P140LVT U45 ( .A1(n14), .B1(i_cmd[3]), .ZN(n15) );
  ND2OPTIBD1BWP30P140LVT U46 ( .A1(n16), .A2(n15), .ZN(n17) );
  INR2D1BWP30P140LVT U47 ( .A1(n20), .B1(n23), .ZN(n21) );
  INVD1BWP30P140LVT U48 ( .I(i_cmd[5]), .ZN(n22) );
  INVD2BWP30P140LVT U49 ( .I(n25), .ZN(n174) );
  NR4D0BWP30P140LVT U50 ( .A1(n220), .A2(n2), .A3(n4), .A4(n3), .ZN(n46) );
  INVD1BWP30P140LVT U51 ( .I(i_cmd[3]), .ZN(n36) );
  ND4D1BWP30P140LVT U52 ( .A1(n28), .A2(n36), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n29) );
  INR2D1BWP30P140LVT U53 ( .A1(n39), .B1(n29), .ZN(n30) );
  INVD1BWP30P140LVT U54 ( .I(n232), .ZN(n77) );
  INVD1BWP30P140LVT U55 ( .I(n31), .ZN(n32) );
  ND3D1BWP30P140LVT U56 ( .A1(n32), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n33)
         );
  INR2D2BWP30P140LVT U57 ( .A1(n39), .B1(n33), .ZN(n34) );
  NR2D1BWP30P140LVT U58 ( .A1(n77), .A2(n221), .ZN(n45) );
  INVD1BWP30P140LVT U59 ( .I(n35), .ZN(n37) );
  ND3D1BWP30P140LVT U60 ( .A1(n37), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n38)
         );
  INR2D1BWP30P140LVT U61 ( .A1(n39), .B1(n38), .ZN(n40) );
  INVD1BWP30P140LVT U62 ( .I(n129), .ZN(n78) );
  IND3D1BWP30P140LVT U63 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n41) );
  INVD1BWP30P140LVT U64 ( .I(n41), .ZN(n42) );
  NR2D1BWP30P140LVT U65 ( .A1(n78), .A2(n1), .ZN(n44) );
  ND3D1BWP30P140LVT U66 ( .A1(n46), .A2(n45), .A3(n44), .ZN(N402) );
  INVD1BWP30P140LVT U67 ( .I(i_data_bus[223]), .ZN(n47) );
  MAOI22D1BWP30P140LVT U68 ( .A1(n3), .A2(i_data_bus[191]), .B1(n212), .B2(n47), .ZN(n48) );
  IOA21D1BWP30P140LVT U69 ( .A1(n2), .A2(i_data_bus[255]), .B(n48), .ZN(n49)
         );
  AOI21D1BWP30P140LVT U70 ( .A1(n5), .A2(i_data_bus[31]), .B(n49), .ZN(n52) );
  AOI22D1BWP30P140LVT U71 ( .A1(n77), .A2(i_data_bus[95]), .B1(n221), .B2(
        i_data_bus[63]), .ZN(n51) );
  AOI22D1BWP30P140LVT U72 ( .A1(n78), .A2(i_data_bus[127]), .B1(n1), .B2(
        i_data_bus[159]), .ZN(n50) );
  ND3D1BWP30P140LVT U73 ( .A1(n52), .A2(n51), .A3(n50), .ZN(N400) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[222]), .ZN(n53) );
  MAOI22D1BWP30P140LVT U75 ( .A1(n3), .A2(i_data_bus[190]), .B1(n212), .B2(n53), .ZN(n54) );
  IOA21D1BWP30P140LVT U76 ( .A1(n2), .A2(i_data_bus[254]), .B(n54), .ZN(n55)
         );
  AOI21D1BWP30P140LVT U77 ( .A1(n5), .A2(i_data_bus[30]), .B(n55), .ZN(n58) );
  AOI22D1BWP30P140LVT U78 ( .A1(n77), .A2(i_data_bus[94]), .B1(n221), .B2(
        i_data_bus[62]), .ZN(n57) );
  AOI22D1BWP30P140LVT U79 ( .A1(n78), .A2(i_data_bus[126]), .B1(n1), .B2(
        i_data_bus[158]), .ZN(n56) );
  ND3D1BWP30P140LVT U80 ( .A1(n58), .A2(n57), .A3(n56), .ZN(N399) );
  AOI22D1BWP30P140LVT U81 ( .A1(n4), .A2(i_data_bus[219]), .B1(n3), .B2(
        i_data_bus[187]), .ZN(n59) );
  IOA21D1BWP30P140LVT U82 ( .A1(n2), .A2(i_data_bus[251]), .B(n59), .ZN(n60)
         );
  AOI21D1BWP30P140LVT U83 ( .A1(n220), .A2(i_data_bus[27]), .B(n60), .ZN(n63)
         );
  AOI22D1BWP30P140LVT U84 ( .A1(n77), .A2(i_data_bus[91]), .B1(n221), .B2(
        i_data_bus[59]), .ZN(n62) );
  AOI22D1BWP30P140LVT U85 ( .A1(n78), .A2(i_data_bus[123]), .B1(n1), .B2(
        i_data_bus[155]), .ZN(n61) );
  ND3D1BWP30P140LVT U86 ( .A1(n63), .A2(n62), .A3(n61), .ZN(N396) );
  AOI22D1BWP30P140LVT U87 ( .A1(n4), .A2(i_data_bus[218]), .B1(n3), .B2(
        i_data_bus[186]), .ZN(n64) );
  IOA21D1BWP30P140LVT U88 ( .A1(n2), .A2(i_data_bus[250]), .B(n64), .ZN(n65)
         );
  AOI21D1BWP30P140LVT U89 ( .A1(n5), .A2(i_data_bus[26]), .B(n65), .ZN(n68) );
  AOI22D1BWP30P140LVT U90 ( .A1(n77), .A2(i_data_bus[90]), .B1(n221), .B2(
        i_data_bus[58]), .ZN(n67) );
  AOI22D1BWP30P140LVT U91 ( .A1(n78), .A2(i_data_bus[122]), .B1(n1), .B2(
        i_data_bus[154]), .ZN(n66) );
  ND3D1BWP30P140LVT U92 ( .A1(n68), .A2(n67), .A3(n66), .ZN(N395) );
  AOI22D1BWP30P140LVT U93 ( .A1(n4), .A2(i_data_bus[220]), .B1(n3), .B2(
        i_data_bus[188]), .ZN(n69) );
  IOA21D1BWP30P140LVT U94 ( .A1(n2), .A2(i_data_bus[252]), .B(n69), .ZN(n70)
         );
  AOI21D1BWP30P140LVT U95 ( .A1(n5), .A2(i_data_bus[28]), .B(n70), .ZN(n73) );
  AOI22D1BWP30P140LVT U96 ( .A1(n77), .A2(i_data_bus[92]), .B1(n221), .B2(
        i_data_bus[60]), .ZN(n72) );
  AOI22D1BWP30P140LVT U97 ( .A1(n78), .A2(i_data_bus[124]), .B1(n1), .B2(
        i_data_bus[156]), .ZN(n71) );
  ND3D1BWP30P140LVT U98 ( .A1(n73), .A2(n72), .A3(n71), .ZN(N397) );
  INVD1BWP30P140LVT U99 ( .I(i_data_bus[221]), .ZN(n74) );
  MAOI22D1BWP30P140LVT U100 ( .A1(n3), .A2(i_data_bus[189]), .B1(n212), .B2(
        n74), .ZN(n75) );
  IOA21D1BWP30P140LVT U101 ( .A1(n2), .A2(i_data_bus[253]), .B(n75), .ZN(n76)
         );
  AOI21D1BWP30P140LVT U102 ( .A1(n220), .A2(i_data_bus[29]), .B(n76), .ZN(n81)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n77), .A2(i_data_bus[93]), .B1(n221), .B2(
        i_data_bus[61]), .ZN(n80) );
  AOI22D1BWP30P140LVT U104 ( .A1(n78), .A2(i_data_bus[125]), .B1(n1), .B2(
        i_data_bus[157]), .ZN(n79) );
  ND3D1BWP30P140LVT U105 ( .A1(n81), .A2(n80), .A3(n79), .ZN(N398) );
  AOI22D1BWP30P140LVT U106 ( .A1(n4), .A2(i_data_bus[196]), .B1(n3), .B2(
        i_data_bus[164]), .ZN(n82) );
  IOA21D1BWP30P140LVT U107 ( .A1(n2), .A2(i_data_bus[228]), .B(n82), .ZN(n83)
         );
  AOI21D1BWP30P140LVT U108 ( .A1(n5), .A2(i_data_bus[4]), .B(n83), .ZN(n86) );
  AOI22D1BWP30P140LVT U109 ( .A1(n206), .A2(i_data_bus[68]), .B1(n205), .B2(
        i_data_bus[36]), .ZN(n85) );
  AOI22D1BWP30P140LVT U110 ( .A1(n207), .A2(i_data_bus[100]), .B1(n1), .B2(
        i_data_bus[132]), .ZN(n84) );
  ND3D1BWP30P140LVT U111 ( .A1(n86), .A2(n85), .A3(n84), .ZN(N373) );
  AOI22D1BWP30P140LVT U112 ( .A1(n4), .A2(i_data_bus[200]), .B1(n3), .B2(
        i_data_bus[168]), .ZN(n87) );
  IOA21D1BWP30P140LVT U113 ( .A1(n2), .A2(i_data_bus[232]), .B(n87), .ZN(n88)
         );
  AOI21D1BWP30P140LVT U114 ( .A1(n5), .A2(i_data_bus[8]), .B(n88), .ZN(n91) );
  AOI22D1BWP30P140LVT U115 ( .A1(n206), .A2(i_data_bus[72]), .B1(n205), .B2(
        i_data_bus[40]), .ZN(n90) );
  AOI22D1BWP30P140LVT U116 ( .A1(n207), .A2(i_data_bus[104]), .B1(n1), .B2(
        i_data_bus[136]), .ZN(n89) );
  ND3D1BWP30P140LVT U117 ( .A1(n91), .A2(n90), .A3(n89), .ZN(N377) );
  AOI22D1BWP30P140LVT U118 ( .A1(n4), .A2(i_data_bus[199]), .B1(n3), .B2(
        i_data_bus[167]), .ZN(n92) );
  IOA21D1BWP30P140LVT U119 ( .A1(n2), .A2(i_data_bus[231]), .B(n92), .ZN(n93)
         );
  AOI21D1BWP30P140LVT U120 ( .A1(n220), .A2(i_data_bus[7]), .B(n93), .ZN(n96)
         );
  AOI22D1BWP30P140LVT U121 ( .A1(n206), .A2(i_data_bus[71]), .B1(n205), .B2(
        i_data_bus[39]), .ZN(n95) );
  AOI22D1BWP30P140LVT U122 ( .A1(n207), .A2(i_data_bus[103]), .B1(n1), .B2(
        i_data_bus[135]), .ZN(n94) );
  ND3D1BWP30P140LVT U123 ( .A1(n96), .A2(n95), .A3(n94), .ZN(N376) );
  AOI22D1BWP30P140LVT U124 ( .A1(n4), .A2(i_data_bus[198]), .B1(n3), .B2(
        i_data_bus[166]), .ZN(n97) );
  IOA21D1BWP30P140LVT U125 ( .A1(n2), .A2(i_data_bus[230]), .B(n97), .ZN(n98)
         );
  AOI21D1BWP30P140LVT U126 ( .A1(n5), .A2(i_data_bus[6]), .B(n98), .ZN(n101)
         );
  AOI22D1BWP30P140LVT U127 ( .A1(n206), .A2(i_data_bus[70]), .B1(n205), .B2(
        i_data_bus[38]), .ZN(n100) );
  AOI22D1BWP30P140LVT U128 ( .A1(n207), .A2(i_data_bus[102]), .B1(n1), .B2(
        i_data_bus[134]), .ZN(n99) );
  ND3D1BWP30P140LVT U129 ( .A1(n101), .A2(n100), .A3(n99), .ZN(N375) );
  AOI22D1BWP30P140LVT U130 ( .A1(n4), .A2(i_data_bus[197]), .B1(n3), .B2(
        i_data_bus[165]), .ZN(n102) );
  IOA21D1BWP30P140LVT U131 ( .A1(n2), .A2(i_data_bus[229]), .B(n102), .ZN(n103) );
  AOI21D1BWP30P140LVT U132 ( .A1(n5), .A2(i_data_bus[5]), .B(n103), .ZN(n106)
         );
  AOI22D1BWP30P140LVT U133 ( .A1(n206), .A2(i_data_bus[69]), .B1(n205), .B2(
        i_data_bus[37]), .ZN(n105) );
  AOI22D1BWP30P140LVT U134 ( .A1(n207), .A2(i_data_bus[101]), .B1(n1), .B2(
        i_data_bus[133]), .ZN(n104) );
  ND3D1BWP30P140LVT U135 ( .A1(n106), .A2(n105), .A3(n104), .ZN(N374) );
  AOI22D1BWP30P140LVT U136 ( .A1(n4), .A2(i_data_bus[203]), .B1(n3), .B2(
        i_data_bus[171]), .ZN(n107) );
  IOA21D1BWP30P140LVT U137 ( .A1(n2), .A2(i_data_bus[235]), .B(n107), .ZN(n108) );
  AOI21D1BWP30P140LVT U138 ( .A1(n220), .A2(i_data_bus[11]), .B(n108), .ZN(
        n111) );
  AOI22D1BWP30P140LVT U139 ( .A1(n206), .A2(i_data_bus[75]), .B1(n205), .B2(
        i_data_bus[43]), .ZN(n110) );
  AOI22D1BWP30P140LVT U140 ( .A1(n207), .A2(i_data_bus[107]), .B1(n1), .B2(
        i_data_bus[139]), .ZN(n109) );
  ND3D1BWP30P140LVT U141 ( .A1(n111), .A2(n110), .A3(n109), .ZN(N380) );
  AOI22D1BWP30P140LVT U142 ( .A1(n4), .A2(i_data_bus[202]), .B1(n3), .B2(
        i_data_bus[170]), .ZN(n112) );
  IOA21D1BWP30P140LVT U143 ( .A1(n2), .A2(i_data_bus[234]), .B(n112), .ZN(n113) );
  AOI21D1BWP30P140LVT U144 ( .A1(n5), .A2(i_data_bus[10]), .B(n113), .ZN(n116)
         );
  AOI22D1BWP30P140LVT U145 ( .A1(n206), .A2(i_data_bus[74]), .B1(n205), .B2(
        i_data_bus[42]), .ZN(n115) );
  AOI22D1BWP30P140LVT U146 ( .A1(n207), .A2(i_data_bus[106]), .B1(n1), .B2(
        i_data_bus[138]), .ZN(n114) );
  ND3D1BWP30P140LVT U147 ( .A1(n116), .A2(n115), .A3(n114), .ZN(N379) );
  AOI22D1BWP30P140LVT U148 ( .A1(n4), .A2(i_data_bus[201]), .B1(n3), .B2(
        i_data_bus[169]), .ZN(n117) );
  IOA21D1BWP30P140LVT U149 ( .A1(n2), .A2(i_data_bus[233]), .B(n117), .ZN(n118) );
  AOI21D1BWP30P140LVT U150 ( .A1(n5), .A2(i_data_bus[9]), .B(n118), .ZN(n121)
         );
  AOI22D1BWP30P140LVT U151 ( .A1(n206), .A2(i_data_bus[73]), .B1(n205), .B2(
        i_data_bus[41]), .ZN(n120) );
  AOI22D1BWP30P140LVT U152 ( .A1(n207), .A2(i_data_bus[105]), .B1(n1), .B2(
        i_data_bus[137]), .ZN(n119) );
  ND3D1BWP30P140LVT U153 ( .A1(n121), .A2(n120), .A3(n119), .ZN(N378) );
  AOI22D1BWP30P140LVT U154 ( .A1(n4), .A2(i_data_bus[204]), .B1(n3), .B2(
        i_data_bus[172]), .ZN(n122) );
  IOA21D1BWP30P140LVT U155 ( .A1(n2), .A2(i_data_bus[236]), .B(n122), .ZN(n123) );
  AOI21D1BWP30P140LVT U156 ( .A1(n220), .A2(i_data_bus[12]), .B(n123), .ZN(
        n126) );
  AOI22D1BWP30P140LVT U157 ( .A1(n206), .A2(i_data_bus[76]), .B1(n205), .B2(
        i_data_bus[44]), .ZN(n125) );
  AOI22D1BWP30P140LVT U158 ( .A1(n207), .A2(i_data_bus[108]), .B1(n1), .B2(
        i_data_bus[140]), .ZN(n124) );
  ND3D1BWP30P140LVT U159 ( .A1(n126), .A2(n125), .A3(n124), .ZN(N381) );
  AOI22D1BWP30P140LVT U160 ( .A1(n4), .A2(i_data_bus[216]), .B1(n3), .B2(
        i_data_bus[184]), .ZN(n127) );
  IOA21D1BWP30P140LVT U161 ( .A1(n2), .A2(i_data_bus[248]), .B(n127), .ZN(n128) );
  AOI21D1BWP30P140LVT U162 ( .A1(n5), .A2(i_data_bus[24]), .B(n128), .ZN(n132)
         );
  AOI22D1BWP30P140LVT U163 ( .A1(n222), .A2(i_data_bus[88]), .B1(n221), .B2(
        i_data_bus[56]), .ZN(n131) );
  AOI22D1BWP30P140LVT U164 ( .A1(n233), .A2(i_data_bus[120]), .B1(n1), .B2(
        i_data_bus[152]), .ZN(n130) );
  ND3D1BWP30P140LVT U165 ( .A1(n132), .A2(n131), .A3(n130), .ZN(N393) );
  AOI22D1BWP30P140LVT U166 ( .A1(n4), .A2(i_data_bus[209]), .B1(n3), .B2(
        i_data_bus[177]), .ZN(n133) );
  IOA21D1BWP30P140LVT U167 ( .A1(n2), .A2(i_data_bus[241]), .B(n133), .ZN(n134) );
  AOI21D1BWP30P140LVT U168 ( .A1(n5), .A2(i_data_bus[17]), .B(n134), .ZN(n137)
         );
  AOI22D1BWP30P140LVT U169 ( .A1(n222), .A2(i_data_bus[81]), .B1(n221), .B2(
        i_data_bus[49]), .ZN(n136) );
  AOI22D1BWP30P140LVT U170 ( .A1(n233), .A2(i_data_bus[113]), .B1(n1), .B2(
        i_data_bus[145]), .ZN(n135) );
  ND3D1BWP30P140LVT U171 ( .A1(n137), .A2(n136), .A3(n135), .ZN(N386) );
  AOI22D1BWP30P140LVT U172 ( .A1(n4), .A2(i_data_bus[215]), .B1(n3), .B2(
        i_data_bus[183]), .ZN(n138) );
  IOA21D1BWP30P140LVT U173 ( .A1(n2), .A2(i_data_bus[247]), .B(n138), .ZN(n139) );
  AOI21D1BWP30P140LVT U174 ( .A1(n220), .A2(i_data_bus[23]), .B(n139), .ZN(
        n142) );
  AOI22D1BWP30P140LVT U175 ( .A1(n222), .A2(i_data_bus[87]), .B1(n221), .B2(
        i_data_bus[55]), .ZN(n141) );
  AOI22D1BWP30P140LVT U176 ( .A1(n233), .A2(i_data_bus[119]), .B1(n1), .B2(
        i_data_bus[151]), .ZN(n140) );
  ND3D1BWP30P140LVT U177 ( .A1(n142), .A2(n141), .A3(n140), .ZN(N392) );
  AOI22D1BWP30P140LVT U178 ( .A1(n4), .A2(i_data_bus[214]), .B1(n3), .B2(
        i_data_bus[182]), .ZN(n143) );
  IOA21D1BWP30P140LVT U179 ( .A1(n2), .A2(i_data_bus[246]), .B(n143), .ZN(n144) );
  AOI21D1BWP30P140LVT U180 ( .A1(n5), .A2(i_data_bus[22]), .B(n144), .ZN(n147)
         );
  AOI22D1BWP30P140LVT U181 ( .A1(n222), .A2(i_data_bus[86]), .B1(n221), .B2(
        i_data_bus[54]), .ZN(n146) );
  AOI22D1BWP30P140LVT U182 ( .A1(n233), .A2(i_data_bus[118]), .B1(n1), .B2(
        i_data_bus[150]), .ZN(n145) );
  ND3D1BWP30P140LVT U183 ( .A1(n147), .A2(n146), .A3(n145), .ZN(N391) );
  AOI22D1BWP30P140LVT U184 ( .A1(n4), .A2(i_data_bus[213]), .B1(n3), .B2(
        i_data_bus[181]), .ZN(n148) );
  IOA21D1BWP30P140LVT U185 ( .A1(n2), .A2(i_data_bus[245]), .B(n148), .ZN(n149) );
  AOI21D1BWP30P140LVT U186 ( .A1(n5), .A2(i_data_bus[21]), .B(n149), .ZN(n152)
         );
  AOI22D1BWP30P140LVT U187 ( .A1(n222), .A2(i_data_bus[85]), .B1(n221), .B2(
        i_data_bus[53]), .ZN(n151) );
  AOI22D1BWP30P140LVT U188 ( .A1(n233), .A2(i_data_bus[117]), .B1(n1), .B2(
        i_data_bus[149]), .ZN(n150) );
  ND3D1BWP30P140LVT U189 ( .A1(n152), .A2(n151), .A3(n150), .ZN(N390) );
  AOI22D1BWP30P140LVT U190 ( .A1(n4), .A2(i_data_bus[212]), .B1(n3), .B2(
        i_data_bus[180]), .ZN(n153) );
  IOA21D1BWP30P140LVT U191 ( .A1(n2), .A2(i_data_bus[244]), .B(n153), .ZN(n154) );
  AOI21D1BWP30P140LVT U192 ( .A1(n220), .A2(i_data_bus[20]), .B(n154), .ZN(
        n157) );
  AOI22D1BWP30P140LVT U193 ( .A1(n222), .A2(i_data_bus[84]), .B1(n221), .B2(
        i_data_bus[52]), .ZN(n156) );
  AOI22D1BWP30P140LVT U194 ( .A1(n233), .A2(i_data_bus[116]), .B1(n1), .B2(
        i_data_bus[148]), .ZN(n155) );
  ND3D1BWP30P140LVT U195 ( .A1(n157), .A2(n156), .A3(n155), .ZN(N389) );
  AOI22D1BWP30P140LVT U196 ( .A1(n4), .A2(i_data_bus[211]), .B1(n3), .B2(
        i_data_bus[179]), .ZN(n158) );
  IOA21D1BWP30P140LVT U197 ( .A1(n2), .A2(i_data_bus[243]), .B(n158), .ZN(n159) );
  AOI21D1BWP30P140LVT U198 ( .A1(n5), .A2(i_data_bus[19]), .B(n159), .ZN(n162)
         );
  AOI22D1BWP30P140LVT U199 ( .A1(n222), .A2(i_data_bus[83]), .B1(n221), .B2(
        i_data_bus[51]), .ZN(n161) );
  AOI22D1BWP30P140LVT U200 ( .A1(n233), .A2(i_data_bus[115]), .B1(n1), .B2(
        i_data_bus[147]), .ZN(n160) );
  ND3D1BWP30P140LVT U201 ( .A1(n162), .A2(n161), .A3(n160), .ZN(N388) );
  AOI22D1BWP30P140LVT U202 ( .A1(n4), .A2(i_data_bus[210]), .B1(n3), .B2(
        i_data_bus[178]), .ZN(n163) );
  IOA21D1BWP30P140LVT U203 ( .A1(n2), .A2(i_data_bus[242]), .B(n163), .ZN(n164) );
  AOI21D1BWP30P140LVT U204 ( .A1(n5), .A2(i_data_bus[18]), .B(n164), .ZN(n167)
         );
  AOI22D1BWP30P140LVT U205 ( .A1(n222), .A2(i_data_bus[82]), .B1(n221), .B2(
        i_data_bus[50]), .ZN(n166) );
  AOI22D1BWP30P140LVT U206 ( .A1(n233), .A2(i_data_bus[114]), .B1(n1), .B2(
        i_data_bus[146]), .ZN(n165) );
  ND3D1BWP30P140LVT U207 ( .A1(n167), .A2(n166), .A3(n165), .ZN(N387) );
  AOI22D1BWP30P140LVT U208 ( .A1(n4), .A2(i_data_bus[206]), .B1(n3), .B2(
        i_data_bus[174]), .ZN(n168) );
  IOA21D1BWP30P140LVT U209 ( .A1(n2), .A2(i_data_bus[238]), .B(n168), .ZN(n169) );
  AOI22D1BWP30P140LVT U210 ( .A1(n222), .A2(i_data_bus[78]), .B1(n221), .B2(
        i_data_bus[46]), .ZN(n171) );
  AOI22D1BWP30P140LVT U211 ( .A1(n233), .A2(i_data_bus[110]), .B1(n1), .B2(
        i_data_bus[142]), .ZN(n170) );
  ND3D1BWP30P140LVT U212 ( .A1(n172), .A2(n171), .A3(n170), .ZN(N383) );
  INVD1BWP30P140LVT U213 ( .I(i_data_bus[173]), .ZN(n173) );
  MAOI22D1BWP30P140LVT U214 ( .A1(n4), .A2(i_data_bus[205]), .B1(n174), .B2(
        n173), .ZN(n175) );
  IOA21D1BWP30P140LVT U215 ( .A1(n2), .A2(i_data_bus[237]), .B(n175), .ZN(n176) );
  AOI21D1BWP30P140LVT U216 ( .A1(n220), .A2(i_data_bus[13]), .B(n176), .ZN(
        n179) );
  AOI22D1BWP30P140LVT U217 ( .A1(n222), .A2(i_data_bus[77]), .B1(n221), .B2(
        i_data_bus[45]), .ZN(n178) );
  AOI22D1BWP30P140LVT U218 ( .A1(n233), .A2(i_data_bus[109]), .B1(n1), .B2(
        i_data_bus[141]), .ZN(n177) );
  ND3D1BWP30P140LVT U219 ( .A1(n179), .A2(n178), .A3(n177), .ZN(N382) );
  INVD1BWP30P140LVT U220 ( .I(i_data_bus[194]), .ZN(n180) );
  MAOI22D1BWP30P140LVT U221 ( .A1(n3), .A2(i_data_bus[162]), .B1(n212), .B2(
        n180), .ZN(n181) );
  IOA21D1BWP30P140LVT U222 ( .A1(n2), .A2(i_data_bus[226]), .B(n181), .ZN(n182) );
  AOI21D1BWP30P140LVT U223 ( .A1(n5), .A2(i_data_bus[2]), .B(n182), .ZN(n185)
         );
  AOI22D1BWP30P140LVT U224 ( .A1(n206), .A2(i_data_bus[66]), .B1(n205), .B2(
        i_data_bus[34]), .ZN(n184) );
  AOI22D1BWP30P140LVT U225 ( .A1(n207), .A2(i_data_bus[98]), .B1(n1), .B2(
        i_data_bus[130]), .ZN(n183) );
  ND3D1BWP30P140LVT U226 ( .A1(n185), .A2(n184), .A3(n183), .ZN(N371) );
  INVD1BWP30P140LVT U227 ( .I(n2), .ZN(n192) );
  INVD1BWP30P140LVT U228 ( .I(i_data_bus[224]), .ZN(n191) );
  INVD1BWP30P140LVT U229 ( .I(i_data_bus[192]), .ZN(n186) );
  MAOI22D1BWP30P140LVT U230 ( .A1(n3), .A2(i_data_bus[160]), .B1(n212), .B2(
        n186), .ZN(n190) );
  INR2D1BWP30P140LVT U231 ( .A1(i_data_bus[0]), .B1(n187), .ZN(n188) );
  INVD1BWP30P140LVT U232 ( .I(n188), .ZN(n189) );
  OA211D1BWP30P140LVT U233 ( .A1(n192), .A2(n191), .B(n190), .C(n189), .Z(n195) );
  AOI22D1BWP30P140LVT U234 ( .A1(n206), .A2(i_data_bus[64]), .B1(n205), .B2(
        i_data_bus[32]), .ZN(n194) );
  AOI22D1BWP30P140LVT U235 ( .A1(n207), .A2(i_data_bus[96]), .B1(n1), .B2(
        i_data_bus[128]), .ZN(n193) );
  ND3D1BWP30P140LVT U236 ( .A1(n195), .A2(n194), .A3(n193), .ZN(N369) );
  INVD1BWP30P140LVT U237 ( .I(i_data_bus[193]), .ZN(n196) );
  MAOI22D1BWP30P140LVT U238 ( .A1(n3), .A2(i_data_bus[161]), .B1(n212), .B2(
        n196), .ZN(n197) );
  IOA21D1BWP30P140LVT U239 ( .A1(n2), .A2(i_data_bus[225]), .B(n197), .ZN(n198) );
  AOI21D1BWP30P140LVT U240 ( .A1(n220), .A2(i_data_bus[1]), .B(n198), .ZN(n201) );
  AOI22D1BWP30P140LVT U241 ( .A1(n206), .A2(i_data_bus[65]), .B1(n205), .B2(
        i_data_bus[33]), .ZN(n200) );
  AOI22D1BWP30P140LVT U242 ( .A1(n207), .A2(i_data_bus[97]), .B1(n1), .B2(
        i_data_bus[129]), .ZN(n199) );
  ND3D1BWP30P140LVT U243 ( .A1(n201), .A2(n200), .A3(n199), .ZN(N370) );
  INVD1BWP30P140LVT U244 ( .I(i_data_bus[195]), .ZN(n202) );
  MAOI22D1BWP30P140LVT U245 ( .A1(n3), .A2(i_data_bus[163]), .B1(n212), .B2(
        n202), .ZN(n203) );
  IOA21D1BWP30P140LVT U246 ( .A1(n2), .A2(i_data_bus[227]), .B(n203), .ZN(n204) );
  AOI21D1BWP30P140LVT U247 ( .A1(n5), .A2(i_data_bus[3]), .B(n204), .ZN(n210)
         );
  AOI22D1BWP30P140LVT U248 ( .A1(n206), .A2(i_data_bus[67]), .B1(n205), .B2(
        i_data_bus[35]), .ZN(n209) );
  AOI22D1BWP30P140LVT U249 ( .A1(n207), .A2(i_data_bus[99]), .B1(n1), .B2(
        i_data_bus[131]), .ZN(n208) );
  ND3D1BWP30P140LVT U250 ( .A1(n210), .A2(n209), .A3(n208), .ZN(N372) );
  INVD1BWP30P140LVT U251 ( .I(i_data_bus[208]), .ZN(n211) );
  MAOI22D1BWP30P140LVT U252 ( .A1(n3), .A2(i_data_bus[176]), .B1(n212), .B2(
        n211), .ZN(n213) );
  IOA21D1BWP30P140LVT U253 ( .A1(n2), .A2(i_data_bus[240]), .B(n213), .ZN(n214) );
  AOI21D1BWP30P140LVT U254 ( .A1(n5), .A2(i_data_bus[16]), .B(n214), .ZN(n217)
         );
  AOI22D1BWP30P140LVT U255 ( .A1(n222), .A2(i_data_bus[80]), .B1(n221), .B2(
        i_data_bus[48]), .ZN(n216) );
  AOI22D1BWP30P140LVT U256 ( .A1(n233), .A2(i_data_bus[112]), .B1(n1), .B2(
        i_data_bus[144]), .ZN(n215) );
  ND3D1BWP30P140LVT U257 ( .A1(n217), .A2(n216), .A3(n215), .ZN(N385) );
  AOI22D1BWP30P140LVT U258 ( .A1(n4), .A2(i_data_bus[217]), .B1(n3), .B2(
        i_data_bus[185]), .ZN(n218) );
  IOA21D1BWP30P140LVT U259 ( .A1(n2), .A2(i_data_bus[249]), .B(n218), .ZN(n219) );
  AOI21D1BWP30P140LVT U260 ( .A1(n5), .A2(i_data_bus[25]), .B(n219), .ZN(n225)
         );
  AOI22D1BWP30P140LVT U261 ( .A1(n222), .A2(i_data_bus[89]), .B1(n221), .B2(
        i_data_bus[57]), .ZN(n224) );
  AOI22D1BWP30P140LVT U262 ( .A1(n233), .A2(i_data_bus[121]), .B1(n1), .B2(
        i_data_bus[153]), .ZN(n223) );
  ND3D1BWP30P140LVT U263 ( .A1(n225), .A2(n224), .A3(n223), .ZN(N394) );
  AOI22D1BWP30P140LVT U264 ( .A1(n4), .A2(i_data_bus[207]), .B1(n3), .B2(
        i_data_bus[175]), .ZN(n226) );
  IOA21D1BWP30P140LVT U265 ( .A1(n2), .A2(i_data_bus[239]), .B(n226), .ZN(n228) );
  AOI21D1BWP30P140LVT U266 ( .A1(n5), .A2(i_data_bus[15]), .B(n228), .ZN(n236)
         );
  INVD1BWP30P140LVT U267 ( .I(i_data_bus[79]), .ZN(n231) );
  INVD1BWP30P140LVT U268 ( .I(i_data_bus[47]), .ZN(n229) );
  OA22D1BWP30P140LVT U269 ( .A1(n232), .A2(n231), .B1(n230), .B2(n229), .Z(
        n235) );
  AOI22D1BWP30P140LVT U270 ( .A1(n233), .A2(i_data_bus[111]), .B1(n1), .B2(
        i_data_bus[143]), .ZN(n234) );
  ND3D1BWP30P140LVT U271 ( .A1(n236), .A2(n235), .A3(n234), .ZN(N384) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_5 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD3BWP30P140LVT U3 ( .I(n184), .ZN(n234) );
  CKND2D2BWP30P140LVT U4 ( .A1(n5), .A2(n4), .ZN(n22) );
  NR2D2BWP30P140LVT U5 ( .A1(i_cmd[7]), .A2(i_cmd[6]), .ZN(n5) );
  OR2D1BWP30P140LVT U6 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n26) );
  IAO21D1BWP30P140LVT U7 ( .A1(n137), .A2(n1), .B(n125), .ZN(n128) );
  INVD1BWP30P140LVT U8 ( .I(i_data_bus[14]), .ZN(n1) );
  INVD1BWP30P140LVT U9 ( .I(n137), .ZN(n233) );
  INVD2BWP30P140LVT U10 ( .I(n186), .ZN(n164) );
  INVD2BWP30P140LVT U11 ( .I(n100), .ZN(n186) );
  NR2D3BWP30P140LVT U12 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n13) );
  BUFFD2BWP30P140LVT U13 ( .I(n52), .Z(n229) );
  INR2D1BWP30P140LVT U14 ( .A1(i_en), .B1(rst), .ZN(n3) );
  NR4D0BWP30P140LVT U15 ( .A1(n17), .A2(n16), .A3(i_cmd[5]), .A4(i_cmd[7]), 
        .ZN(n18) );
  INVD1BWP30P140LVT U16 ( .I(i_valid[6]), .ZN(n16) );
  INVD1BWP30P140LVT U17 ( .I(n34), .ZN(n78) );
  INVD1BWP30P140LVT U18 ( .I(n186), .ZN(n235) );
  INVD1BWP30P140LVT U19 ( .I(n78), .ZN(n237) );
  INVD1BWP30P140LVT U20 ( .I(i_cmd[5]), .ZN(n19) );
  NR2OPTPAD1BWP30P140LVT U21 ( .A1(n6), .A2(n22), .ZN(n37) );
  INVD1BWP30P140LVT U22 ( .I(n231), .ZN(n142) );
  INR2D1BWP30P140LVT U23 ( .A1(n33), .B1(n28), .ZN(n163) );
  INVD1BWP30P140LVT U24 ( .I(n79), .ZN(n165) );
  INR2D1BWP30P140LVT U25 ( .A1(n33), .B1(n25), .ZN(n100) );
  INVD1BWP30P140LVT U26 ( .I(n163), .ZN(n184) );
  INVD1BWP30P140LVT U27 ( .I(n78), .ZN(n224) );
  ND2D1BWP30P140LVT U28 ( .A1(n175), .A2(n174), .ZN(n176) );
  ND2D1BWP30P140LVT U29 ( .A1(n228), .A2(i_data_bus[185]), .ZN(n175) );
  AOI22D1BWP30P140LVT U30 ( .A1(n229), .A2(i_data_bus[217]), .B1(
        i_data_bus[249]), .B2(n231), .ZN(n174) );
  NR4D0BWP30P140LVT U31 ( .A1(n9), .A2(n8), .A3(i_cmd[6]), .A4(i_cmd[5]), .ZN(
        n15) );
  INVD1BWP30P140LVT U32 ( .I(i_valid[7]), .ZN(n9) );
  INVD1BWP30P140LVT U33 ( .I(i_cmd[7]), .ZN(n8) );
  NR2D1BWP30P140LVT U34 ( .A1(n164), .A2(n234), .ZN(n39) );
  NR2D1BWP30P140LVT U35 ( .A1(n237), .A2(n236), .ZN(n38) );
  INVD1BWP30P140LVT U36 ( .I(i_cmd[3]), .ZN(n30) );
  OR2D4BWP30P140LVT U37 ( .A1(n29), .A2(n14), .Z(n20) );
  INR2D1BWP30P140LVT U38 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n2) );
  INVD1BWP30P140LVT U39 ( .I(n2), .ZN(n7) );
  OR2D1BWP30P140LVT U40 ( .A1(n26), .A2(i_cmd[1]), .Z(n6) );
  INR2D2BWP30P140LVT U41 ( .A1(n3), .B1(i_cmd[5]), .ZN(n4) );
  IND3D2BWP30P140LVT U42 ( .A1(n7), .B1(i_cmd[0]), .B2(n37), .ZN(n137) );
  INVD1BWP30P140LVT U43 ( .I(i_cmd[2]), .ZN(n10) );
  INVD2BWP30P140LVT U44 ( .I(i_cmd[1]), .ZN(n24) );
  ND2OPTIBD2BWP30P140LVT U45 ( .A1(n10), .A2(n24), .ZN(n29) );
  INR2D1BWP30P140LVT U46 ( .A1(i_en), .B1(rst), .ZN(n11) );
  INR2D4BWP30P140LVT U47 ( .A1(n11), .B1(i_cmd[3]), .ZN(n12) );
  ND2OPTPAD2BWP30P140LVT U48 ( .A1(n13), .A2(n12), .ZN(n14) );
  INR2D4BWP30P140LVT U49 ( .A1(n15), .B1(n20), .ZN(n231) );
  INVD1BWP30P140LVT U50 ( .I(i_cmd[6]), .ZN(n17) );
  INR2D2BWP30P140LVT U51 ( .A1(n18), .B1(n20), .ZN(n52) );
  INR4D1BWP30P140LVT U52 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n19), .ZN(n21) );
  INR2D1BWP30P140LVT U53 ( .A1(n21), .B1(n20), .ZN(n41) );
  INVD2BWP30P140LVT U54 ( .I(n41), .ZN(n130) );
  INVD4BWP30P140LVT U55 ( .I(n130), .ZN(n159) );
  NR4D0BWP30P140LVT U56 ( .A1(n162), .A2(n231), .A3(n229), .A4(n159), .ZN(n40)
         );
  NR2OPTPAD1BWP30P140LVT U57 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n23) );
  INR2D2BWP30P140LVT U58 ( .A1(n23), .B1(n22), .ZN(n33) );
  ND4D1BWP30P140LVT U59 ( .A1(n24), .A2(n30), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n25) );
  INVD1BWP30P140LVT U60 ( .I(n26), .ZN(n27) );
  ND3D1BWP30P140LVT U61 ( .A1(n27), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n28)
         );
  INVD1BWP30P140LVT U62 ( .I(n29), .ZN(n31) );
  ND3D1BWP30P140LVT U63 ( .A1(n31), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n32)
         );
  INR2D1BWP30P140LVT U64 ( .A1(n33), .B1(n32), .ZN(n34) );
  IND3D1BWP30P140LVT U65 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n35) );
  INVD1BWP30P140LVT U66 ( .I(n35), .ZN(n36) );
  ND2OPTIBD2BWP30P140LVT U67 ( .A1(n37), .A2(n36), .ZN(n79) );
  INVD2BWP30P140LVT U68 ( .I(n79), .ZN(n236) );
  ND3D1BWP30P140LVT U69 ( .A1(n40), .A2(n39), .A3(n38), .ZN(N402) );
  BUFFD4BWP30P140LVT U70 ( .I(n41), .Z(n228) );
  AOI22D1BWP30P140LVT U71 ( .A1(n229), .A2(i_data_bus[219]), .B1(n228), .B2(
        i_data_bus[187]), .ZN(n42) );
  IOA21D1BWP30P140LVT U72 ( .A1(n231), .A2(i_data_bus[251]), .B(n42), .ZN(n43)
         );
  AOI21D1BWP30P140LVT U73 ( .A1(n162), .A2(i_data_bus[27]), .B(n43), .ZN(n46)
         );
  AOI22D1BWP30P140LVT U74 ( .A1(n164), .A2(i_data_bus[91]), .B1(n234), .B2(
        i_data_bus[59]), .ZN(n45) );
  AOI22D1BWP30P140LVT U75 ( .A1(n237), .A2(i_data_bus[123]), .B1(n236), .B2(
        i_data_bus[155]), .ZN(n44) );
  ND3D1BWP30P140LVT U76 ( .A1(n46), .A2(n45), .A3(n44), .ZN(N396) );
  AOI22D1BWP30P140LVT U77 ( .A1(n229), .A2(i_data_bus[218]), .B1(n228), .B2(
        i_data_bus[186]), .ZN(n47) );
  IOA21D1BWP30P140LVT U78 ( .A1(n231), .A2(i_data_bus[250]), .B(n47), .ZN(n48)
         );
  AOI21D1BWP30P140LVT U79 ( .A1(n162), .A2(i_data_bus[26]), .B(n48), .ZN(n51)
         );
  AOI22D1BWP30P140LVT U80 ( .A1(n164), .A2(i_data_bus[90]), .B1(n234), .B2(
        i_data_bus[58]), .ZN(n50) );
  AOI22D1BWP30P140LVT U81 ( .A1(n237), .A2(i_data_bus[122]), .B1(n236), .B2(
        i_data_bus[154]), .ZN(n49) );
  ND3D1BWP30P140LVT U82 ( .A1(n51), .A2(n50), .A3(n49), .ZN(N395) );
  INVD2BWP30P140LVT U83 ( .I(n52), .ZN(n191) );
  INVD1BWP30P140LVT U84 ( .I(i_data_bus[223]), .ZN(n53) );
  MAOI22D1BWP30P140LVT U85 ( .A1(n159), .A2(i_data_bus[191]), .B1(n191), .B2(
        n53), .ZN(n54) );
  IOA21D1BWP30P140LVT U86 ( .A1(n231), .A2(i_data_bus[255]), .B(n54), .ZN(n55)
         );
  AOI21D1BWP30P140LVT U87 ( .A1(n162), .A2(i_data_bus[31]), .B(n55), .ZN(n58)
         );
  AOI22D1BWP30P140LVT U88 ( .A1(n164), .A2(i_data_bus[95]), .B1(n234), .B2(
        i_data_bus[63]), .ZN(n57) );
  AOI22D1BWP30P140LVT U89 ( .A1(n237), .A2(i_data_bus[127]), .B1(n236), .B2(
        i_data_bus[159]), .ZN(n56) );
  ND3D1BWP30P140LVT U90 ( .A1(n58), .A2(n57), .A3(n56), .ZN(N400) );
  INVD1BWP30P140LVT U91 ( .I(i_data_bus[222]), .ZN(n59) );
  MAOI22D1BWP30P140LVT U92 ( .A1(n159), .A2(i_data_bus[190]), .B1(n191), .B2(
        n59), .ZN(n60) );
  IOA21D1BWP30P140LVT U93 ( .A1(n231), .A2(i_data_bus[254]), .B(n60), .ZN(n61)
         );
  AOI21D1BWP30P140LVT U94 ( .A1(n162), .A2(i_data_bus[30]), .B(n61), .ZN(n64)
         );
  AOI22D1BWP30P140LVT U95 ( .A1(n164), .A2(i_data_bus[94]), .B1(n234), .B2(
        i_data_bus[62]), .ZN(n63) );
  AOI22D1BWP30P140LVT U96 ( .A1(n237), .A2(i_data_bus[126]), .B1(n236), .B2(
        i_data_bus[158]), .ZN(n62) );
  ND3D1BWP30P140LVT U97 ( .A1(n64), .A2(n63), .A3(n62), .ZN(N399) );
  AOI22D1BWP30P140LVT U98 ( .A1(n229), .A2(i_data_bus[220]), .B1(n228), .B2(
        i_data_bus[188]), .ZN(n65) );
  IOA21D1BWP30P140LVT U99 ( .A1(n231), .A2(i_data_bus[252]), .B(n65), .ZN(n66)
         );
  AOI21D1BWP30P140LVT U100 ( .A1(n162), .A2(i_data_bus[28]), .B(n66), .ZN(n69)
         );
  AOI22D1BWP30P140LVT U101 ( .A1(n164), .A2(i_data_bus[92]), .B1(n234), .B2(
        i_data_bus[60]), .ZN(n68) );
  AOI22D1BWP30P140LVT U102 ( .A1(n237), .A2(i_data_bus[124]), .B1(n236), .B2(
        i_data_bus[156]), .ZN(n67) );
  ND3D1BWP30P140LVT U103 ( .A1(n69), .A2(n68), .A3(n67), .ZN(N397) );
  INVD1BWP30P140LVT U104 ( .I(i_data_bus[221]), .ZN(n70) );
  MAOI22D1BWP30P140LVT U105 ( .A1(n159), .A2(i_data_bus[189]), .B1(n191), .B2(
        n70), .ZN(n71) );
  IOA21D1BWP30P140LVT U106 ( .A1(n231), .A2(i_data_bus[253]), .B(n71), .ZN(n72) );
  AOI21D1BWP30P140LVT U107 ( .A1(n162), .A2(i_data_bus[29]), .B(n72), .ZN(n75)
         );
  AOI22D1BWP30P140LVT U108 ( .A1(n164), .A2(i_data_bus[93]), .B1(n234), .B2(
        i_data_bus[61]), .ZN(n74) );
  AOI22D1BWP30P140LVT U109 ( .A1(n237), .A2(i_data_bus[125]), .B1(n236), .B2(
        i_data_bus[157]), .ZN(n73) );
  ND3D1BWP30P140LVT U110 ( .A1(n75), .A2(n74), .A3(n73), .ZN(N398) );
  INVD2BWP30P140LVT U111 ( .I(n137), .ZN(n162) );
  INVD2BWP30P140LVT U112 ( .I(n191), .ZN(n180) );
  AOI22D1BWP30P140LVT U113 ( .A1(n180), .A2(i_data_bus[201]), .B1(n159), .B2(
        i_data_bus[169]), .ZN(n76) );
  IOA21D1BWP30P140LVT U114 ( .A1(n231), .A2(i_data_bus[233]), .B(n76), .ZN(n77) );
  AOI21D1BWP30P140LVT U115 ( .A1(n162), .A2(i_data_bus[9]), .B(n77), .ZN(n82)
         );
  AOI22D1BWP30P140LVT U116 ( .A1(n164), .A2(i_data_bus[73]), .B1(n234), .B2(
        i_data_bus[41]), .ZN(n81) );
  AOI22D1BWP30P140LVT U117 ( .A1(n224), .A2(i_data_bus[105]), .B1(n165), .B2(
        i_data_bus[137]), .ZN(n80) );
  ND3D1BWP30P140LVT U118 ( .A1(n82), .A2(n81), .A3(n80), .ZN(N378) );
  AOI22D1BWP30P140LVT U119 ( .A1(n180), .A2(i_data_bus[202]), .B1(n159), .B2(
        i_data_bus[170]), .ZN(n83) );
  IOA21D1BWP30P140LVT U120 ( .A1(n231), .A2(i_data_bus[234]), .B(n83), .ZN(n84) );
  AOI21D1BWP30P140LVT U121 ( .A1(n162), .A2(i_data_bus[10]), .B(n84), .ZN(n87)
         );
  AOI22D1BWP30P140LVT U122 ( .A1(n235), .A2(i_data_bus[74]), .B1(n234), .B2(
        i_data_bus[42]), .ZN(n86) );
  AOI22D1BWP30P140LVT U123 ( .A1(n224), .A2(i_data_bus[106]), .B1(n165), .B2(
        i_data_bus[138]), .ZN(n85) );
  ND3D1BWP30P140LVT U124 ( .A1(n87), .A2(n86), .A3(n85), .ZN(N379) );
  AOI22D1BWP30P140LVT U125 ( .A1(n180), .A2(i_data_bus[196]), .B1(n159), .B2(
        i_data_bus[164]), .ZN(n88) );
  IOA21D1BWP30P140LVT U126 ( .A1(n231), .A2(i_data_bus[228]), .B(n88), .ZN(n89) );
  AOI21D1BWP30P140LVT U127 ( .A1(n162), .A2(i_data_bus[4]), .B(n89), .ZN(n92)
         );
  AOI22D1BWP30P140LVT U128 ( .A1(n164), .A2(i_data_bus[68]), .B1(n234), .B2(
        i_data_bus[36]), .ZN(n91) );
  AOI22D1BWP30P140LVT U129 ( .A1(n224), .A2(i_data_bus[100]), .B1(n165), .B2(
        i_data_bus[132]), .ZN(n90) );
  ND3D1BWP30P140LVT U130 ( .A1(n92), .A2(n91), .A3(n90), .ZN(N373) );
  AOI22D1BWP30P140LVT U131 ( .A1(n180), .A2(i_data_bus[200]), .B1(n159), .B2(
        i_data_bus[168]), .ZN(n93) );
  IOA21D1BWP30P140LVT U132 ( .A1(n231), .A2(i_data_bus[232]), .B(n93), .ZN(n94) );
  AOI21D1BWP30P140LVT U133 ( .A1(n162), .A2(i_data_bus[8]), .B(n94), .ZN(n97)
         );
  AOI22D1BWP30P140LVT U134 ( .A1(n235), .A2(i_data_bus[72]), .B1(n234), .B2(
        i_data_bus[40]), .ZN(n96) );
  AOI22D1BWP30P140LVT U135 ( .A1(n224), .A2(i_data_bus[104]), .B1(n165), .B2(
        i_data_bus[136]), .ZN(n95) );
  ND3D1BWP30P140LVT U136 ( .A1(n97), .A2(n96), .A3(n95), .ZN(N377) );
  AOI22D1BWP30P140LVT U137 ( .A1(n180), .A2(i_data_bus[204]), .B1(n159), .B2(
        i_data_bus[172]), .ZN(n98) );
  IOA21D1BWP30P140LVT U138 ( .A1(n231), .A2(i_data_bus[236]), .B(n98), .ZN(n99) );
  AOI21D1BWP30P140LVT U139 ( .A1(n162), .A2(i_data_bus[12]), .B(n99), .ZN(n103) );
  AOI22D1BWP30P140LVT U140 ( .A1(n100), .A2(i_data_bus[76]), .B1(n234), .B2(
        i_data_bus[44]), .ZN(n102) );
  AOI22D1BWP30P140LVT U141 ( .A1(n224), .A2(i_data_bus[108]), .B1(n165), .B2(
        i_data_bus[140]), .ZN(n101) );
  ND3D1BWP30P140LVT U142 ( .A1(n103), .A2(n102), .A3(n101), .ZN(N381) );
  AOI22D1BWP30P140LVT U143 ( .A1(n180), .A2(i_data_bus[203]), .B1(n159), .B2(
        i_data_bus[171]), .ZN(n104) );
  IOA21D1BWP30P140LVT U144 ( .A1(n231), .A2(i_data_bus[235]), .B(n104), .ZN(
        n105) );
  AOI21D1BWP30P140LVT U145 ( .A1(n162), .A2(i_data_bus[11]), .B(n105), .ZN(
        n108) );
  AOI22D1BWP30P140LVT U146 ( .A1(n164), .A2(i_data_bus[75]), .B1(n234), .B2(
        i_data_bus[43]), .ZN(n107) );
  AOI22D1BWP30P140LVT U147 ( .A1(n224), .A2(i_data_bus[107]), .B1(n165), .B2(
        i_data_bus[139]), .ZN(n106) );
  ND3D1BWP30P140LVT U148 ( .A1(n108), .A2(n107), .A3(n106), .ZN(N380) );
  AOI22D1BWP30P140LVT U149 ( .A1(n180), .A2(i_data_bus[197]), .B1(n159), .B2(
        i_data_bus[165]), .ZN(n109) );
  IOA21D1BWP30P140LVT U150 ( .A1(n231), .A2(i_data_bus[229]), .B(n109), .ZN(
        n110) );
  AOI21D1BWP30P140LVT U151 ( .A1(n162), .A2(i_data_bus[5]), .B(n110), .ZN(n113) );
  AOI22D1BWP30P140LVT U152 ( .A1(n164), .A2(i_data_bus[69]), .B1(n234), .B2(
        i_data_bus[37]), .ZN(n112) );
  AOI22D1BWP30P140LVT U153 ( .A1(n224), .A2(i_data_bus[101]), .B1(n165), .B2(
        i_data_bus[133]), .ZN(n111) );
  ND3D1BWP30P140LVT U154 ( .A1(n113), .A2(n112), .A3(n111), .ZN(N374) );
  AOI22D1BWP30P140LVT U155 ( .A1(n180), .A2(i_data_bus[199]), .B1(n159), .B2(
        i_data_bus[167]), .ZN(n114) );
  IOA21D1BWP30P140LVT U156 ( .A1(n231), .A2(i_data_bus[231]), .B(n114), .ZN(
        n115) );
  AOI21D1BWP30P140LVT U157 ( .A1(n162), .A2(i_data_bus[7]), .B(n115), .ZN(n118) );
  AOI22D1BWP30P140LVT U158 ( .A1(n164), .A2(i_data_bus[71]), .B1(n234), .B2(
        i_data_bus[39]), .ZN(n117) );
  AOI22D1BWP30P140LVT U159 ( .A1(n224), .A2(i_data_bus[103]), .B1(n165), .B2(
        i_data_bus[135]), .ZN(n116) );
  ND3D1BWP30P140LVT U160 ( .A1(n118), .A2(n117), .A3(n116), .ZN(N376) );
  AOI22D1BWP30P140LVT U161 ( .A1(n180), .A2(i_data_bus[198]), .B1(n159), .B2(
        i_data_bus[166]), .ZN(n119) );
  IOA21D1BWP30P140LVT U162 ( .A1(n231), .A2(i_data_bus[230]), .B(n119), .ZN(
        n120) );
  AOI21D1BWP30P140LVT U163 ( .A1(n162), .A2(i_data_bus[6]), .B(n120), .ZN(n123) );
  AOI22D1BWP30P140LVT U164 ( .A1(n164), .A2(i_data_bus[70]), .B1(n234), .B2(
        i_data_bus[38]), .ZN(n122) );
  AOI22D1BWP30P140LVT U165 ( .A1(n224), .A2(i_data_bus[102]), .B1(n165), .B2(
        i_data_bus[134]), .ZN(n121) );
  ND3D1BWP30P140LVT U166 ( .A1(n123), .A2(n122), .A3(n121), .ZN(N375) );
  AOI22D1BWP30P140LVT U167 ( .A1(n180), .A2(i_data_bus[206]), .B1(n159), .B2(
        i_data_bus[174]), .ZN(n124) );
  IOA21D1BWP30P140LVT U168 ( .A1(n231), .A2(i_data_bus[238]), .B(n124), .ZN(
        n125) );
  AOI22D1BWP30P140LVT U169 ( .A1(n235), .A2(i_data_bus[78]), .B1(n234), .B2(
        i_data_bus[46]), .ZN(n127) );
  AOI22D1BWP30P140LVT U170 ( .A1(n237), .A2(i_data_bus[110]), .B1(n236), .B2(
        i_data_bus[142]), .ZN(n126) );
  ND3D1BWP30P140LVT U171 ( .A1(n128), .A2(n127), .A3(n126), .ZN(N383) );
  INVD1BWP30P140LVT U172 ( .I(i_data_bus[173]), .ZN(n129) );
  MAOI22D1BWP30P140LVT U173 ( .A1(n180), .A2(i_data_bus[205]), .B1(n130), .B2(
        n129), .ZN(n131) );
  IOA21D1BWP30P140LVT U174 ( .A1(n231), .A2(i_data_bus[237]), .B(n131), .ZN(
        n132) );
  AOI21D1BWP30P140LVT U175 ( .A1(n233), .A2(i_data_bus[13]), .B(n132), .ZN(
        n135) );
  AOI22D1BWP30P140LVT U176 ( .A1(n235), .A2(i_data_bus[77]), .B1(n234), .B2(
        i_data_bus[45]), .ZN(n134) );
  AOI22D1BWP30P140LVT U177 ( .A1(n237), .A2(i_data_bus[109]), .B1(n236), .B2(
        i_data_bus[141]), .ZN(n133) );
  ND3D1BWP30P140LVT U178 ( .A1(n135), .A2(n134), .A3(n133), .ZN(N382) );
  INVD1BWP30P140LVT U179 ( .I(i_data_bus[224]), .ZN(n141) );
  INVD1BWP30P140LVT U180 ( .I(i_data_bus[192]), .ZN(n136) );
  MAOI22D1BWP30P140LVT U181 ( .A1(n228), .A2(i_data_bus[160]), .B1(n191), .B2(
        n136), .ZN(n140) );
  INR2D1BWP30P140LVT U182 ( .A1(i_data_bus[0]), .B1(n137), .ZN(n138) );
  INVD1BWP30P140LVT U183 ( .I(n138), .ZN(n139) );
  OA211D1BWP30P140LVT U184 ( .A1(n142), .A2(n141), .B(n140), .C(n139), .Z(n145) );
  AOI22D1BWP30P140LVT U185 ( .A1(n164), .A2(i_data_bus[64]), .B1(n234), .B2(
        i_data_bus[32]), .ZN(n144) );
  AOI22D1BWP30P140LVT U186 ( .A1(n224), .A2(i_data_bus[96]), .B1(n165), .B2(
        i_data_bus[128]), .ZN(n143) );
  ND3D1BWP30P140LVT U187 ( .A1(n145), .A2(n144), .A3(n143), .ZN(N369) );
  INVD1BWP30P140LVT U188 ( .I(i_data_bus[193]), .ZN(n146) );
  MAOI22D1BWP30P140LVT U189 ( .A1(n159), .A2(i_data_bus[161]), .B1(n191), .B2(
        n146), .ZN(n147) );
  IOA21D1BWP30P140LVT U190 ( .A1(n231), .A2(i_data_bus[225]), .B(n147), .ZN(
        n148) );
  AOI21D1BWP30P140LVT U191 ( .A1(n162), .A2(i_data_bus[1]), .B(n148), .ZN(n151) );
  AOI22D1BWP30P140LVT U192 ( .A1(n164), .A2(i_data_bus[65]), .B1(n234), .B2(
        i_data_bus[33]), .ZN(n150) );
  AOI22D1BWP30P140LVT U193 ( .A1(n224), .A2(i_data_bus[97]), .B1(n165), .B2(
        i_data_bus[129]), .ZN(n149) );
  ND3D1BWP30P140LVT U194 ( .A1(n151), .A2(n150), .A3(n149), .ZN(N370) );
  INVD1BWP30P140LVT U195 ( .I(i_data_bus[194]), .ZN(n152) );
  MAOI22D1BWP30P140LVT U196 ( .A1(n159), .A2(i_data_bus[162]), .B1(n191), .B2(
        n152), .ZN(n153) );
  IOA21D1BWP30P140LVT U197 ( .A1(n231), .A2(i_data_bus[226]), .B(n153), .ZN(
        n154) );
  AOI21D1BWP30P140LVT U198 ( .A1(n162), .A2(i_data_bus[2]), .B(n154), .ZN(n157) );
  AOI22D1BWP30P140LVT U199 ( .A1(n235), .A2(i_data_bus[66]), .B1(n234), .B2(
        i_data_bus[34]), .ZN(n156) );
  AOI22D1BWP30P140LVT U200 ( .A1(n224), .A2(i_data_bus[98]), .B1(n165), .B2(
        i_data_bus[130]), .ZN(n155) );
  ND3D1BWP30P140LVT U201 ( .A1(n157), .A2(n156), .A3(n155), .ZN(N371) );
  INVD1BWP30P140LVT U202 ( .I(i_data_bus[195]), .ZN(n158) );
  MAOI22D1BWP30P140LVT U203 ( .A1(n159), .A2(i_data_bus[163]), .B1(n191), .B2(
        n158), .ZN(n160) );
  IOA21D1BWP30P140LVT U204 ( .A1(n231), .A2(i_data_bus[227]), .B(n160), .ZN(
        n161) );
  AOI21D1BWP30P140LVT U205 ( .A1(n162), .A2(i_data_bus[3]), .B(n161), .ZN(n168) );
  AOI22D1BWP30P140LVT U206 ( .A1(n164), .A2(i_data_bus[67]), .B1(n163), .B2(
        i_data_bus[35]), .ZN(n167) );
  AOI22D1BWP30P140LVT U207 ( .A1(n224), .A2(i_data_bus[99]), .B1(n165), .B2(
        i_data_bus[131]), .ZN(n166) );
  ND3D1BWP30P140LVT U208 ( .A1(n168), .A2(n167), .A3(n166), .ZN(N372) );
  AOI22D1BWP30P140LVT U209 ( .A1(n229), .A2(i_data_bus[216]), .B1(n228), .B2(
        i_data_bus[184]), .ZN(n169) );
  IOA21D1BWP30P140LVT U210 ( .A1(n231), .A2(i_data_bus[248]), .B(n169), .ZN(
        n170) );
  AOI21D1BWP30P140LVT U211 ( .A1(n233), .A2(i_data_bus[24]), .B(n170), .ZN(
        n173) );
  AOI22D1BWP30P140LVT U212 ( .A1(n235), .A2(i_data_bus[88]), .B1(n234), .B2(
        i_data_bus[56]), .ZN(n172) );
  AOI22D1BWP30P140LVT U213 ( .A1(n237), .A2(i_data_bus[120]), .B1(n236), .B2(
        i_data_bus[152]), .ZN(n171) );
  ND3D1BWP30P140LVT U214 ( .A1(n173), .A2(n172), .A3(n171), .ZN(N393) );
  AOI21D1BWP30P140LVT U215 ( .A1(n162), .A2(i_data_bus[25]), .B(n176), .ZN(
        n179) );
  AOI22D1BWP30P140LVT U216 ( .A1(n235), .A2(i_data_bus[89]), .B1(n234), .B2(
        i_data_bus[57]), .ZN(n178) );
  AOI22D1BWP30P140LVT U217 ( .A1(n237), .A2(i_data_bus[121]), .B1(n236), .B2(
        i_data_bus[153]), .ZN(n177) );
  ND3D1BWP30P140LVT U218 ( .A1(n179), .A2(n178), .A3(n177), .ZN(N394) );
  AOI22D1BWP30P140LVT U219 ( .A1(n180), .A2(i_data_bus[207]), .B1(n228), .B2(
        i_data_bus[175]), .ZN(n181) );
  IOA21D1BWP30P140LVT U220 ( .A1(n231), .A2(i_data_bus[239]), .B(n181), .ZN(
        n182) );
  AOI21D1BWP30P140LVT U221 ( .A1(n233), .A2(i_data_bus[15]), .B(n182), .ZN(
        n189) );
  INVD1BWP30P140LVT U222 ( .I(i_data_bus[79]), .ZN(n185) );
  INVD1BWP30P140LVT U223 ( .I(i_data_bus[47]), .ZN(n183) );
  OA22D1BWP30P140LVT U224 ( .A1(n186), .A2(n185), .B1(n184), .B2(n183), .Z(
        n188) );
  AOI22D1BWP30P140LVT U225 ( .A1(n237), .A2(i_data_bus[111]), .B1(n236), .B2(
        i_data_bus[143]), .ZN(n187) );
  ND3D1BWP30P140LVT U226 ( .A1(n189), .A2(n188), .A3(n187), .ZN(N384) );
  INVD1BWP30P140LVT U227 ( .I(i_data_bus[208]), .ZN(n190) );
  MAOI22D1BWP30P140LVT U228 ( .A1(n228), .A2(i_data_bus[176]), .B1(n191), .B2(
        n190), .ZN(n192) );
  IOA21D1BWP30P140LVT U229 ( .A1(n231), .A2(i_data_bus[240]), .B(n192), .ZN(
        n193) );
  AOI21D1BWP30P140LVT U230 ( .A1(n233), .A2(i_data_bus[16]), .B(n193), .ZN(
        n196) );
  AOI22D1BWP30P140LVT U231 ( .A1(n235), .A2(i_data_bus[80]), .B1(n234), .B2(
        i_data_bus[48]), .ZN(n195) );
  AOI22D1BWP30P140LVT U232 ( .A1(n237), .A2(i_data_bus[112]), .B1(n236), .B2(
        i_data_bus[144]), .ZN(n194) );
  ND3D1BWP30P140LVT U233 ( .A1(n196), .A2(n195), .A3(n194), .ZN(N385) );
  AOI22D1BWP30P140LVT U234 ( .A1(n229), .A2(i_data_bus[212]), .B1(n228), .B2(
        i_data_bus[180]), .ZN(n197) );
  IOA21D1BWP30P140LVT U235 ( .A1(n231), .A2(i_data_bus[244]), .B(n197), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U236 ( .A1(n233), .A2(i_data_bus[20]), .B(n198), .ZN(
        n201) );
  AOI22D1BWP30P140LVT U237 ( .A1(n235), .A2(i_data_bus[84]), .B1(n234), .B2(
        i_data_bus[52]), .ZN(n200) );
  AOI22D1BWP30P140LVT U238 ( .A1(n237), .A2(i_data_bus[116]), .B1(n236), .B2(
        i_data_bus[148]), .ZN(n199) );
  ND3D1BWP30P140LVT U239 ( .A1(n201), .A2(n200), .A3(n199), .ZN(N389) );
  AOI22D1BWP30P140LVT U240 ( .A1(n229), .A2(i_data_bus[209]), .B1(n228), .B2(
        i_data_bus[177]), .ZN(n202) );
  IOA21D1BWP30P140LVT U241 ( .A1(n231), .A2(i_data_bus[241]), .B(n202), .ZN(
        n203) );
  AOI21D1BWP30P140LVT U242 ( .A1(n233), .A2(i_data_bus[17]), .B(n203), .ZN(
        n206) );
  AOI22D1BWP30P140LVT U243 ( .A1(n235), .A2(i_data_bus[81]), .B1(n234), .B2(
        i_data_bus[49]), .ZN(n205) );
  AOI22D1BWP30P140LVT U244 ( .A1(n224), .A2(i_data_bus[113]), .B1(n236), .B2(
        i_data_bus[145]), .ZN(n204) );
  ND3D1BWP30P140LVT U245 ( .A1(n206), .A2(n205), .A3(n204), .ZN(N386) );
  AOI22D1BWP30P140LVT U246 ( .A1(n229), .A2(i_data_bus[211]), .B1(n228), .B2(
        i_data_bus[179]), .ZN(n207) );
  IOA21D1BWP30P140LVT U247 ( .A1(n231), .A2(i_data_bus[243]), .B(n207), .ZN(
        n208) );
  AOI21D1BWP30P140LVT U248 ( .A1(n233), .A2(i_data_bus[19]), .B(n208), .ZN(
        n211) );
  AOI22D1BWP30P140LVT U249 ( .A1(n235), .A2(i_data_bus[83]), .B1(n234), .B2(
        i_data_bus[51]), .ZN(n210) );
  AOI22D1BWP30P140LVT U250 ( .A1(n237), .A2(i_data_bus[115]), .B1(n236), .B2(
        i_data_bus[147]), .ZN(n209) );
  ND3D1BWP30P140LVT U251 ( .A1(n211), .A2(n210), .A3(n209), .ZN(N388) );
  AOI22D1BWP30P140LVT U252 ( .A1(n229), .A2(i_data_bus[213]), .B1(n228), .B2(
        i_data_bus[181]), .ZN(n212) );
  IOA21D1BWP30P140LVT U253 ( .A1(n231), .A2(i_data_bus[245]), .B(n212), .ZN(
        n213) );
  AOI21D1BWP30P140LVT U254 ( .A1(n233), .A2(i_data_bus[21]), .B(n213), .ZN(
        n216) );
  AOI22D1BWP30P140LVT U255 ( .A1(n235), .A2(i_data_bus[85]), .B1(n234), .B2(
        i_data_bus[53]), .ZN(n215) );
  AOI22D1BWP30P140LVT U256 ( .A1(n224), .A2(i_data_bus[117]), .B1(n236), .B2(
        i_data_bus[149]), .ZN(n214) );
  ND3D1BWP30P140LVT U257 ( .A1(n216), .A2(n215), .A3(n214), .ZN(N390) );
  AOI22D1BWP30P140LVT U258 ( .A1(n229), .A2(i_data_bus[214]), .B1(n228), .B2(
        i_data_bus[182]), .ZN(n217) );
  IOA21D1BWP30P140LVT U259 ( .A1(n231), .A2(i_data_bus[246]), .B(n217), .ZN(
        n218) );
  AOI21D1BWP30P140LVT U260 ( .A1(n233), .A2(i_data_bus[22]), .B(n218), .ZN(
        n221) );
  AOI22D1BWP30P140LVT U261 ( .A1(n235), .A2(i_data_bus[86]), .B1(n234), .B2(
        i_data_bus[54]), .ZN(n220) );
  AOI22D1BWP30P140LVT U262 ( .A1(n237), .A2(i_data_bus[118]), .B1(n236), .B2(
        i_data_bus[150]), .ZN(n219) );
  ND3D1BWP30P140LVT U263 ( .A1(n221), .A2(n220), .A3(n219), .ZN(N391) );
  AOI22D1BWP30P140LVT U264 ( .A1(n229), .A2(i_data_bus[215]), .B1(n228), .B2(
        i_data_bus[183]), .ZN(n222) );
  IOA21D1BWP30P140LVT U265 ( .A1(n231), .A2(i_data_bus[247]), .B(n222), .ZN(
        n223) );
  AOI21D1BWP30P140LVT U266 ( .A1(n233), .A2(i_data_bus[23]), .B(n223), .ZN(
        n227) );
  AOI22D1BWP30P140LVT U267 ( .A1(n235), .A2(i_data_bus[87]), .B1(n234), .B2(
        i_data_bus[55]), .ZN(n226) );
  AOI22D1BWP30P140LVT U268 ( .A1(n224), .A2(i_data_bus[119]), .B1(n236), .B2(
        i_data_bus[151]), .ZN(n225) );
  ND3D1BWP30P140LVT U269 ( .A1(n227), .A2(n226), .A3(n225), .ZN(N392) );
  AOI22D1BWP30P140LVT U270 ( .A1(n229), .A2(i_data_bus[210]), .B1(n228), .B2(
        i_data_bus[178]), .ZN(n230) );
  IOA21D1BWP30P140LVT U271 ( .A1(n231), .A2(i_data_bus[242]), .B(n230), .ZN(
        n232) );
  AOI21D1BWP30P140LVT U272 ( .A1(n233), .A2(i_data_bus[18]), .B(n232), .ZN(
        n240) );
  AOI22D1BWP30P140LVT U273 ( .A1(n235), .A2(i_data_bus[82]), .B1(n234), .B2(
        i_data_bus[50]), .ZN(n239) );
  AOI22D1BWP30P140LVT U274 ( .A1(n237), .A2(i_data_bus[114]), .B1(n236), .B2(
        i_data_bus[146]), .ZN(n238) );
  ND3D1BWP30P140LVT U275 ( .A1(n240), .A2(n239), .A3(n238), .ZN(N387) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_6 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD6BWP30P140LVT U3 ( .I(n229), .ZN(n2) );
  NR2OPTPAD1BWP30P140LVT U4 ( .A1(n6), .A2(n27), .ZN(n43) );
  NR2OPTPAD1BWP30P140LVT U5 ( .A1(i_cmd[0]), .A2(n15), .ZN(n16) );
  INR2D1BWP30P140LVT U6 ( .A1(n39), .B1(n34), .ZN(n35) );
  INVD8BWP30P140LVT U7 ( .I(n136), .ZN(n1) );
  INVD2BWP30P140LVT U8 ( .I(n161), .ZN(n3) );
  INVD3BWP30P140LVT U9 ( .I(n24), .ZN(n4) );
  INVD1BWP30P140LVT U10 ( .I(n131), .ZN(n78) );
  INVD2BWP30P140LVT U11 ( .I(n40), .ZN(n131) );
  IND3D6BWP30P140LVT U12 ( .A1(rst), .B1(n5), .B2(i_en), .ZN(n27) );
  NR3D4BWP30P140LVT U13 ( .A1(i_cmd[6]), .A2(i_cmd[5]), .A3(i_cmd[7]), .ZN(n5)
         );
  ND2OPTIBD1BWP30P140LVT U14 ( .A1(n13), .A2(n12), .ZN(n36) );
  INVD1BWP30P140LVT U15 ( .I(i_cmd[2]), .ZN(n13) );
  INVD1BWP30P140LVT U16 ( .I(i_cmd[1]), .ZN(n12) );
  ND2D1BWP30P140LVT U17 ( .A1(n43), .A2(n10), .ZN(n161) );
  NR2D1BWP30P140LVT U18 ( .A1(n9), .A2(n8), .ZN(n10) );
  INVD1BWP30P140LVT U19 ( .I(i_cmd[0]), .ZN(n8) );
  INVD1BWP30P140LVT U20 ( .I(n36), .ZN(n37) );
  ND2OPTIBD1BWP30P140LVT U21 ( .A1(n43), .A2(n42), .ZN(n84) );
  INVD1BWP30P140LVT U22 ( .I(n231), .ZN(n77) );
  INVD2BWP30P140LVT U23 ( .I(n84), .ZN(n232) );
  ND2D1BWP30P140LVT U24 ( .A1(n14), .A2(i_en), .ZN(n15) );
  NR2D1BWP30P140LVT U25 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n28) );
  OR2D2BWP30P140LVT U26 ( .A1(n36), .A2(n18), .Z(n24) );
  ND2OPTIBD1BWP30P140LVT U27 ( .A1(n17), .A2(n16), .ZN(n18) );
  MAOI22D1BWP30P140LVT U28 ( .A1(n1), .A2(i_data_bus[167]), .B1(n219), .B2(
        n123), .ZN(n124) );
  INVD1BWP30P140LVT U29 ( .I(i_data_bus[199]), .ZN(n123) );
  NR2D1BWP30P140LVT U30 ( .A1(n77), .A2(n2), .ZN(n45) );
  INVD4BWP30P140LVT U31 ( .I(n219), .ZN(n212) );
  INR2D4BWP30P140LVT U32 ( .A1(n19), .B1(n24), .ZN(n20) );
  ND2OPTIBD6BWP30P140LVT U33 ( .A1(n4), .A2(n23), .ZN(n219) );
  INVD1BWP30P140LVT U34 ( .I(n20), .ZN(n21) );
  OR2D1BWP30P140LVT U35 ( .A1(i_cmd[3]), .A2(i_cmd[2]), .Z(n32) );
  OR2D1BWP30P140LVT U36 ( .A1(n32), .A2(i_cmd[1]), .Z(n6) );
  INR2D1BWP30P140LVT U37 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n7) );
  INVD1BWP30P140LVT U38 ( .I(n7), .ZN(n9) );
  ND2D1BWP30P140LVT U39 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n11) );
  NR3D0P7BWP30P140LVT U40 ( .A1(n11), .A2(i_cmd[5]), .A3(i_cmd[6]), .ZN(n19)
         );
  NR2OPTPAD1BWP30P140LVT U41 ( .A1(i_cmd[3]), .A2(i_cmd[4]), .ZN(n17) );
  INVD1BWP30P140LVT U42 ( .I(rst), .ZN(n14) );
  INVD1BWP30P140LVT U43 ( .I(i_cmd[6]), .ZN(n22) );
  INR4D1BWP30P140LVT U44 ( .A1(i_valid[6]), .B1(i_cmd[5]), .B2(i_cmd[7]), .B3(
        n22), .ZN(n23) );
  INVD1BWP30P140LVT U45 ( .I(i_cmd[5]), .ZN(n25) );
  INR4D1BWP30P140LVT U46 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n25), .ZN(n26) );
  ND2OPTIBD4BWP30P140LVT U47 ( .A1(n4), .A2(n26), .ZN(n136) );
  NR4D0BWP30P140LVT U48 ( .A1(n3), .A2(n20), .A3(n212), .A4(n1), .ZN(n46) );
  INR2D2BWP30P140LVT U49 ( .A1(n28), .B1(n27), .ZN(n39) );
  INVD1BWP30P140LVT U50 ( .I(i_cmd[3]), .ZN(n29) );
  ND4D1BWP30P140LVT U51 ( .A1(n12), .A2(n29), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n30) );
  INR2D1BWP30P140LVT U52 ( .A1(n39), .B1(n30), .ZN(n31) );
  INVD2BWP30P140LVT U53 ( .I(n31), .ZN(n231) );
  INVD1BWP30P140LVT U54 ( .I(n32), .ZN(n33) );
  ND3D1BWP30P140LVT U55 ( .A1(n33), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n34)
         );
  INVD2BWP30P140LVT U56 ( .I(n35), .ZN(n229) );
  ND3D1BWP30P140LVT U57 ( .A1(n37), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n38)
         );
  INR2D1BWP30P140LVT U58 ( .A1(n39), .B1(n38), .ZN(n40) );
  IND3D1BWP30P140LVT U59 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n41) );
  INVD1BWP30P140LVT U60 ( .I(n41), .ZN(n42) );
  NR2D1BWP30P140LVT U61 ( .A1(n78), .A2(n232), .ZN(n44) );
  ND3D1BWP30P140LVT U62 ( .A1(n46), .A2(n45), .A3(n44), .ZN(N402) );
  AOI22D1BWP30P140LVT U63 ( .A1(n212), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n47) );
  IOA21D1BWP30P140LVT U64 ( .A1(n20), .A2(i_data_bus[252]), .B(n47), .ZN(n48)
         );
  AOI21D1BWP30P140LVT U65 ( .A1(n3), .A2(i_data_bus[28]), .B(n48), .ZN(n51) );
  AOI22D1BWP30P140LVT U66 ( .A1(n77), .A2(i_data_bus[92]), .B1(n2), .B2(
        i_data_bus[60]), .ZN(n50) );
  AOI22D1BWP30P140LVT U67 ( .A1(n78), .A2(i_data_bus[124]), .B1(n232), .B2(
        i_data_bus[156]), .ZN(n49) );
  ND3D1BWP30P140LVT U68 ( .A1(n51), .A2(n50), .A3(n49), .ZN(N397) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[221]), .ZN(n52) );
  MAOI22D1BWP30P140LVT U70 ( .A1(n1), .A2(i_data_bus[189]), .B1(n219), .B2(n52), .ZN(n53) );
  IOA21D1BWP30P140LVT U71 ( .A1(n20), .A2(i_data_bus[253]), .B(n53), .ZN(n54)
         );
  AOI21D1BWP30P140LVT U72 ( .A1(n3), .A2(i_data_bus[29]), .B(n54), .ZN(n57) );
  AOI22D1BWP30P140LVT U73 ( .A1(n77), .A2(i_data_bus[93]), .B1(n2), .B2(
        i_data_bus[61]), .ZN(n56) );
  AOI22D1BWP30P140LVT U74 ( .A1(n78), .A2(i_data_bus[125]), .B1(n232), .B2(
        i_data_bus[157]), .ZN(n55) );
  ND3D1BWP30P140LVT U75 ( .A1(n57), .A2(n56), .A3(n55), .ZN(N398) );
  INVD1BWP30P140LVT U76 ( .I(i_data_bus[222]), .ZN(n58) );
  MAOI22D1BWP30P140LVT U77 ( .A1(n1), .A2(i_data_bus[190]), .B1(n219), .B2(n58), .ZN(n59) );
  IOA21D1BWP30P140LVT U78 ( .A1(n20), .A2(i_data_bus[254]), .B(n59), .ZN(n60)
         );
  AOI21D1BWP30P140LVT U79 ( .A1(n3), .A2(i_data_bus[30]), .B(n60), .ZN(n63) );
  AOI22D1BWP30P140LVT U80 ( .A1(n77), .A2(i_data_bus[94]), .B1(n2), .B2(
        i_data_bus[62]), .ZN(n62) );
  AOI22D1BWP30P140LVT U81 ( .A1(n78), .A2(i_data_bus[126]), .B1(n232), .B2(
        i_data_bus[158]), .ZN(n61) );
  ND3D1BWP30P140LVT U82 ( .A1(n63), .A2(n62), .A3(n61), .ZN(N399) );
  INVD1BWP30P140LVT U83 ( .I(i_data_bus[223]), .ZN(n64) );
  MAOI22D1BWP30P140LVT U84 ( .A1(n1), .A2(i_data_bus[191]), .B1(n219), .B2(n64), .ZN(n65) );
  IOA21D1BWP30P140LVT U85 ( .A1(n20), .A2(i_data_bus[255]), .B(n65), .ZN(n66)
         );
  AOI21D1BWP30P140LVT U86 ( .A1(n3), .A2(i_data_bus[31]), .B(n66), .ZN(n69) );
  AOI22D1BWP30P140LVT U87 ( .A1(n77), .A2(i_data_bus[95]), .B1(n2), .B2(
        i_data_bus[63]), .ZN(n68) );
  AOI22D1BWP30P140LVT U88 ( .A1(n78), .A2(i_data_bus[127]), .B1(n232), .B2(
        i_data_bus[159]), .ZN(n67) );
  ND3D1BWP30P140LVT U89 ( .A1(n69), .A2(n68), .A3(n67), .ZN(N400) );
  AOI22D1BWP30P140LVT U90 ( .A1(n212), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n70) );
  IOA21D1BWP30P140LVT U91 ( .A1(n20), .A2(i_data_bus[251]), .B(n70), .ZN(n71)
         );
  AOI21D1BWP30P140LVT U92 ( .A1(n3), .A2(i_data_bus[27]), .B(n71), .ZN(n74) );
  AOI22D1BWP30P140LVT U93 ( .A1(n77), .A2(i_data_bus[91]), .B1(n2), .B2(
        i_data_bus[59]), .ZN(n73) );
  AOI22D1BWP30P140LVT U94 ( .A1(n78), .A2(i_data_bus[123]), .B1(n232), .B2(
        i_data_bus[155]), .ZN(n72) );
  ND3D1BWP30P140LVT U95 ( .A1(n74), .A2(n73), .A3(n72), .ZN(N396) );
  AOI22D1BWP30P140LVT U96 ( .A1(n212), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n75) );
  IOA21D1BWP30P140LVT U97 ( .A1(n20), .A2(i_data_bus[250]), .B(n75), .ZN(n76)
         );
  AOI21D1BWP30P140LVT U98 ( .A1(n3), .A2(i_data_bus[26]), .B(n76), .ZN(n81) );
  AOI22D1BWP30P140LVT U99 ( .A1(n77), .A2(i_data_bus[90]), .B1(n2), .B2(
        i_data_bus[58]), .ZN(n80) );
  AOI22D1BWP30P140LVT U100 ( .A1(n78), .A2(i_data_bus[122]), .B1(n232), .B2(
        i_data_bus[154]), .ZN(n79) );
  ND3D1BWP30P140LVT U101 ( .A1(n81), .A2(n80), .A3(n79), .ZN(N395) );
  AOI22D1BWP30P140LVT U102 ( .A1(n212), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n82) );
  IOA21D1BWP30P140LVT U103 ( .A1(n20), .A2(i_data_bus[236]), .B(n82), .ZN(n83)
         );
  AOI21D1BWP30P140LVT U104 ( .A1(n3), .A2(i_data_bus[12]), .B(n83), .ZN(n87)
         );
  INVD2BWP30P140LVT U105 ( .I(n231), .ZN(n166) );
  AOI22D1BWP30P140LVT U106 ( .A1(n166), .A2(i_data_bus[76]), .B1(n2), .B2(
        i_data_bus[44]), .ZN(n86) );
  INVD2BWP30P140LVT U107 ( .I(n131), .ZN(n168) );
  INVD2BWP30P140LVT U108 ( .I(n84), .ZN(n167) );
  AOI22D1BWP30P140LVT U109 ( .A1(n168), .A2(i_data_bus[108]), .B1(n167), .B2(
        i_data_bus[140]), .ZN(n85) );
  ND3D1BWP30P140LVT U110 ( .A1(n87), .A2(n86), .A3(n85), .ZN(N381) );
  AOI22D1BWP30P140LVT U111 ( .A1(n212), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n88) );
  IOA21D1BWP30P140LVT U112 ( .A1(n20), .A2(i_data_bus[233]), .B(n88), .ZN(n89)
         );
  AOI21D1BWP30P140LVT U113 ( .A1(n3), .A2(i_data_bus[9]), .B(n89), .ZN(n92) );
  AOI22D1BWP30P140LVT U114 ( .A1(n166), .A2(i_data_bus[73]), .B1(n2), .B2(
        i_data_bus[41]), .ZN(n91) );
  AOI22D1BWP30P140LVT U115 ( .A1(n168), .A2(i_data_bus[105]), .B1(n167), .B2(
        i_data_bus[137]), .ZN(n90) );
  ND3D1BWP30P140LVT U116 ( .A1(n92), .A2(n91), .A3(n90), .ZN(N378) );
  AOI22D1BWP30P140LVT U117 ( .A1(n212), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n93) );
  IOA21D1BWP30P140LVT U118 ( .A1(n20), .A2(i_data_bus[228]), .B(n93), .ZN(n94)
         );
  AOI21D1BWP30P140LVT U119 ( .A1(n3), .A2(i_data_bus[4]), .B(n94), .ZN(n97) );
  AOI22D1BWP30P140LVT U120 ( .A1(n166), .A2(i_data_bus[68]), .B1(n2), .B2(
        i_data_bus[36]), .ZN(n96) );
  AOI22D1BWP30P140LVT U121 ( .A1(n168), .A2(i_data_bus[100]), .B1(n167), .B2(
        i_data_bus[132]), .ZN(n95) );
  ND3D1BWP30P140LVT U122 ( .A1(n97), .A2(n96), .A3(n95), .ZN(N373) );
  AOI22D1BWP30P140LVT U123 ( .A1(n212), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n98) );
  IOA21D1BWP30P140LVT U124 ( .A1(n20), .A2(i_data_bus[235]), .B(n98), .ZN(n99)
         );
  AOI21D1BWP30P140LVT U125 ( .A1(n3), .A2(i_data_bus[11]), .B(n99), .ZN(n102)
         );
  AOI22D1BWP30P140LVT U126 ( .A1(n166), .A2(i_data_bus[75]), .B1(n2), .B2(
        i_data_bus[43]), .ZN(n101) );
  AOI22D1BWP30P140LVT U127 ( .A1(n168), .A2(i_data_bus[107]), .B1(n167), .B2(
        i_data_bus[139]), .ZN(n100) );
  ND3D1BWP30P140LVT U128 ( .A1(n102), .A2(n101), .A3(n100), .ZN(N380) );
  AOI22D1BWP30P140LVT U129 ( .A1(n212), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n103) );
  IOA21D1BWP30P140LVT U130 ( .A1(n20), .A2(i_data_bus[234]), .B(n103), .ZN(
        n104) );
  AOI21D1BWP30P140LVT U131 ( .A1(n3), .A2(i_data_bus[10]), .B(n104), .ZN(n107)
         );
  AOI22D1BWP30P140LVT U132 ( .A1(n166), .A2(i_data_bus[74]), .B1(n2), .B2(
        i_data_bus[42]), .ZN(n106) );
  AOI22D1BWP30P140LVT U133 ( .A1(n168), .A2(i_data_bus[106]), .B1(n167), .B2(
        i_data_bus[138]), .ZN(n105) );
  ND3D1BWP30P140LVT U134 ( .A1(n107), .A2(n106), .A3(n105), .ZN(N379) );
  AOI22D1BWP30P140LVT U135 ( .A1(n212), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n108) );
  IOA21D1BWP30P140LVT U136 ( .A1(n20), .A2(i_data_bus[232]), .B(n108), .ZN(
        n109) );
  AOI21D1BWP30P140LVT U137 ( .A1(n3), .A2(i_data_bus[8]), .B(n109), .ZN(n112)
         );
  AOI22D1BWP30P140LVT U138 ( .A1(n166), .A2(i_data_bus[72]), .B1(n2), .B2(
        i_data_bus[40]), .ZN(n111) );
  AOI22D1BWP30P140LVT U139 ( .A1(n168), .A2(i_data_bus[104]), .B1(n167), .B2(
        i_data_bus[136]), .ZN(n110) );
  ND3D1BWP30P140LVT U140 ( .A1(n112), .A2(n111), .A3(n110), .ZN(N377) );
  AOI22D1BWP30P140LVT U141 ( .A1(n212), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n113) );
  IOA21D1BWP30P140LVT U142 ( .A1(n20), .A2(i_data_bus[229]), .B(n113), .ZN(
        n114) );
  AOI21D1BWP30P140LVT U143 ( .A1(n3), .A2(i_data_bus[5]), .B(n114), .ZN(n117)
         );
  AOI22D1BWP30P140LVT U144 ( .A1(n166), .A2(i_data_bus[69]), .B1(n2), .B2(
        i_data_bus[37]), .ZN(n116) );
  AOI22D1BWP30P140LVT U145 ( .A1(n168), .A2(i_data_bus[101]), .B1(n167), .B2(
        i_data_bus[133]), .ZN(n115) );
  ND3D1BWP30P140LVT U146 ( .A1(n117), .A2(n116), .A3(n115), .ZN(N374) );
  AOI22D1BWP30P140LVT U147 ( .A1(n212), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n118) );
  IOA21D1BWP30P140LVT U148 ( .A1(n20), .A2(i_data_bus[230]), .B(n118), .ZN(
        n119) );
  AOI21D1BWP30P140LVT U149 ( .A1(n3), .A2(i_data_bus[6]), .B(n119), .ZN(n122)
         );
  AOI22D1BWP30P140LVT U150 ( .A1(n166), .A2(i_data_bus[70]), .B1(n2), .B2(
        i_data_bus[38]), .ZN(n121) );
  AOI22D1BWP30P140LVT U151 ( .A1(n168), .A2(i_data_bus[102]), .B1(n167), .B2(
        i_data_bus[134]), .ZN(n120) );
  ND3D1BWP30P140LVT U152 ( .A1(n122), .A2(n121), .A3(n120), .ZN(N375) );
  IOA21D1BWP30P140LVT U153 ( .A1(n20), .A2(i_data_bus[231]), .B(n124), .ZN(
        n125) );
  AOI21D1BWP30P140LVT U154 ( .A1(n3), .A2(i_data_bus[7]), .B(n125), .ZN(n128)
         );
  AOI22D1BWP30P140LVT U155 ( .A1(n166), .A2(i_data_bus[71]), .B1(n2), .B2(
        i_data_bus[39]), .ZN(n127) );
  AOI22D1BWP30P140LVT U156 ( .A1(n168), .A2(i_data_bus[103]), .B1(n167), .B2(
        i_data_bus[135]), .ZN(n126) );
  ND3D1BWP30P140LVT U157 ( .A1(n128), .A2(n127), .A3(n126), .ZN(N376) );
  AOI22D1BWP30P140LVT U158 ( .A1(n212), .A2(i_data_bus[206]), .B1(n1), .B2(
        i_data_bus[174]), .ZN(n129) );
  IOA21D1BWP30P140LVT U159 ( .A1(n20), .A2(i_data_bus[238]), .B(n129), .ZN(
        n130) );
  AOI21D1BWP30P140LVT U160 ( .A1(n3), .A2(i_data_bus[14]), .B(n130), .ZN(n134)
         );
  INVD2BWP30P140LVT U161 ( .I(n231), .ZN(n222) );
  AOI22D1BWP30P140LVT U162 ( .A1(n222), .A2(i_data_bus[78]), .B1(n2), .B2(
        i_data_bus[46]), .ZN(n133) );
  INVD2BWP30P140LVT U163 ( .I(n131), .ZN(n233) );
  AOI22D1BWP30P140LVT U164 ( .A1(n233), .A2(i_data_bus[110]), .B1(n232), .B2(
        i_data_bus[142]), .ZN(n132) );
  ND3D1BWP30P140LVT U165 ( .A1(n134), .A2(n133), .A3(n132), .ZN(N383) );
  INVD1BWP30P140LVT U166 ( .I(i_data_bus[173]), .ZN(n135) );
  MAOI22D1BWP30P140LVT U167 ( .A1(n212), .A2(i_data_bus[205]), .B1(n136), .B2(
        n135), .ZN(n137) );
  IOA21D1BWP30P140LVT U168 ( .A1(n20), .A2(i_data_bus[237]), .B(n137), .ZN(
        n138) );
  AOI21D1BWP30P140LVT U169 ( .A1(n3), .A2(i_data_bus[13]), .B(n138), .ZN(n141)
         );
  AOI22D1BWP30P140LVT U170 ( .A1(n222), .A2(i_data_bus[77]), .B1(n2), .B2(
        i_data_bus[45]), .ZN(n140) );
  AOI22D1BWP30P140LVT U171 ( .A1(n233), .A2(i_data_bus[109]), .B1(n232), .B2(
        i_data_bus[141]), .ZN(n139) );
  ND3D1BWP30P140LVT U172 ( .A1(n141), .A2(n140), .A3(n139), .ZN(N382) );
  INVD1BWP30P140LVT U173 ( .I(i_data_bus[194]), .ZN(n142) );
  MAOI22D1BWP30P140LVT U174 ( .A1(n1), .A2(i_data_bus[162]), .B1(n219), .B2(
        n142), .ZN(n143) );
  IOA21D1BWP30P140LVT U175 ( .A1(n20), .A2(i_data_bus[226]), .B(n143), .ZN(
        n144) );
  AOI21D1BWP30P140LVT U176 ( .A1(n3), .A2(i_data_bus[2]), .B(n144), .ZN(n147)
         );
  AOI22D1BWP30P140LVT U177 ( .A1(n166), .A2(i_data_bus[66]), .B1(n2), .B2(
        i_data_bus[34]), .ZN(n146) );
  AOI22D1BWP30P140LVT U178 ( .A1(n168), .A2(i_data_bus[98]), .B1(n167), .B2(
        i_data_bus[130]), .ZN(n145) );
  ND3D1BWP30P140LVT U179 ( .A1(n147), .A2(n146), .A3(n145), .ZN(N371) );
  INVD1BWP30P140LVT U180 ( .I(i_data_bus[195]), .ZN(n148) );
  MAOI22D1BWP30P140LVT U181 ( .A1(n1), .A2(i_data_bus[163]), .B1(n219), .B2(
        n148), .ZN(n149) );
  IOA21D1BWP30P140LVT U182 ( .A1(n20), .A2(i_data_bus[227]), .B(n149), .ZN(
        n150) );
  AOI21D1BWP30P140LVT U183 ( .A1(n3), .A2(i_data_bus[3]), .B(n150), .ZN(n153)
         );
  AOI22D1BWP30P140LVT U184 ( .A1(n166), .A2(i_data_bus[67]), .B1(n2), .B2(
        i_data_bus[35]), .ZN(n152) );
  AOI22D1BWP30P140LVT U185 ( .A1(n168), .A2(i_data_bus[99]), .B1(n167), .B2(
        i_data_bus[131]), .ZN(n151) );
  ND3D1BWP30P140LVT U186 ( .A1(n153), .A2(n152), .A3(n151), .ZN(N372) );
  INVD1BWP30P140LVT U187 ( .I(i_data_bus[193]), .ZN(n154) );
  MAOI22D1BWP30P140LVT U188 ( .A1(n1), .A2(i_data_bus[161]), .B1(n219), .B2(
        n154), .ZN(n155) );
  IOA21D1BWP30P140LVT U189 ( .A1(n20), .A2(i_data_bus[225]), .B(n155), .ZN(
        n156) );
  AOI21D1BWP30P140LVT U190 ( .A1(n3), .A2(i_data_bus[1]), .B(n156), .ZN(n159)
         );
  AOI22D1BWP30P140LVT U191 ( .A1(n166), .A2(i_data_bus[65]), .B1(n2), .B2(
        i_data_bus[33]), .ZN(n158) );
  AOI22D1BWP30P140LVT U192 ( .A1(n168), .A2(i_data_bus[97]), .B1(n167), .B2(
        i_data_bus[129]), .ZN(n157) );
  ND3D1BWP30P140LVT U193 ( .A1(n159), .A2(n158), .A3(n157), .ZN(N370) );
  INVD1BWP30P140LVT U194 ( .I(i_data_bus[224]), .ZN(n165) );
  INVD1BWP30P140LVT U195 ( .I(i_data_bus[192]), .ZN(n160) );
  MAOI22D1BWP30P140LVT U196 ( .A1(n1), .A2(i_data_bus[160]), .B1(n219), .B2(
        n160), .ZN(n164) );
  INR2D1BWP30P140LVT U197 ( .A1(i_data_bus[0]), .B1(n161), .ZN(n162) );
  INVD1BWP30P140LVT U198 ( .I(n162), .ZN(n163) );
  OA211D1BWP30P140LVT U199 ( .A1(n21), .A2(n165), .B(n164), .C(n163), .Z(n171)
         );
  AOI22D1BWP30P140LVT U200 ( .A1(n166), .A2(i_data_bus[64]), .B1(n2), .B2(
        i_data_bus[32]), .ZN(n170) );
  AOI22D1BWP30P140LVT U201 ( .A1(n168), .A2(i_data_bus[96]), .B1(n167), .B2(
        i_data_bus[128]), .ZN(n169) );
  ND3D1BWP30P140LVT U202 ( .A1(n171), .A2(n170), .A3(n169), .ZN(N369) );
  AOI22D1BWP30P140LVT U203 ( .A1(n212), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n172) );
  IOA21D1BWP30P140LVT U204 ( .A1(n20), .A2(i_data_bus[248]), .B(n172), .ZN(
        n173) );
  AOI21D1BWP30P140LVT U205 ( .A1(n3), .A2(i_data_bus[24]), .B(n173), .ZN(n176)
         );
  AOI22D1BWP30P140LVT U206 ( .A1(n222), .A2(i_data_bus[88]), .B1(n2), .B2(
        i_data_bus[56]), .ZN(n175) );
  AOI22D1BWP30P140LVT U207 ( .A1(n233), .A2(i_data_bus[120]), .B1(n232), .B2(
        i_data_bus[152]), .ZN(n174) );
  ND3D1BWP30P140LVT U208 ( .A1(n176), .A2(n175), .A3(n174), .ZN(N393) );
  AOI22D1BWP30P140LVT U209 ( .A1(n212), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n177) );
  IOA21D1BWP30P140LVT U210 ( .A1(n20), .A2(i_data_bus[249]), .B(n177), .ZN(
        n178) );
  AOI21D1BWP30P140LVT U211 ( .A1(n3), .A2(i_data_bus[25]), .B(n178), .ZN(n181)
         );
  AOI22D1BWP30P140LVT U212 ( .A1(n222), .A2(i_data_bus[89]), .B1(n2), .B2(
        i_data_bus[57]), .ZN(n180) );
  AOI22D1BWP30P140LVT U213 ( .A1(n233), .A2(i_data_bus[121]), .B1(n232), .B2(
        i_data_bus[153]), .ZN(n179) );
  ND3D1BWP30P140LVT U214 ( .A1(n181), .A2(n180), .A3(n179), .ZN(N394) );
  AOI22D1BWP30P140LVT U215 ( .A1(n212), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n182) );
  IOA21D1BWP30P140LVT U216 ( .A1(n20), .A2(i_data_bus[247]), .B(n182), .ZN(
        n183) );
  AOI21D1BWP30P140LVT U217 ( .A1(n3), .A2(i_data_bus[23]), .B(n183), .ZN(n186)
         );
  AOI22D1BWP30P140LVT U218 ( .A1(n222), .A2(i_data_bus[87]), .B1(n2), .B2(
        i_data_bus[55]), .ZN(n185) );
  AOI22D1BWP30P140LVT U219 ( .A1(n233), .A2(i_data_bus[119]), .B1(n232), .B2(
        i_data_bus[151]), .ZN(n184) );
  ND3D1BWP30P140LVT U220 ( .A1(n186), .A2(n185), .A3(n184), .ZN(N392) );
  AOI22D1BWP30P140LVT U221 ( .A1(n212), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n187) );
  IOA21D1BWP30P140LVT U222 ( .A1(n20), .A2(i_data_bus[246]), .B(n187), .ZN(
        n188) );
  AOI21D1BWP30P140LVT U223 ( .A1(n3), .A2(i_data_bus[22]), .B(n188), .ZN(n191)
         );
  AOI22D1BWP30P140LVT U224 ( .A1(n222), .A2(i_data_bus[86]), .B1(n2), .B2(
        i_data_bus[54]), .ZN(n190) );
  AOI22D1BWP30P140LVT U225 ( .A1(n233), .A2(i_data_bus[118]), .B1(n232), .B2(
        i_data_bus[150]), .ZN(n189) );
  ND3D1BWP30P140LVT U226 ( .A1(n191), .A2(n190), .A3(n189), .ZN(N391) );
  AOI22D1BWP30P140LVT U227 ( .A1(n212), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n192) );
  IOA21D1BWP30P140LVT U228 ( .A1(n20), .A2(i_data_bus[245]), .B(n192), .ZN(
        n193) );
  AOI21D1BWP30P140LVT U229 ( .A1(n3), .A2(i_data_bus[21]), .B(n193), .ZN(n196)
         );
  AOI22D1BWP30P140LVT U230 ( .A1(n222), .A2(i_data_bus[85]), .B1(n2), .B2(
        i_data_bus[53]), .ZN(n195) );
  AOI22D1BWP30P140LVT U231 ( .A1(n233), .A2(i_data_bus[117]), .B1(n232), .B2(
        i_data_bus[149]), .ZN(n194) );
  ND3D1BWP30P140LVT U232 ( .A1(n196), .A2(n195), .A3(n194), .ZN(N390) );
  AOI22D1BWP30P140LVT U233 ( .A1(n212), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n197) );
  IOA21D1BWP30P140LVT U234 ( .A1(n20), .A2(i_data_bus[244]), .B(n197), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U235 ( .A1(n3), .A2(i_data_bus[20]), .B(n198), .ZN(n201)
         );
  AOI22D1BWP30P140LVT U236 ( .A1(n222), .A2(i_data_bus[84]), .B1(n2), .B2(
        i_data_bus[52]), .ZN(n200) );
  AOI22D1BWP30P140LVT U237 ( .A1(n233), .A2(i_data_bus[116]), .B1(n232), .B2(
        i_data_bus[148]), .ZN(n199) );
  ND3D1BWP30P140LVT U238 ( .A1(n201), .A2(n200), .A3(n199), .ZN(N389) );
  AOI22D1BWP30P140LVT U239 ( .A1(n212), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n202) );
  IOA21D1BWP30P140LVT U240 ( .A1(n20), .A2(i_data_bus[243]), .B(n202), .ZN(
        n203) );
  AOI21D1BWP30P140LVT U241 ( .A1(n3), .A2(i_data_bus[19]), .B(n203), .ZN(n206)
         );
  AOI22D1BWP30P140LVT U242 ( .A1(n222), .A2(i_data_bus[83]), .B1(n2), .B2(
        i_data_bus[51]), .ZN(n205) );
  AOI22D1BWP30P140LVT U243 ( .A1(n233), .A2(i_data_bus[115]), .B1(n232), .B2(
        i_data_bus[147]), .ZN(n204) );
  ND3D1BWP30P140LVT U244 ( .A1(n206), .A2(n205), .A3(n204), .ZN(N388) );
  AOI22D1BWP30P140LVT U245 ( .A1(n212), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n207) );
  IOA21D1BWP30P140LVT U246 ( .A1(n20), .A2(i_data_bus[242]), .B(n207), .ZN(
        n208) );
  AOI21D1BWP30P140LVT U247 ( .A1(n3), .A2(i_data_bus[18]), .B(n208), .ZN(n211)
         );
  AOI22D1BWP30P140LVT U248 ( .A1(n222), .A2(i_data_bus[82]), .B1(n2), .B2(
        i_data_bus[50]), .ZN(n210) );
  AOI22D1BWP30P140LVT U249 ( .A1(n233), .A2(i_data_bus[114]), .B1(n232), .B2(
        i_data_bus[146]), .ZN(n209) );
  ND3D1BWP30P140LVT U250 ( .A1(n211), .A2(n210), .A3(n209), .ZN(N387) );
  AOI22D1BWP30P140LVT U251 ( .A1(n212), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n213) );
  IOA21D1BWP30P140LVT U252 ( .A1(n20), .A2(i_data_bus[241]), .B(n213), .ZN(
        n214) );
  AOI21D1BWP30P140LVT U253 ( .A1(n3), .A2(i_data_bus[17]), .B(n214), .ZN(n217)
         );
  AOI22D1BWP30P140LVT U254 ( .A1(n222), .A2(i_data_bus[81]), .B1(n2), .B2(
        i_data_bus[49]), .ZN(n216) );
  AOI22D1BWP30P140LVT U255 ( .A1(n233), .A2(i_data_bus[113]), .B1(n232), .B2(
        i_data_bus[145]), .ZN(n215) );
  ND3D1BWP30P140LVT U256 ( .A1(n217), .A2(n216), .A3(n215), .ZN(N386) );
  INVD1BWP30P140LVT U257 ( .I(i_data_bus[208]), .ZN(n218) );
  MAOI22D1BWP30P140LVT U258 ( .A1(n1), .A2(i_data_bus[176]), .B1(n219), .B2(
        n218), .ZN(n220) );
  IOA21D1BWP30P140LVT U259 ( .A1(n20), .A2(i_data_bus[240]), .B(n220), .ZN(
        n221) );
  AOI21D1BWP30P140LVT U260 ( .A1(n3), .A2(i_data_bus[16]), .B(n221), .ZN(n225)
         );
  AOI22D1BWP30P140LVT U261 ( .A1(n222), .A2(i_data_bus[80]), .B1(n2), .B2(
        i_data_bus[48]), .ZN(n224) );
  AOI22D1BWP30P140LVT U262 ( .A1(n233), .A2(i_data_bus[112]), .B1(n232), .B2(
        i_data_bus[144]), .ZN(n223) );
  ND3D1BWP30P140LVT U263 ( .A1(n225), .A2(n224), .A3(n223), .ZN(N385) );
  AOI22D1BWP30P140LVT U264 ( .A1(n212), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n226) );
  IOA21D1BWP30P140LVT U265 ( .A1(n20), .A2(i_data_bus[239]), .B(n226), .ZN(
        n227) );
  AOI21D1BWP30P140LVT U266 ( .A1(n3), .A2(i_data_bus[15]), .B(n227), .ZN(n236)
         );
  INVD1BWP30P140LVT U267 ( .I(i_data_bus[79]), .ZN(n230) );
  INVD1BWP30P140LVT U268 ( .I(i_data_bus[47]), .ZN(n228) );
  OA22D1BWP30P140LVT U269 ( .A1(n231), .A2(n230), .B1(n229), .B2(n228), .Z(
        n235) );
  AOI22D1BWP30P140LVT U270 ( .A1(n233), .A2(i_data_bus[111]), .B1(n232), .B2(
        i_data_bus[143]), .ZN(n234) );
  ND3D1BWP30P140LVT U271 ( .A1(n236), .A2(n235), .A3(n234), .ZN(N384) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_7 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  NR2D1BWP30P140LVT U3 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n26) );
  CKND2D2BWP30P140LVT U4 ( .A1(n7), .A2(n6), .ZN(n25) );
  INR2D1BWP30P140LVT U5 ( .A1(n13), .B1(i_cmd[0]), .ZN(n14) );
  INR2D1BWP30P140LVT U6 ( .A1(n5), .B1(i_cmd[6]), .ZN(n6) );
  INVD1BWP30P140LVT U7 ( .I(n28), .ZN(n52) );
  ND3D2BWP30P140LVT U8 ( .A1(n39), .A2(i_cmd[0]), .A3(n9), .ZN(n59) );
  INVD2BWP30P140LVT U9 ( .I(n59), .ZN(n1) );
  INVD1BWP30P140LVT U10 ( .I(i_cmd[2]), .ZN(n12) );
  INVD1BWP30P140LVT U11 ( .I(n225), .ZN(n64) );
  INVD4BWP30P140LVT U12 ( .I(n43), .ZN(n225) );
  CKAN2D4BWP30P140LVT U13 ( .A1(n35), .A2(n31), .Z(n2) );
  INR2D2BWP30P140LVT U14 ( .A1(n22), .B1(n21), .ZN(n47) );
  INVD3BWP30P140LVT U15 ( .I(n69), .ZN(n176) );
  INVD2BWP30P140LVT U16 ( .I(n47), .ZN(n69) );
  INVD2BWP30P140LVT U17 ( .I(i_cmd[3]), .ZN(n4) );
  INVD1BWP30P140LVT U18 ( .I(n32), .ZN(n33) );
  ND2OPTIBD1BWP30P140LVT U19 ( .A1(n12), .A2(n11), .ZN(n32) );
  ND2OPTIBD2BWP30P140LVT U20 ( .A1(n12), .A2(n4), .ZN(n30) );
  INR2D1BWP30P140LVT U21 ( .A1(n26), .B1(n25), .ZN(n35) );
  INR2D1BWP30P140LVT U22 ( .A1(i_en), .B1(rst), .ZN(n13) );
  INVD2BWP30P140LVT U23 ( .I(n175), .ZN(n223) );
  INR2D1BWP30P140LVT U24 ( .A1(n8), .B1(n25), .ZN(n39) );
  NR2D1BWP30P140LVT U25 ( .A1(n30), .A2(i_cmd[1]), .ZN(n8) );
  ND2D1BWP30P140LVT U26 ( .A1(n116), .A2(i_data_bus[207]), .ZN(n49) );
  ND2D1BWP30P140LVT U27 ( .A1(n222), .A2(i_data_bus[175]), .ZN(n48) );
  NR2D1BWP30P140LVT U28 ( .A1(n30), .A2(n29), .ZN(n31) );
  ND2OPTIBD1BWP30P140LVT U29 ( .A1(i_valid[1]), .A2(i_cmd[1]), .ZN(n29) );
  OR2D1BWP30P140LVT U30 ( .A1(n17), .A2(n21), .Z(n43) );
  AOI21D1BWP30P140LVT U31 ( .A1(n1), .A2(i_data_bus[6]), .B(n24), .ZN(n42) );
  AOI22D1BWP30P140LVT U32 ( .A1(n228), .A2(i_data_bus[125]), .B1(n3), .B2(
        i_data_bus[157]), .ZN(n179) );
  NR2D1BWP30P140LVT U33 ( .A1(n28), .A2(n2), .ZN(n45) );
  NR2D1BWP30P140LVT U34 ( .A1(n138), .A2(n3), .ZN(n44) );
  AOI21D1BWP30P140LVT U35 ( .A1(n1), .A2(i_data_bus[14]), .B(n118), .ZN(n121)
         );
  CKAN2D4BWP30P140LVT U36 ( .A1(n39), .A2(n38), .Z(n3) );
  INVD1BWP30P140LVT U37 ( .I(n36), .ZN(n53) );
  INVD2BWP30P140LVT U38 ( .I(n53), .ZN(n138) );
  INVD2BWP30P140LVT U39 ( .I(n53), .ZN(n228) );
  INVD1BWP30P140LVT U40 ( .I(i_cmd[1]), .ZN(n11) );
  NR2OPTPAD1BWP30P140LVT U41 ( .A1(i_cmd[5]), .A2(i_cmd[7]), .ZN(n7) );
  INR2D1BWP30P140LVT U42 ( .A1(i_en), .B1(rst), .ZN(n5) );
  INR2D1BWP30P140LVT U43 ( .A1(i_valid[0]), .B1(i_cmd[4]), .ZN(n9) );
  ND2D1BWP30P140LVT U44 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n10) );
  OR3D1BWP30P140LVT U45 ( .A1(n10), .A2(i_cmd[5]), .A3(i_cmd[6]), .Z(n17) );
  NR2OPTPAD1BWP30P140LVT U46 ( .A1(i_cmd[3]), .A2(i_cmd[4]), .ZN(n15) );
  ND2OPTIBD1BWP30P140LVT U47 ( .A1(n15), .A2(n14), .ZN(n16) );
  OR2D2BWP30P140LVT U48 ( .A1(n32), .A2(n16), .Z(n21) );
  ND2D1BWP30P140LVT U49 ( .A1(i_valid[6]), .A2(i_cmd[6]), .ZN(n18) );
  NR3D0P7BWP30P140LVT U50 ( .A1(n18), .A2(i_cmd[5]), .A3(i_cmd[7]), .ZN(n19)
         );
  INR2D2BWP30P140LVT U51 ( .A1(n19), .B1(n21), .ZN(n57) );
  BUFFD2BWP30P140LVT U52 ( .I(n57), .Z(n116) );
  INVD1BWP30P140LVT U53 ( .I(i_cmd[5]), .ZN(n20) );
  INR4D1BWP30P140LVT U54 ( .A1(i_valid[5]), .B1(i_cmd[6]), .B2(i_cmd[7]), .B3(
        n20), .ZN(n22) );
  AOI22D1BWP30P140LVT U55 ( .A1(n116), .A2(i_data_bus[198]), .B1(n176), .B2(
        i_data_bus[166]), .ZN(n23) );
  IOA21D1BWP30P140LVT U56 ( .A1(n225), .A2(i_data_bus[230]), .B(n23), .ZN(n24)
         );
  ND4D1BWP30P140LVT U57 ( .A1(n11), .A2(n4), .A3(i_cmd[2]), .A4(i_valid[2]), 
        .ZN(n27) );
  INR2D1BWP30P140LVT U58 ( .A1(n35), .B1(n27), .ZN(n28) );
  INVD2BWP30P140LVT U59 ( .I(n52), .ZN(n137) );
  AOI22D1BWP30P140LVT U60 ( .A1(n137), .A2(i_data_bus[70]), .B1(n2), .B2(
        i_data_bus[38]), .ZN(n41) );
  ND3D1BWP30P140LVT U61 ( .A1(n33), .A2(i_cmd[3]), .A3(i_valid[3]), .ZN(n34)
         );
  INR2D1BWP30P140LVT U62 ( .A1(n35), .B1(n34), .ZN(n36) );
  IND3D1BWP30P140LVT U63 ( .A1(i_cmd[0]), .B1(i_cmd[4]), .B2(i_valid[4]), .ZN(
        n37) );
  INVD1BWP30P140LVT U64 ( .I(n37), .ZN(n38) );
  AOI22D1BWP30P140LVT U65 ( .A1(n138), .A2(i_data_bus[102]), .B1(n3), .B2(
        i_data_bus[134]), .ZN(n40) );
  ND3D1BWP30P140LVT U66 ( .A1(n42), .A2(n41), .A3(n40), .ZN(N375) );
  NR4D0BWP30P140LVT U67 ( .A1(n1), .A2(n225), .A3(n116), .A4(n176), .ZN(n46)
         );
  ND3D1BWP30P140LVT U68 ( .A1(n46), .A2(n45), .A3(n44), .ZN(N402) );
  INVD1BWP30P140LVT U69 ( .I(i_data_bus[239]), .ZN(n50) );
  BUFFD4BWP30P140LVT U70 ( .I(n47), .Z(n222) );
  OAI211D1BWP30P140LVT U71 ( .A1(n64), .A2(n50), .B(n49), .C(n48), .ZN(n51) );
  AOI21D1BWP30P140LVT U72 ( .A1(n1), .A2(i_data_bus[15]), .B(n51), .ZN(n56) );
  INVD2BWP30P140LVT U73 ( .I(n52), .ZN(n227) );
  AOI22D1BWP30P140LVT U74 ( .A1(n227), .A2(i_data_bus[79]), .B1(n2), .B2(
        i_data_bus[47]), .ZN(n55) );
  AOI22D1BWP30P140LVT U75 ( .A1(n228), .A2(i_data_bus[111]), .B1(n3), .B2(
        i_data_bus[143]), .ZN(n54) );
  ND3D1BWP30P140LVT U76 ( .A1(n56), .A2(n55), .A3(n54), .ZN(N384) );
  INVD1BWP30P140LVT U77 ( .I(i_data_bus[224]), .ZN(n63) );
  INVD2BWP30P140LVT U78 ( .I(n57), .ZN(n175) );
  INVD1BWP30P140LVT U79 ( .I(i_data_bus[192]), .ZN(n58) );
  MAOI22D1BWP30P140LVT U80 ( .A1(n222), .A2(i_data_bus[160]), .B1(n175), .B2(
        n58), .ZN(n62) );
  INR2D1BWP30P140LVT U81 ( .A1(i_data_bus[0]), .B1(n59), .ZN(n60) );
  INVD1BWP30P140LVT U82 ( .I(n60), .ZN(n61) );
  OA211D1BWP30P140LVT U83 ( .A1(n64), .A2(n63), .B(n62), .C(n61), .Z(n67) );
  AOI22D1BWP30P140LVT U84 ( .A1(n137), .A2(i_data_bus[64]), .B1(n2), .B2(
        i_data_bus[32]), .ZN(n66) );
  AOI22D1BWP30P140LVT U85 ( .A1(n138), .A2(i_data_bus[96]), .B1(n3), .B2(
        i_data_bus[128]), .ZN(n65) );
  ND3D1BWP30P140LVT U86 ( .A1(n66), .A2(n67), .A3(n65), .ZN(N369) );
  INVD1BWP30P140LVT U87 ( .I(i_data_bus[173]), .ZN(n68) );
  MAOI22D1BWP30P140LVT U88 ( .A1(n116), .A2(i_data_bus[205]), .B1(n69), .B2(
        n68), .ZN(n70) );
  IOA21D1BWP30P140LVT U89 ( .A1(n225), .A2(i_data_bus[237]), .B(n70), .ZN(n71)
         );
  AOI21D1BWP30P140LVT U90 ( .A1(n1), .A2(i_data_bus[13]), .B(n71), .ZN(n74) );
  AOI22D1BWP30P140LVT U91 ( .A1(n227), .A2(i_data_bus[77]), .B1(n2), .B2(
        i_data_bus[45]), .ZN(n73) );
  AOI22D1BWP30P140LVT U92 ( .A1(n228), .A2(i_data_bus[109]), .B1(n3), .B2(
        i_data_bus[141]), .ZN(n72) );
  ND3D1BWP30P140LVT U93 ( .A1(n74), .A2(n73), .A3(n72), .ZN(N382) );
  INVD1BWP30P140LVT U94 ( .I(i_data_bus[8]), .ZN(n77) );
  AOI22D1BWP30P140LVT U95 ( .A1(n116), .A2(i_data_bus[200]), .B1(n176), .B2(
        i_data_bus[168]), .ZN(n75) );
  IOA21D1BWP30P140LVT U96 ( .A1(n225), .A2(i_data_bus[232]), .B(n75), .ZN(n76)
         );
  IAO21D1BWP30P140LVT U97 ( .A1(n59), .A2(n77), .B(n76), .ZN(n80) );
  AOI22D1BWP30P140LVT U98 ( .A1(n137), .A2(i_data_bus[72]), .B1(n2), .B2(
        i_data_bus[40]), .ZN(n79) );
  AOI22D1BWP30P140LVT U99 ( .A1(n138), .A2(i_data_bus[104]), .B1(n3), .B2(
        i_data_bus[136]), .ZN(n78) );
  ND3D1BWP30P140LVT U100 ( .A1(n80), .A2(n79), .A3(n78), .ZN(N377) );
  AOI22D1BWP30P140LVT U101 ( .A1(n116), .A2(i_data_bus[199]), .B1(n176), .B2(
        i_data_bus[167]), .ZN(n81) );
  IOA21D1BWP30P140LVT U102 ( .A1(n225), .A2(i_data_bus[231]), .B(n81), .ZN(n82) );
  AOI21D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[7]), .B(n82), .ZN(n85) );
  AOI22D1BWP30P140LVT U104 ( .A1(n137), .A2(i_data_bus[71]), .B1(n2), .B2(
        i_data_bus[39]), .ZN(n84) );
  AOI22D1BWP30P140LVT U105 ( .A1(n138), .A2(i_data_bus[103]), .B1(n3), .B2(
        i_data_bus[135]), .ZN(n83) );
  ND3D1BWP30P140LVT U106 ( .A1(n85), .A2(n84), .A3(n83), .ZN(N376) );
  AOI22D1BWP30P140LVT U107 ( .A1(n116), .A2(i_data_bus[204]), .B1(n176), .B2(
        i_data_bus[172]), .ZN(n86) );
  IOA21D1BWP30P140LVT U108 ( .A1(n225), .A2(i_data_bus[236]), .B(n86), .ZN(n87) );
  AOI21D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[12]), .B(n87), .ZN(n90)
         );
  AOI22D1BWP30P140LVT U110 ( .A1(n137), .A2(i_data_bus[76]), .B1(n2), .B2(
        i_data_bus[44]), .ZN(n89) );
  AOI22D1BWP30P140LVT U111 ( .A1(n138), .A2(i_data_bus[108]), .B1(n3), .B2(
        i_data_bus[140]), .ZN(n88) );
  ND3D1BWP30P140LVT U112 ( .A1(n90), .A2(n89), .A3(n88), .ZN(N381) );
  AOI22D1BWP30P140LVT U113 ( .A1(n116), .A2(i_data_bus[197]), .B1(n176), .B2(
        i_data_bus[165]), .ZN(n91) );
  IOA21D1BWP30P140LVT U114 ( .A1(n225), .A2(i_data_bus[229]), .B(n91), .ZN(n92) );
  AOI21D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[5]), .B(n92), .ZN(n95) );
  AOI22D1BWP30P140LVT U116 ( .A1(n137), .A2(i_data_bus[69]), .B1(n2), .B2(
        i_data_bus[37]), .ZN(n94) );
  AOI22D1BWP30P140LVT U117 ( .A1(n138), .A2(i_data_bus[101]), .B1(n3), .B2(
        i_data_bus[133]), .ZN(n93) );
  ND3D1BWP30P140LVT U118 ( .A1(n95), .A2(n94), .A3(n93), .ZN(N374) );
  AOI22D1BWP30P140LVT U119 ( .A1(n116), .A2(i_data_bus[203]), .B1(n176), .B2(
        i_data_bus[171]), .ZN(n96) );
  IOA21D1BWP30P140LVT U120 ( .A1(n225), .A2(i_data_bus[235]), .B(n96), .ZN(n97) );
  AOI21D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[11]), .B(n97), .ZN(n100)
         );
  AOI22D1BWP30P140LVT U122 ( .A1(n137), .A2(i_data_bus[75]), .B1(n2), .B2(
        i_data_bus[43]), .ZN(n99) );
  AOI22D1BWP30P140LVT U123 ( .A1(n138), .A2(i_data_bus[107]), .B1(n3), .B2(
        i_data_bus[139]), .ZN(n98) );
  ND3D1BWP30P140LVT U124 ( .A1(n100), .A2(n99), .A3(n98), .ZN(N380) );
  AOI22D1BWP30P140LVT U125 ( .A1(n116), .A2(i_data_bus[201]), .B1(n176), .B2(
        i_data_bus[169]), .ZN(n101) );
  IOA21D1BWP30P140LVT U126 ( .A1(n225), .A2(i_data_bus[233]), .B(n101), .ZN(
        n102) );
  AOI21D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[9]), .B(n102), .ZN(n105)
         );
  AOI22D1BWP30P140LVT U128 ( .A1(n137), .A2(i_data_bus[73]), .B1(n2), .B2(
        i_data_bus[41]), .ZN(n104) );
  AOI22D1BWP30P140LVT U129 ( .A1(n138), .A2(i_data_bus[105]), .B1(n3), .B2(
        i_data_bus[137]), .ZN(n103) );
  ND3D1BWP30P140LVT U130 ( .A1(n105), .A2(n104), .A3(n103), .ZN(N378) );
  AOI22D1BWP30P140LVT U131 ( .A1(n116), .A2(i_data_bus[196]), .B1(n176), .B2(
        i_data_bus[164]), .ZN(n106) );
  IOA21D1BWP30P140LVT U132 ( .A1(n225), .A2(i_data_bus[228]), .B(n106), .ZN(
        n107) );
  AOI21D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[4]), .B(n107), .ZN(n110)
         );
  AOI22D1BWP30P140LVT U134 ( .A1(n137), .A2(i_data_bus[68]), .B1(n2), .B2(
        i_data_bus[36]), .ZN(n109) );
  AOI22D1BWP30P140LVT U135 ( .A1(n138), .A2(i_data_bus[100]), .B1(n3), .B2(
        i_data_bus[132]), .ZN(n108) );
  ND3D1BWP30P140LVT U136 ( .A1(n110), .A2(n109), .A3(n108), .ZN(N373) );
  AOI22D1BWP30P140LVT U137 ( .A1(n116), .A2(i_data_bus[202]), .B1(n176), .B2(
        i_data_bus[170]), .ZN(n111) );
  IOA21D1BWP30P140LVT U138 ( .A1(n225), .A2(i_data_bus[234]), .B(n111), .ZN(
        n112) );
  AOI21D1BWP30P140LVT U139 ( .A1(n1), .A2(i_data_bus[10]), .B(n112), .ZN(n115)
         );
  AOI22D1BWP30P140LVT U140 ( .A1(n137), .A2(i_data_bus[74]), .B1(n2), .B2(
        i_data_bus[42]), .ZN(n114) );
  AOI22D1BWP30P140LVT U141 ( .A1(n138), .A2(i_data_bus[106]), .B1(n3), .B2(
        i_data_bus[138]), .ZN(n113) );
  ND3D1BWP30P140LVT U142 ( .A1(n115), .A2(n114), .A3(n113), .ZN(N379) );
  AOI22D1BWP30P140LVT U143 ( .A1(n116), .A2(i_data_bus[206]), .B1(n176), .B2(
        i_data_bus[174]), .ZN(n117) );
  IOA21D1BWP30P140LVT U144 ( .A1(n225), .A2(i_data_bus[238]), .B(n117), .ZN(
        n118) );
  AOI22D1BWP30P140LVT U145 ( .A1(n227), .A2(i_data_bus[78]), .B1(n2), .B2(
        i_data_bus[46]), .ZN(n120) );
  AOI22D1BWP30P140LVT U146 ( .A1(n228), .A2(i_data_bus[110]), .B1(n3), .B2(
        i_data_bus[142]), .ZN(n119) );
  ND3D1BWP30P140LVT U147 ( .A1(n121), .A2(n120), .A3(n119), .ZN(N383) );
  INVD1BWP30P140LVT U148 ( .I(i_data_bus[195]), .ZN(n122) );
  MAOI22D1BWP30P140LVT U149 ( .A1(n176), .A2(i_data_bus[163]), .B1(n175), .B2(
        n122), .ZN(n123) );
  IOA21D1BWP30P140LVT U150 ( .A1(n225), .A2(i_data_bus[227]), .B(n123), .ZN(
        n124) );
  AOI21D1BWP30P140LVT U151 ( .A1(n1), .A2(i_data_bus[3]), .B(n124), .ZN(n127)
         );
  AOI22D1BWP30P140LVT U152 ( .A1(n137), .A2(i_data_bus[67]), .B1(n2), .B2(
        i_data_bus[35]), .ZN(n126) );
  AOI22D1BWP30P140LVT U153 ( .A1(n138), .A2(i_data_bus[99]), .B1(n3), .B2(
        i_data_bus[131]), .ZN(n125) );
  ND3D1BWP30P140LVT U154 ( .A1(n127), .A2(n126), .A3(n125), .ZN(N372) );
  INVD1BWP30P140LVT U155 ( .I(i_data_bus[194]), .ZN(n128) );
  MAOI22D1BWP30P140LVT U156 ( .A1(n176), .A2(i_data_bus[162]), .B1(n175), .B2(
        n128), .ZN(n129) );
  IOA21D1BWP30P140LVT U157 ( .A1(n225), .A2(i_data_bus[226]), .B(n129), .ZN(
        n130) );
  AOI21D1BWP30P140LVT U158 ( .A1(n1), .A2(i_data_bus[2]), .B(n130), .ZN(n133)
         );
  AOI22D1BWP30P140LVT U159 ( .A1(n137), .A2(i_data_bus[66]), .B1(n2), .B2(
        i_data_bus[34]), .ZN(n132) );
  AOI22D1BWP30P140LVT U160 ( .A1(n138), .A2(i_data_bus[98]), .B1(n3), .B2(
        i_data_bus[130]), .ZN(n131) );
  ND3D1BWP30P140LVT U161 ( .A1(n133), .A2(n132), .A3(n131), .ZN(N371) );
  INVD1BWP30P140LVT U162 ( .I(i_data_bus[193]), .ZN(n134) );
  MAOI22D1BWP30P140LVT U163 ( .A1(n176), .A2(i_data_bus[161]), .B1(n175), .B2(
        n134), .ZN(n135) );
  IOA21D1BWP30P140LVT U164 ( .A1(n225), .A2(i_data_bus[225]), .B(n135), .ZN(
        n136) );
  AOI21D1BWP30P140LVT U165 ( .A1(n1), .A2(i_data_bus[1]), .B(n136), .ZN(n141)
         );
  AOI22D1BWP30P140LVT U166 ( .A1(n137), .A2(i_data_bus[65]), .B1(n2), .B2(
        i_data_bus[33]), .ZN(n140) );
  AOI22D1BWP30P140LVT U167 ( .A1(n138), .A2(i_data_bus[97]), .B1(n3), .B2(
        i_data_bus[129]), .ZN(n139) );
  ND3D1BWP30P140LVT U168 ( .A1(n141), .A2(n140), .A3(n139), .ZN(N370) );
  AOI22D1BWP30P140LVT U169 ( .A1(n223), .A2(i_data_bus[220]), .B1(n222), .B2(
        i_data_bus[188]), .ZN(n142) );
  IOA21D1BWP30P140LVT U170 ( .A1(n225), .A2(i_data_bus[252]), .B(n142), .ZN(
        n143) );
  AOI21D1BWP30P140LVT U171 ( .A1(n1), .A2(i_data_bus[28]), .B(n143), .ZN(n146)
         );
  AOI22D1BWP30P140LVT U172 ( .A1(n227), .A2(i_data_bus[92]), .B1(n2), .B2(
        i_data_bus[60]), .ZN(n145) );
  AOI22D1BWP30P140LVT U173 ( .A1(n138), .A2(i_data_bus[124]), .B1(n3), .B2(
        i_data_bus[156]), .ZN(n144) );
  ND3D1BWP30P140LVT U174 ( .A1(n146), .A2(n145), .A3(n144), .ZN(N397) );
  AOI22D1BWP30P140LVT U175 ( .A1(n223), .A2(i_data_bus[219]), .B1(n222), .B2(
        i_data_bus[187]), .ZN(n147) );
  IOA21D1BWP30P140LVT U176 ( .A1(n225), .A2(i_data_bus[251]), .B(n147), .ZN(
        n148) );
  AOI21D1BWP30P140LVT U177 ( .A1(n1), .A2(i_data_bus[27]), .B(n148), .ZN(n151)
         );
  AOI22D1BWP30P140LVT U178 ( .A1(n137), .A2(i_data_bus[91]), .B1(n2), .B2(
        i_data_bus[59]), .ZN(n150) );
  AOI22D1BWP30P140LVT U179 ( .A1(n228), .A2(i_data_bus[123]), .B1(n3), .B2(
        i_data_bus[155]), .ZN(n149) );
  ND3D1BWP30P140LVT U180 ( .A1(n151), .A2(n150), .A3(n149), .ZN(N396) );
  AOI22D1BWP30P140LVT U181 ( .A1(n223), .A2(i_data_bus[218]), .B1(n222), .B2(
        i_data_bus[186]), .ZN(n152) );
  IOA21D1BWP30P140LVT U182 ( .A1(n225), .A2(i_data_bus[250]), .B(n152), .ZN(
        n153) );
  AOI21D1BWP30P140LVT U183 ( .A1(n1), .A2(i_data_bus[26]), .B(n153), .ZN(n156)
         );
  AOI22D1BWP30P140LVT U184 ( .A1(n227), .A2(i_data_bus[90]), .B1(n2), .B2(
        i_data_bus[58]), .ZN(n155) );
  AOI22D1BWP30P140LVT U185 ( .A1(n138), .A2(i_data_bus[122]), .B1(n3), .B2(
        i_data_bus[154]), .ZN(n154) );
  ND3D1BWP30P140LVT U186 ( .A1(n156), .A2(n155), .A3(n154), .ZN(N395) );
  AOI22D1BWP30P140LVT U187 ( .A1(n223), .A2(i_data_bus[217]), .B1(n222), .B2(
        i_data_bus[185]), .ZN(n157) );
  IOA21D1BWP30P140LVT U188 ( .A1(n225), .A2(i_data_bus[249]), .B(n157), .ZN(
        n158) );
  AOI21D1BWP30P140LVT U189 ( .A1(n1), .A2(i_data_bus[25]), .B(n158), .ZN(n161)
         );
  AOI22D1BWP30P140LVT U190 ( .A1(n227), .A2(i_data_bus[89]), .B1(n2), .B2(
        i_data_bus[57]), .ZN(n160) );
  AOI22D1BWP30P140LVT U191 ( .A1(n228), .A2(i_data_bus[121]), .B1(n3), .B2(
        i_data_bus[153]), .ZN(n159) );
  ND3D1BWP30P140LVT U192 ( .A1(n161), .A2(n160), .A3(n159), .ZN(N394) );
  INVD1BWP30P140LVT U193 ( .I(i_data_bus[222]), .ZN(n162) );
  MAOI22D1BWP30P140LVT U194 ( .A1(n176), .A2(i_data_bus[190]), .B1(n175), .B2(
        n162), .ZN(n163) );
  IOA21D1BWP30P140LVT U195 ( .A1(n225), .A2(i_data_bus[254]), .B(n163), .ZN(
        n164) );
  AOI21D1BWP30P140LVT U196 ( .A1(n1), .A2(i_data_bus[30]), .B(n164), .ZN(n167)
         );
  AOI22D1BWP30P140LVT U197 ( .A1(n137), .A2(i_data_bus[94]), .B1(n2), .B2(
        i_data_bus[62]), .ZN(n166) );
  AOI22D1BWP30P140LVT U198 ( .A1(n228), .A2(i_data_bus[126]), .B1(n3), .B2(
        i_data_bus[158]), .ZN(n165) );
  ND3D1BWP30P140LVT U199 ( .A1(n167), .A2(n166), .A3(n165), .ZN(N399) );
  INVD1BWP30P140LVT U200 ( .I(i_data_bus[223]), .ZN(n168) );
  MAOI22D1BWP30P140LVT U201 ( .A1(n176), .A2(i_data_bus[191]), .B1(n175), .B2(
        n168), .ZN(n169) );
  IOA21D1BWP30P140LVT U202 ( .A1(n225), .A2(i_data_bus[255]), .B(n169), .ZN(
        n170) );
  AOI21D1BWP30P140LVT U203 ( .A1(n1), .A2(i_data_bus[31]), .B(n170), .ZN(n173)
         );
  AOI22D1BWP30P140LVT U204 ( .A1(n227), .A2(i_data_bus[95]), .B1(n2), .B2(
        i_data_bus[63]), .ZN(n172) );
  AOI22D1BWP30P140LVT U205 ( .A1(n138), .A2(i_data_bus[127]), .B1(n3), .B2(
        i_data_bus[159]), .ZN(n171) );
  ND3D1BWP30P140LVT U206 ( .A1(n173), .A2(n172), .A3(n171), .ZN(N400) );
  INVD1BWP30P140LVT U207 ( .I(i_data_bus[221]), .ZN(n174) );
  MAOI22D1BWP30P140LVT U208 ( .A1(n176), .A2(i_data_bus[189]), .B1(n175), .B2(
        n174), .ZN(n177) );
  IOA21D1BWP30P140LVT U209 ( .A1(n225), .A2(i_data_bus[253]), .B(n177), .ZN(
        n178) );
  AOI21D1BWP30P140LVT U210 ( .A1(n1), .A2(i_data_bus[29]), .B(n178), .ZN(n181)
         );
  AOI22D1BWP30P140LVT U211 ( .A1(n137), .A2(i_data_bus[93]), .B1(n2), .B2(
        i_data_bus[61]), .ZN(n180) );
  ND3D1BWP30P140LVT U212 ( .A1(n181), .A2(n180), .A3(n179), .ZN(N398) );
  AOI22D1BWP30P140LVT U213 ( .A1(n223), .A2(i_data_bus[211]), .B1(n222), .B2(
        i_data_bus[179]), .ZN(n182) );
  IOA21D1BWP30P140LVT U214 ( .A1(n225), .A2(i_data_bus[243]), .B(n182), .ZN(
        n183) );
  AOI21D1BWP30P140LVT U215 ( .A1(n1), .A2(i_data_bus[19]), .B(n183), .ZN(n186)
         );
  AOI22D1BWP30P140LVT U216 ( .A1(n227), .A2(i_data_bus[83]), .B1(n2), .B2(
        i_data_bus[51]), .ZN(n185) );
  AOI22D1BWP30P140LVT U217 ( .A1(n228), .A2(i_data_bus[115]), .B1(n3), .B2(
        i_data_bus[147]), .ZN(n184) );
  ND3D1BWP30P140LVT U218 ( .A1(n186), .A2(n185), .A3(n184), .ZN(N388) );
  AOI22D1BWP30P140LVT U219 ( .A1(n223), .A2(i_data_bus[212]), .B1(n222), .B2(
        i_data_bus[180]), .ZN(n187) );
  IOA21D1BWP30P140LVT U220 ( .A1(n225), .A2(i_data_bus[244]), .B(n187), .ZN(
        n188) );
  AOI21D1BWP30P140LVT U221 ( .A1(n1), .A2(i_data_bus[20]), .B(n188), .ZN(n191)
         );
  AOI22D1BWP30P140LVT U222 ( .A1(n227), .A2(i_data_bus[84]), .B1(n2), .B2(
        i_data_bus[52]), .ZN(n190) );
  AOI22D1BWP30P140LVT U223 ( .A1(n228), .A2(i_data_bus[116]), .B1(n3), .B2(
        i_data_bus[148]), .ZN(n189) );
  ND3D1BWP30P140LVT U224 ( .A1(n191), .A2(n190), .A3(n189), .ZN(N389) );
  AOI22D1BWP30P140LVT U225 ( .A1(n223), .A2(i_data_bus[208]), .B1(n222), .B2(
        i_data_bus[176]), .ZN(n192) );
  IOA21D1BWP30P140LVT U226 ( .A1(n225), .A2(i_data_bus[240]), .B(n192), .ZN(
        n193) );
  AOI21D1BWP30P140LVT U227 ( .A1(n1), .A2(i_data_bus[16]), .B(n193), .ZN(n196)
         );
  AOI22D1BWP30P140LVT U228 ( .A1(n227), .A2(i_data_bus[80]), .B1(n2), .B2(
        i_data_bus[48]), .ZN(n195) );
  AOI22D1BWP30P140LVT U229 ( .A1(n228), .A2(i_data_bus[112]), .B1(n3), .B2(
        i_data_bus[144]), .ZN(n194) );
  ND3D1BWP30P140LVT U230 ( .A1(n196), .A2(n195), .A3(n194), .ZN(N385) );
  AOI22D1BWP30P140LVT U231 ( .A1(n223), .A2(i_data_bus[216]), .B1(n222), .B2(
        i_data_bus[184]), .ZN(n197) );
  IOA21D1BWP30P140LVT U232 ( .A1(n225), .A2(i_data_bus[248]), .B(n197), .ZN(
        n198) );
  AOI21D1BWP30P140LVT U233 ( .A1(n1), .A2(i_data_bus[24]), .B(n198), .ZN(n201)
         );
  AOI22D1BWP30P140LVT U234 ( .A1(n227), .A2(i_data_bus[88]), .B1(n2), .B2(
        i_data_bus[56]), .ZN(n200) );
  AOI22D1BWP30P140LVT U235 ( .A1(n228), .A2(i_data_bus[120]), .B1(n3), .B2(
        i_data_bus[152]), .ZN(n199) );
  ND3D1BWP30P140LVT U236 ( .A1(n201), .A2(n200), .A3(n199), .ZN(N393) );
  AOI22D1BWP30P140LVT U237 ( .A1(n223), .A2(i_data_bus[215]), .B1(n222), .B2(
        i_data_bus[183]), .ZN(n202) );
  IOA21D1BWP30P140LVT U238 ( .A1(n225), .A2(i_data_bus[247]), .B(n202), .ZN(
        n203) );
  AOI21D1BWP30P140LVT U239 ( .A1(n1), .A2(i_data_bus[23]), .B(n203), .ZN(n206)
         );
  AOI22D1BWP30P140LVT U240 ( .A1(n227), .A2(i_data_bus[87]), .B1(n2), .B2(
        i_data_bus[55]), .ZN(n205) );
  AOI22D1BWP30P140LVT U241 ( .A1(n228), .A2(i_data_bus[119]), .B1(n3), .B2(
        i_data_bus[151]), .ZN(n204) );
  ND3D1BWP30P140LVT U242 ( .A1(n206), .A2(n205), .A3(n204), .ZN(N392) );
  AOI22D1BWP30P140LVT U243 ( .A1(n223), .A2(i_data_bus[214]), .B1(n222), .B2(
        i_data_bus[182]), .ZN(n207) );
  IOA21D1BWP30P140LVT U244 ( .A1(n225), .A2(i_data_bus[246]), .B(n207), .ZN(
        n208) );
  AOI21D1BWP30P140LVT U245 ( .A1(n1), .A2(i_data_bus[22]), .B(n208), .ZN(n211)
         );
  AOI22D1BWP30P140LVT U246 ( .A1(n227), .A2(i_data_bus[86]), .B1(n2), .B2(
        i_data_bus[54]), .ZN(n210) );
  AOI22D1BWP30P140LVT U247 ( .A1(n228), .A2(i_data_bus[118]), .B1(n3), .B2(
        i_data_bus[150]), .ZN(n209) );
  ND3D1BWP30P140LVT U248 ( .A1(n211), .A2(n210), .A3(n209), .ZN(N391) );
  AOI22D1BWP30P140LVT U249 ( .A1(n223), .A2(i_data_bus[210]), .B1(n222), .B2(
        i_data_bus[178]), .ZN(n212) );
  IOA21D1BWP30P140LVT U250 ( .A1(n225), .A2(i_data_bus[242]), .B(n212), .ZN(
        n213) );
  AOI21D1BWP30P140LVT U251 ( .A1(n1), .A2(i_data_bus[18]), .B(n213), .ZN(n216)
         );
  AOI22D1BWP30P140LVT U252 ( .A1(n227), .A2(i_data_bus[82]), .B1(n2), .B2(
        i_data_bus[50]), .ZN(n215) );
  AOI22D1BWP30P140LVT U253 ( .A1(n228), .A2(i_data_bus[114]), .B1(n3), .B2(
        i_data_bus[146]), .ZN(n214) );
  ND3D1BWP30P140LVT U254 ( .A1(n216), .A2(n215), .A3(n214), .ZN(N387) );
  AOI22D1BWP30P140LVT U255 ( .A1(n223), .A2(i_data_bus[209]), .B1(n222), .B2(
        i_data_bus[177]), .ZN(n217) );
  IOA21D1BWP30P140LVT U256 ( .A1(n225), .A2(i_data_bus[241]), .B(n217), .ZN(
        n218) );
  AOI21D1BWP30P140LVT U257 ( .A1(n1), .A2(i_data_bus[17]), .B(n218), .ZN(n221)
         );
  AOI22D1BWP30P140LVT U258 ( .A1(n227), .A2(i_data_bus[81]), .B1(n2), .B2(
        i_data_bus[49]), .ZN(n220) );
  AOI22D1BWP30P140LVT U259 ( .A1(n228), .A2(i_data_bus[113]), .B1(n3), .B2(
        i_data_bus[145]), .ZN(n219) );
  ND3D1BWP30P140LVT U260 ( .A1(n221), .A2(n220), .A3(n219), .ZN(N386) );
  AOI22D1BWP30P140LVT U261 ( .A1(n223), .A2(i_data_bus[213]), .B1(n222), .B2(
        i_data_bus[181]), .ZN(n224) );
  IOA21D1BWP30P140LVT U262 ( .A1(n225), .A2(i_data_bus[245]), .B(n224), .ZN(
        n226) );
  AOI21D1BWP30P140LVT U263 ( .A1(n1), .A2(i_data_bus[21]), .B(n226), .ZN(n231)
         );
  AOI22D1BWP30P140LVT U264 ( .A1(n227), .A2(i_data_bus[85]), .B1(n2), .B2(
        i_data_bus[53]), .ZN(n230) );
  AOI22D1BWP30P140LVT U265 ( .A1(n228), .A2(i_data_bus[117]), .B1(n3), .B2(
        i_data_bus[149]), .ZN(n229) );
  ND3D1BWP30P140LVT U266 ( .A1(n231), .A2(n230), .A3(n229), .ZN(N390) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        CLK, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input CLK, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;
  wire   [127:0] buf_in_last_level_0__i_data_o_buf;
  wire   [127:0] buf_in_last_level_1__i_data_o_buf;
  wire   [127:0] buf_in_last_level_2__i_data_o_buf;
  wire   [127:0] buf_in_last_level_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[0]), .Z(
        buf_in_last_level_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[0]), .Z(
        buf_in_last_level_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[0]), .Z(
        buf_in_last_level_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[0]), .Z(
        buf_in_last_level_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[1]), .Z(
        buf_in_last_level_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[1]), .Z(
        buf_in_last_level_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[1]), .Z(
        buf_in_last_level_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[1]), .Z(
        buf_in_last_level_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[2]), .Z(
        buf_in_last_level_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[2]), .Z(
        buf_in_last_level_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[2]), .Z(
        buf_in_last_level_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[2]), .Z(
        buf_in_last_level_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[3]), .Z(
        buf_in_last_level_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[3]), .Z(
        buf_in_last_level_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[3]), .Z(
        buf_in_last_level_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[3]), .Z(
        buf_in_last_level_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[4]), .Z(
        buf_in_last_level_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[4]), .Z(
        buf_in_last_level_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[4]), .Z(
        buf_in_last_level_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[4]), .Z(
        buf_in_last_level_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[5]), .Z(
        buf_in_last_level_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[5]), .Z(
        buf_in_last_level_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[5]), .Z(
        buf_in_last_level_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[5]), .Z(
        buf_in_last_level_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[6]), .Z(
        buf_in_last_level_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[6]), .Z(
        buf_in_last_level_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[6]), .Z(
        buf_in_last_level_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[6]), .Z(
        buf_in_last_level_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[7]), .Z(
        buf_in_last_level_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[7]), .Z(
        buf_in_last_level_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[7]), .Z(
        buf_in_last_level_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[7]), .Z(
        buf_in_last_level_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[8]), .Z(
        buf_in_last_level_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[8]), .Z(
        buf_in_last_level_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[8]), .Z(
        buf_in_last_level_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[8]), .Z(
        buf_in_last_level_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[9]), .Z(
        buf_in_last_level_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[9]), .Z(
        buf_in_last_level_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[9]), .Z(
        buf_in_last_level_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[9]), .Z(
        buf_in_last_level_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[10]), .Z(
        buf_in_last_level_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[10]), .Z(
        buf_in_last_level_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[10]), .Z(
        buf_in_last_level_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[10]), .Z(
        buf_in_last_level_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[11]), .Z(
        buf_in_last_level_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[11]), .Z(
        buf_in_last_level_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[11]), .Z(
        buf_in_last_level_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[11]), .Z(
        buf_in_last_level_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[12]), .Z(
        buf_in_last_level_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[12]), .Z(
        buf_in_last_level_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[12]), .Z(
        buf_in_last_level_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[12]), .Z(
        buf_in_last_level_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[13]), .Z(
        buf_in_last_level_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[13]), .Z(
        buf_in_last_level_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[13]), .Z(
        buf_in_last_level_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[13]), .Z(
        buf_in_last_level_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[14]), .Z(
        buf_in_last_level_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[14]), .Z(
        buf_in_last_level_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[14]), .Z(
        buf_in_last_level_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[14]), .Z(
        buf_in_last_level_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[15]), .Z(
        buf_in_last_level_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[15]), .Z(
        buf_in_last_level_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[15]), .Z(
        buf_in_last_level_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[15]), .Z(
        buf_in_last_level_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[16]), .Z(
        buf_in_last_level_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[16]), .Z(
        buf_in_last_level_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[16]), .Z(
        buf_in_last_level_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[16]), .Z(
        buf_in_last_level_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[17]), .Z(
        buf_in_last_level_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[17]), .Z(
        buf_in_last_level_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[17]), .Z(
        buf_in_last_level_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[17]), .Z(
        buf_in_last_level_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[18]), .Z(
        buf_in_last_level_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[18]), .Z(
        buf_in_last_level_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[18]), .Z(
        buf_in_last_level_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[18]), .Z(
        buf_in_last_level_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[19]), .Z(
        buf_in_last_level_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[19]), .Z(
        buf_in_last_level_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[19]), .Z(
        buf_in_last_level_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[19]), .Z(
        buf_in_last_level_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[20]), .Z(
        buf_in_last_level_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[20]), .Z(
        buf_in_last_level_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[20]), .Z(
        buf_in_last_level_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[20]), .Z(
        buf_in_last_level_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[21]), .Z(
        buf_in_last_level_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[21]), .Z(
        buf_in_last_level_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[21]), .Z(
        buf_in_last_level_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[21]), .Z(
        buf_in_last_level_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[22]), .Z(
        buf_in_last_level_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[22]), .Z(
        buf_in_last_level_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[22]), .Z(
        buf_in_last_level_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[22]), .Z(
        buf_in_last_level_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[23]), .Z(
        buf_in_last_level_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[23]), .Z(
        buf_in_last_level_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[23]), .Z(
        buf_in_last_level_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[23]), .Z(
        buf_in_last_level_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[24]), .Z(
        buf_in_last_level_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[24]), .Z(
        buf_in_last_level_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[24]), .Z(
        buf_in_last_level_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[24]), .Z(
        buf_in_last_level_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[25]), .Z(
        buf_in_last_level_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[25]), .Z(
        buf_in_last_level_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[25]), .Z(
        buf_in_last_level_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[25]), .Z(
        buf_in_last_level_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[26]), .Z(
        buf_in_last_level_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[26]), .Z(
        buf_in_last_level_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[26]), .Z(
        buf_in_last_level_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[26]), .Z(
        buf_in_last_level_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[27]), .Z(
        buf_in_last_level_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[27]), .Z(
        buf_in_last_level_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[27]), .Z(
        buf_in_last_level_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[27]), .Z(
        buf_in_last_level_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[28]), .Z(
        buf_in_last_level_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[28]), .Z(
        buf_in_last_level_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[28]), .Z(
        buf_in_last_level_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[28]), .Z(
        buf_in_last_level_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[29]), .Z(
        buf_in_last_level_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[29]), .Z(
        buf_in_last_level_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[29]), .Z(
        buf_in_last_level_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[29]), .Z(
        buf_in_last_level_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[30]), .Z(
        buf_in_last_level_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[30]), .Z(
        buf_in_last_level_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[30]), .Z(
        buf_in_last_level_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[30]), .Z(
        buf_in_last_level_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[31]), .Z(
        buf_in_last_level_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[31]), .Z(
        buf_in_last_level_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[31]), .Z(
        buf_in_last_level_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[31]), .Z(
        buf_in_last_level_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[32]), .Z(
        buf_in_last_level_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[32]), .Z(
        buf_in_last_level_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[32]), .Z(
        buf_in_last_level_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[32]), .Z(
        buf_in_last_level_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[33]), .Z(
        buf_in_last_level_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[33]), .Z(
        buf_in_last_level_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[33]), .Z(
        buf_in_last_level_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[33]), .Z(
        buf_in_last_level_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[34]), .Z(
        buf_in_last_level_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[34]), .Z(
        buf_in_last_level_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[34]), .Z(
        buf_in_last_level_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[34]), .Z(
        buf_in_last_level_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[35]), .Z(
        buf_in_last_level_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[35]), .Z(
        buf_in_last_level_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[35]), .Z(
        buf_in_last_level_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[35]), .Z(
        buf_in_last_level_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[36]), .Z(
        buf_in_last_level_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[36]), .Z(
        buf_in_last_level_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[36]), .Z(
        buf_in_last_level_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[36]), .Z(
        buf_in_last_level_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[37]), .Z(
        buf_in_last_level_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[37]), .Z(
        buf_in_last_level_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[37]), .Z(
        buf_in_last_level_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[37]), .Z(
        buf_in_last_level_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[38]), .Z(
        buf_in_last_level_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[38]), .Z(
        buf_in_last_level_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[38]), .Z(
        buf_in_last_level_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[38]), .Z(
        buf_in_last_level_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[39]), .Z(
        buf_in_last_level_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[39]), .Z(
        buf_in_last_level_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[39]), .Z(
        buf_in_last_level_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[39]), .Z(
        buf_in_last_level_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[40]), .Z(
        buf_in_last_level_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[40]), .Z(
        buf_in_last_level_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[40]), .Z(
        buf_in_last_level_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[40]), .Z(
        buf_in_last_level_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[41]), .Z(
        buf_in_last_level_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[41]), .Z(
        buf_in_last_level_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[41]), .Z(
        buf_in_last_level_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[41]), .Z(
        buf_in_last_level_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[42]), .Z(
        buf_in_last_level_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[42]), .Z(
        buf_in_last_level_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[42]), .Z(
        buf_in_last_level_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[42]), .Z(
        buf_in_last_level_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[43]), .Z(
        buf_in_last_level_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[43]), .Z(
        buf_in_last_level_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[43]), .Z(
        buf_in_last_level_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[43]), .Z(
        buf_in_last_level_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[44]), .Z(
        buf_in_last_level_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[44]), .Z(
        buf_in_last_level_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[44]), .Z(
        buf_in_last_level_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[44]), .Z(
        buf_in_last_level_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[45]), .Z(
        buf_in_last_level_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[45]), .Z(
        buf_in_last_level_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[45]), .Z(
        buf_in_last_level_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[45]), .Z(
        buf_in_last_level_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[46]), .Z(
        buf_in_last_level_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[46]), .Z(
        buf_in_last_level_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[46]), .Z(
        buf_in_last_level_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[46]), .Z(
        buf_in_last_level_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[47]), .Z(
        buf_in_last_level_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[47]), .Z(
        buf_in_last_level_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[47]), .Z(
        buf_in_last_level_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[47]), .Z(
        buf_in_last_level_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[48]), .Z(
        buf_in_last_level_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[48]), .Z(
        buf_in_last_level_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[48]), .Z(
        buf_in_last_level_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[48]), .Z(
        buf_in_last_level_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[49]), .Z(
        buf_in_last_level_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[49]), .Z(
        buf_in_last_level_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[49]), .Z(
        buf_in_last_level_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[49]), .Z(
        buf_in_last_level_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[50]), .Z(
        buf_in_last_level_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[50]), .Z(
        buf_in_last_level_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[50]), .Z(
        buf_in_last_level_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[50]), .Z(
        buf_in_last_level_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[51]), .Z(
        buf_in_last_level_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[51]), .Z(
        buf_in_last_level_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[51]), .Z(
        buf_in_last_level_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[51]), .Z(
        buf_in_last_level_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[52]), .Z(
        buf_in_last_level_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[52]), .Z(
        buf_in_last_level_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[52]), .Z(
        buf_in_last_level_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[52]), .Z(
        buf_in_last_level_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[53]), .Z(
        buf_in_last_level_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[53]), .Z(
        buf_in_last_level_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[53]), .Z(
        buf_in_last_level_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[53]), .Z(
        buf_in_last_level_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[54]), .Z(
        buf_in_last_level_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[54]), .Z(
        buf_in_last_level_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[54]), .Z(
        buf_in_last_level_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[54]), .Z(
        buf_in_last_level_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[55]), .Z(
        buf_in_last_level_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[55]), .Z(
        buf_in_last_level_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[55]), .Z(
        buf_in_last_level_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[55]), .Z(
        buf_in_last_level_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[56]), .Z(
        buf_in_last_level_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[56]), .Z(
        buf_in_last_level_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[56]), .Z(
        buf_in_last_level_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[56]), .Z(
        buf_in_last_level_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[57]), .Z(
        buf_in_last_level_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[57]), .Z(
        buf_in_last_level_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[57]), .Z(
        buf_in_last_level_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[57]), .Z(
        buf_in_last_level_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[58]), .Z(
        buf_in_last_level_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[58]), .Z(
        buf_in_last_level_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[58]), .Z(
        buf_in_last_level_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[58]), .Z(
        buf_in_last_level_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[59]), .Z(
        buf_in_last_level_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[59]), .Z(
        buf_in_last_level_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[59]), .Z(
        buf_in_last_level_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[59]), .Z(
        buf_in_last_level_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[60]), .Z(
        buf_in_last_level_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[60]), .Z(
        buf_in_last_level_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[60]), .Z(
        buf_in_last_level_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[60]), .Z(
        buf_in_last_level_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[61]), .Z(
        buf_in_last_level_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[61]), .Z(
        buf_in_last_level_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[61]), .Z(
        buf_in_last_level_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[61]), .Z(
        buf_in_last_level_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[62]), .Z(
        buf_in_last_level_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[62]), .Z(
        buf_in_last_level_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[62]), .Z(
        buf_in_last_level_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[62]), .Z(
        buf_in_last_level_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[63]), .Z(
        buf_in_last_level_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[63]), .Z(
        buf_in_last_level_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[63]), .Z(
        buf_in_last_level_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[63]), .Z(
        buf_in_last_level_3__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[64]), .Z(
        buf_in_last_level_0__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[64]), .Z(
        buf_in_last_level_1__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[64]), .Z(
        buf_in_last_level_2__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[64]), .Z(
        buf_in_last_level_3__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[65]), .Z(
        buf_in_last_level_0__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[65]), .Z(
        buf_in_last_level_1__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[65]), .Z(
        buf_in_last_level_2__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[65]), .Z(
        buf_in_last_level_3__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[66]), .Z(
        buf_in_last_level_0__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[66]), .Z(
        buf_in_last_level_1__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[66]), .Z(
        buf_in_last_level_2__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[66]), .Z(
        buf_in_last_level_3__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[67]), .Z(
        buf_in_last_level_0__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[67]), .Z(
        buf_in_last_level_1__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[67]), .Z(
        buf_in_last_level_2__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[67]), .Z(
        buf_in_last_level_3__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[68]), .Z(
        buf_in_last_level_0__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[68]), .Z(
        buf_in_last_level_1__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[68]), .Z(
        buf_in_last_level_2__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[68]), .Z(
        buf_in_last_level_3__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[69]), .Z(
        buf_in_last_level_0__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[69]), .Z(
        buf_in_last_level_1__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[69]), .Z(
        buf_in_last_level_2__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[69]), .Z(
        buf_in_last_level_3__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[70]), .Z(
        buf_in_last_level_0__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[70]), .Z(
        buf_in_last_level_1__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[70]), .Z(
        buf_in_last_level_2__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[70]), .Z(
        buf_in_last_level_3__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[71]), .Z(
        buf_in_last_level_0__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[71]), .Z(
        buf_in_last_level_1__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[71]), .Z(
        buf_in_last_level_2__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[71]), .Z(
        buf_in_last_level_3__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[72]), .Z(
        buf_in_last_level_0__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[72]), .Z(
        buf_in_last_level_1__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[72]), .Z(
        buf_in_last_level_2__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[72]), .Z(
        buf_in_last_level_3__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[73]), .Z(
        buf_in_last_level_0__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[73]), .Z(
        buf_in_last_level_1__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[73]), .Z(
        buf_in_last_level_2__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[73]), .Z(
        buf_in_last_level_3__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[74]), .Z(
        buf_in_last_level_0__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[74]), .Z(
        buf_in_last_level_1__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[74]), .Z(
        buf_in_last_level_2__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[74]), .Z(
        buf_in_last_level_3__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[75]), .Z(
        buf_in_last_level_0__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[75]), .Z(
        buf_in_last_level_1__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[75]), .Z(
        buf_in_last_level_2__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[75]), .Z(
        buf_in_last_level_3__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[76]), .Z(
        buf_in_last_level_0__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[76]), .Z(
        buf_in_last_level_1__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[76]), .Z(
        buf_in_last_level_2__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[76]), .Z(
        buf_in_last_level_3__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[77]), .Z(
        buf_in_last_level_0__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[77]), .Z(
        buf_in_last_level_1__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[77]), .Z(
        buf_in_last_level_2__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[77]), .Z(
        buf_in_last_level_3__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[78]), .Z(
        buf_in_last_level_0__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[78]), .Z(
        buf_in_last_level_1__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[78]), .Z(
        buf_in_last_level_2__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[78]), .Z(
        buf_in_last_level_3__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[79]), .Z(
        buf_in_last_level_0__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[79]), .Z(
        buf_in_last_level_1__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[79]), .Z(
        buf_in_last_level_2__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[79]), .Z(
        buf_in_last_level_3__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[80]), .Z(
        buf_in_last_level_0__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[80]), .Z(
        buf_in_last_level_1__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[80]), .Z(
        buf_in_last_level_2__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[80]), .Z(
        buf_in_last_level_3__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[81]), .Z(
        buf_in_last_level_0__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[81]), .Z(
        buf_in_last_level_1__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[81]), .Z(
        buf_in_last_level_2__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[81]), .Z(
        buf_in_last_level_3__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[82]), .Z(
        buf_in_last_level_0__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[82]), .Z(
        buf_in_last_level_1__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[82]), .Z(
        buf_in_last_level_2__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[82]), .Z(
        buf_in_last_level_3__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[83]), .Z(
        buf_in_last_level_0__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[83]), .Z(
        buf_in_last_level_1__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[83]), .Z(
        buf_in_last_level_2__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[83]), .Z(
        buf_in_last_level_3__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[84]), .Z(
        buf_in_last_level_0__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[84]), .Z(
        buf_in_last_level_1__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[84]), .Z(
        buf_in_last_level_2__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[84]), .Z(
        buf_in_last_level_3__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[85]), .Z(
        buf_in_last_level_0__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[85]), .Z(
        buf_in_last_level_1__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[85]), .Z(
        buf_in_last_level_2__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[85]), .Z(
        buf_in_last_level_3__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[86]), .Z(
        buf_in_last_level_0__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[86]), .Z(
        buf_in_last_level_1__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[86]), .Z(
        buf_in_last_level_2__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[86]), .Z(
        buf_in_last_level_3__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[87]), .Z(
        buf_in_last_level_0__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[87]), .Z(
        buf_in_last_level_1__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[87]), .Z(
        buf_in_last_level_2__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[87]), .Z(
        buf_in_last_level_3__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[88]), .Z(
        buf_in_last_level_0__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[88]), .Z(
        buf_in_last_level_1__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[88]), .Z(
        buf_in_last_level_2__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[88]), .Z(
        buf_in_last_level_3__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[89]), .Z(
        buf_in_last_level_0__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[89]), .Z(
        buf_in_last_level_1__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[89]), .Z(
        buf_in_last_level_2__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[89]), .Z(
        buf_in_last_level_3__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[90]), .Z(
        buf_in_last_level_0__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[90]), .Z(
        buf_in_last_level_1__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[90]), .Z(
        buf_in_last_level_2__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[90]), .Z(
        buf_in_last_level_3__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[91]), .Z(
        buf_in_last_level_0__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[91]), .Z(
        buf_in_last_level_1__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[91]), .Z(
        buf_in_last_level_2__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[91]), .Z(
        buf_in_last_level_3__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[92]), .Z(
        buf_in_last_level_0__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[92]), .Z(
        buf_in_last_level_1__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[92]), .Z(
        buf_in_last_level_2__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[92]), .Z(
        buf_in_last_level_3__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[93]), .Z(
        buf_in_last_level_0__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[93]), .Z(
        buf_in_last_level_1__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[93]), .Z(
        buf_in_last_level_2__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[93]), .Z(
        buf_in_last_level_3__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[94]), .Z(
        buf_in_last_level_0__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[94]), .Z(
        buf_in_last_level_1__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[94]), .Z(
        buf_in_last_level_2__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[94]), .Z(
        buf_in_last_level_3__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[95]), .Z(
        buf_in_last_level_0__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[95]), .Z(
        buf_in_last_level_1__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[95]), .Z(
        buf_in_last_level_2__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[95]), .Z(
        buf_in_last_level_3__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[96]), .Z(
        buf_in_last_level_0__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[96]), .Z(
        buf_in_last_level_1__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[96]), .Z(
        buf_in_last_level_2__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[96]), .Z(
        buf_in_last_level_3__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[97]), .Z(
        buf_in_last_level_0__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[97]), .Z(
        buf_in_last_level_1__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[97]), .Z(
        buf_in_last_level_2__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[97]), .Z(
        buf_in_last_level_3__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[98]), .Z(
        buf_in_last_level_0__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[98]), .Z(
        buf_in_last_level_1__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[98]), .Z(
        buf_in_last_level_2__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[98]), .Z(
        buf_in_last_level_3__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[99]), .Z(
        buf_in_last_level_0__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[99]), .Z(
        buf_in_last_level_1__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[99]), .Z(
        buf_in_last_level_2__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[99]), .Z(
        buf_in_last_level_3__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[100]), .Z(
        buf_in_last_level_0__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[100]), .Z(
        buf_in_last_level_1__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[100]), .Z(
        buf_in_last_level_2__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[100]), .Z(
        buf_in_last_level_3__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[101]), .Z(
        buf_in_last_level_0__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[101]), .Z(
        buf_in_last_level_1__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[101]), .Z(
        buf_in_last_level_2__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[101]), .Z(
        buf_in_last_level_3__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[102]), .Z(
        buf_in_last_level_0__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[102]), .Z(
        buf_in_last_level_1__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[102]), .Z(
        buf_in_last_level_2__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[102]), .Z(
        buf_in_last_level_3__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[103]), .Z(
        buf_in_last_level_0__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[103]), .Z(
        buf_in_last_level_1__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[103]), .Z(
        buf_in_last_level_2__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[103]), .Z(
        buf_in_last_level_3__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[104]), .Z(
        buf_in_last_level_0__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[104]), .Z(
        buf_in_last_level_1__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[104]), .Z(
        buf_in_last_level_2__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[104]), .Z(
        buf_in_last_level_3__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[105]), .Z(
        buf_in_last_level_0__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[105]), .Z(
        buf_in_last_level_1__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[105]), .Z(
        buf_in_last_level_2__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[105]), .Z(
        buf_in_last_level_3__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[106]), .Z(
        buf_in_last_level_0__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[106]), .Z(
        buf_in_last_level_1__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[106]), .Z(
        buf_in_last_level_2__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[106]), .Z(
        buf_in_last_level_3__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[107]), .Z(
        buf_in_last_level_0__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[107]), .Z(
        buf_in_last_level_1__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[107]), .Z(
        buf_in_last_level_2__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[107]), .Z(
        buf_in_last_level_3__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[108]), .Z(
        buf_in_last_level_0__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[108]), .Z(
        buf_in_last_level_1__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[108]), .Z(
        buf_in_last_level_2__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[108]), .Z(
        buf_in_last_level_3__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[109]), .Z(
        buf_in_last_level_0__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[109]), .Z(
        buf_in_last_level_1__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[109]), .Z(
        buf_in_last_level_2__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[109]), .Z(
        buf_in_last_level_3__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[110]), .Z(
        buf_in_last_level_0__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[110]), .Z(
        buf_in_last_level_1__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[110]), .Z(
        buf_in_last_level_2__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[110]), .Z(
        buf_in_last_level_3__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[111]), .Z(
        buf_in_last_level_0__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[111]), .Z(
        buf_in_last_level_1__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[111]), .Z(
        buf_in_last_level_2__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[111]), .Z(
        buf_in_last_level_3__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[112]), .Z(
        buf_in_last_level_0__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[112]), .Z(
        buf_in_last_level_1__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[112]), .Z(
        buf_in_last_level_2__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[112]), .Z(
        buf_in_last_level_3__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[113]), .Z(
        buf_in_last_level_0__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[113]), .Z(
        buf_in_last_level_1__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[113]), .Z(
        buf_in_last_level_2__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[113]), .Z(
        buf_in_last_level_3__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[114]), .Z(
        buf_in_last_level_0__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[114]), .Z(
        buf_in_last_level_1__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[114]), .Z(
        buf_in_last_level_2__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[114]), .Z(
        buf_in_last_level_3__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[115]), .Z(
        buf_in_last_level_0__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[115]), .Z(
        buf_in_last_level_1__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[115]), .Z(
        buf_in_last_level_2__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[115]), .Z(
        buf_in_last_level_3__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[116]), .Z(
        buf_in_last_level_0__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[116]), .Z(
        buf_in_last_level_1__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[116]), .Z(
        buf_in_last_level_2__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[116]), .Z(
        buf_in_last_level_3__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[117]), .Z(
        buf_in_last_level_0__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[117]), .Z(
        buf_in_last_level_1__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[117]), .Z(
        buf_in_last_level_2__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[117]), .Z(
        buf_in_last_level_3__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[118]), .Z(
        buf_in_last_level_0__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[118]), .Z(
        buf_in_last_level_1__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[118]), .Z(
        buf_in_last_level_2__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[118]), .Z(
        buf_in_last_level_3__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[119]), .Z(
        buf_in_last_level_0__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[119]), .Z(
        buf_in_last_level_1__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[119]), .Z(
        buf_in_last_level_2__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[119]), .Z(
        buf_in_last_level_3__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[120]), .Z(
        buf_in_last_level_0__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[120]), .Z(
        buf_in_last_level_1__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[120]), .Z(
        buf_in_last_level_2__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[120]), .Z(
        buf_in_last_level_3__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[121]), .Z(
        buf_in_last_level_0__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[121]), .Z(
        buf_in_last_level_1__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[121]), .Z(
        buf_in_last_level_2__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[121]), .Z(
        buf_in_last_level_3__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[122]), .Z(
        buf_in_last_level_0__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[122]), .Z(
        buf_in_last_level_1__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[122]), .Z(
        buf_in_last_level_2__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[122]), .Z(
        buf_in_last_level_3__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[123]), .Z(
        buf_in_last_level_0__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[123]), .Z(
        buf_in_last_level_1__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[123]), .Z(
        buf_in_last_level_2__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[123]), .Z(
        buf_in_last_level_3__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[124]), .Z(
        buf_in_last_level_0__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[124]), .Z(
        buf_in_last_level_1__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[124]), .Z(
        buf_in_last_level_2__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[124]), .Z(
        buf_in_last_level_3__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[125]), .Z(
        buf_in_last_level_0__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[125]), .Z(
        buf_in_last_level_1__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[125]), .Z(
        buf_in_last_level_2__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[125]), .Z(
        buf_in_last_level_3__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[126]), .Z(
        buf_in_last_level_0__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[126]), .Z(
        buf_in_last_level_1__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[126]), .Z(
        buf_in_last_level_2__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[126]), .Z(
        buf_in_last_level_3__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[127]), .Z(
        buf_in_last_level_0__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[127]), .Z(
        buf_in_last_level_1__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[127]), .Z(
        buf_in_last_level_2__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[127]), .Z(
        buf_in_last_level_3__i_data_o_buf[127]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(CLK), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(CLK), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(CLK), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(CLK), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(CLK), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(CLK), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(CLK), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(CLK), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[101]), .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[102]), .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[105]), .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[107]), .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[109]), .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[110]), .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[111]), .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[112]), .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[115]), .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[82]), .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[86]), .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[61]), .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[63]), .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[31]), .Z(N297) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[30]), .Z(N296) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[28]), .Z(N294) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[27]), .Z(N293) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[26]), .Z(N292) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[25]), .Z(N291) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[24]), .Z(N290) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[23]), .Z(N289) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[22]), .Z(N288) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[21]), .Z(N287) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[20]), .Z(N286) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[29]), .Z(N295) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[19]), .Z(N285) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[18]), .Z(N284) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[17]), .Z(N283) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[16]), .Z(N282) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[15]), .Z(N281) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[14]), .Z(N280) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[13]), .Z(N279) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[12]), .Z(N278) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[11]), .Z(N277) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[10]), .Z(N276) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[9]), .Z(N275) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[8]), .Z(N274) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[7]), .Z(N273) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[5]), .Z(N271) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[4]), .Z(N270) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[3]), .Z(N269) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[1]), .Z(N267) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[0]), .Z(N266) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[62]), .Z(N362) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[60]), .Z(N360) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[59]), .Z(N359) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[58]), .Z(N358) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[57]), .Z(N357) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[56]), .Z(N356) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[55]), .Z(N355) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[54]), .Z(N354) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[53]), .Z(N353) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[52]), .Z(N352) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[51]), .Z(N351) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[50]), .Z(N350) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[49]), .Z(N349) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[48]), .Z(N348) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[47]), .Z(N347) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[46]), .Z(N346) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[45]), .Z(N345) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[44]), .Z(N344) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[43]), .Z(N343) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[42]), .Z(N342) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[41]), .Z(N341) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[40]), .Z(N340) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[39]), .Z(N339) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[38]), .Z(N338) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[37]), .Z(N337) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[36]), .Z(N336) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[35]), .Z(N335) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[34]), .Z(N334) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[33]), .Z(N333) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[32]), .Z(N332) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[71]), .Z(N405) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[72]), .Z(N406) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[70]), .Z(N404) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[80]), .Z(N414) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[81]), .Z(N415) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[69]), .Z(N403) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[68]), .Z(N402) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[67]), .Z(N401) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[66]), .Z(N400) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[65]), .Z(N399) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[64]), .Z(N398) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[95]), .Z(N429) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[94]), .Z(N428) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[93]), .Z(N427) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[83]), .Z(N417) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[84]), .Z(N418) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[85]), .Z(N419) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[87]), .Z(N421) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[88]), .Z(N422) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[89]), .Z(N423) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[90]), .Z(N424) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[92]), .Z(N426) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[91]), .Z(N425) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[79]), .Z(N413) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[78]), .Z(N412) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[77]), .Z(N411) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[76]), .Z(N410) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[75]), .Z(N409) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[74]), .Z(N408) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[73]), .Z(N407) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        CLK, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input CLK, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;
  wire   [127:0] buf_in_last_level_0__i_data_o_buf;
  wire   [127:0] buf_in_last_level_1__i_data_o_buf;
  wire   [127:0] buf_in_last_level_2__i_data_o_buf;
  wire   [127:0] buf_in_last_level_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[0]), .Z(
        buf_in_last_level_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[0]), .Z(
        buf_in_last_level_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[0]), .Z(
        buf_in_last_level_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[0]), .Z(
        buf_in_last_level_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[1]), .Z(
        buf_in_last_level_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[1]), .Z(
        buf_in_last_level_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[1]), .Z(
        buf_in_last_level_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[1]), .Z(
        buf_in_last_level_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[2]), .Z(
        buf_in_last_level_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[2]), .Z(
        buf_in_last_level_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[2]), .Z(
        buf_in_last_level_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[2]), .Z(
        buf_in_last_level_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[3]), .Z(
        buf_in_last_level_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[3]), .Z(
        buf_in_last_level_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[3]), .Z(
        buf_in_last_level_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[3]), .Z(
        buf_in_last_level_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[4]), .Z(
        buf_in_last_level_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[4]), .Z(
        buf_in_last_level_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[4]), .Z(
        buf_in_last_level_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[4]), .Z(
        buf_in_last_level_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[5]), .Z(
        buf_in_last_level_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[5]), .Z(
        buf_in_last_level_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[5]), .Z(
        buf_in_last_level_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[5]), .Z(
        buf_in_last_level_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[6]), .Z(
        buf_in_last_level_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[6]), .Z(
        buf_in_last_level_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[6]), .Z(
        buf_in_last_level_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[6]), .Z(
        buf_in_last_level_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[7]), .Z(
        buf_in_last_level_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[7]), .Z(
        buf_in_last_level_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[7]), .Z(
        buf_in_last_level_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[7]), .Z(
        buf_in_last_level_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[8]), .Z(
        buf_in_last_level_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[8]), .Z(
        buf_in_last_level_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[8]), .Z(
        buf_in_last_level_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[8]), .Z(
        buf_in_last_level_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[9]), .Z(
        buf_in_last_level_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[9]), .Z(
        buf_in_last_level_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[9]), .Z(
        buf_in_last_level_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[9]), .Z(
        buf_in_last_level_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[10]), .Z(
        buf_in_last_level_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[10]), .Z(
        buf_in_last_level_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[10]), .Z(
        buf_in_last_level_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[10]), .Z(
        buf_in_last_level_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[11]), .Z(
        buf_in_last_level_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[11]), .Z(
        buf_in_last_level_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[11]), .Z(
        buf_in_last_level_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[11]), .Z(
        buf_in_last_level_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[12]), .Z(
        buf_in_last_level_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[12]), .Z(
        buf_in_last_level_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[12]), .Z(
        buf_in_last_level_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[12]), .Z(
        buf_in_last_level_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[13]), .Z(
        buf_in_last_level_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[13]), .Z(
        buf_in_last_level_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[13]), .Z(
        buf_in_last_level_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[13]), .Z(
        buf_in_last_level_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[14]), .Z(
        buf_in_last_level_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[14]), .Z(
        buf_in_last_level_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[14]), .Z(
        buf_in_last_level_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[14]), .Z(
        buf_in_last_level_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[15]), .Z(
        buf_in_last_level_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[15]), .Z(
        buf_in_last_level_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[15]), .Z(
        buf_in_last_level_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[15]), .Z(
        buf_in_last_level_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[16]), .Z(
        buf_in_last_level_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[16]), .Z(
        buf_in_last_level_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[16]), .Z(
        buf_in_last_level_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[16]), .Z(
        buf_in_last_level_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[17]), .Z(
        buf_in_last_level_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[17]), .Z(
        buf_in_last_level_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[17]), .Z(
        buf_in_last_level_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[17]), .Z(
        buf_in_last_level_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[18]), .Z(
        buf_in_last_level_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[18]), .Z(
        buf_in_last_level_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[18]), .Z(
        buf_in_last_level_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[18]), .Z(
        buf_in_last_level_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[19]), .Z(
        buf_in_last_level_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[19]), .Z(
        buf_in_last_level_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[19]), .Z(
        buf_in_last_level_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[19]), .Z(
        buf_in_last_level_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[20]), .Z(
        buf_in_last_level_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[20]), .Z(
        buf_in_last_level_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[20]), .Z(
        buf_in_last_level_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[20]), .Z(
        buf_in_last_level_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[21]), .Z(
        buf_in_last_level_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[21]), .Z(
        buf_in_last_level_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[21]), .Z(
        buf_in_last_level_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[21]), .Z(
        buf_in_last_level_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[22]), .Z(
        buf_in_last_level_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[22]), .Z(
        buf_in_last_level_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[22]), .Z(
        buf_in_last_level_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[22]), .Z(
        buf_in_last_level_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[23]), .Z(
        buf_in_last_level_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[23]), .Z(
        buf_in_last_level_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[23]), .Z(
        buf_in_last_level_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[23]), .Z(
        buf_in_last_level_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[24]), .Z(
        buf_in_last_level_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[24]), .Z(
        buf_in_last_level_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[24]), .Z(
        buf_in_last_level_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[24]), .Z(
        buf_in_last_level_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[25]), .Z(
        buf_in_last_level_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[25]), .Z(
        buf_in_last_level_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[25]), .Z(
        buf_in_last_level_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[25]), .Z(
        buf_in_last_level_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[26]), .Z(
        buf_in_last_level_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[26]), .Z(
        buf_in_last_level_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[26]), .Z(
        buf_in_last_level_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[26]), .Z(
        buf_in_last_level_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[27]), .Z(
        buf_in_last_level_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[27]), .Z(
        buf_in_last_level_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[27]), .Z(
        buf_in_last_level_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[27]), .Z(
        buf_in_last_level_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[28]), .Z(
        buf_in_last_level_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[28]), .Z(
        buf_in_last_level_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[28]), .Z(
        buf_in_last_level_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[28]), .Z(
        buf_in_last_level_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[29]), .Z(
        buf_in_last_level_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[29]), .Z(
        buf_in_last_level_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[29]), .Z(
        buf_in_last_level_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[29]), .Z(
        buf_in_last_level_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[30]), .Z(
        buf_in_last_level_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[30]), .Z(
        buf_in_last_level_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[30]), .Z(
        buf_in_last_level_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[30]), .Z(
        buf_in_last_level_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[31]), .Z(
        buf_in_last_level_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[31]), .Z(
        buf_in_last_level_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[31]), .Z(
        buf_in_last_level_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[31]), .Z(
        buf_in_last_level_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[32]), .Z(
        buf_in_last_level_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[32]), .Z(
        buf_in_last_level_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[32]), .Z(
        buf_in_last_level_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[32]), .Z(
        buf_in_last_level_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[33]), .Z(
        buf_in_last_level_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[33]), .Z(
        buf_in_last_level_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[33]), .Z(
        buf_in_last_level_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[33]), .Z(
        buf_in_last_level_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[34]), .Z(
        buf_in_last_level_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[34]), .Z(
        buf_in_last_level_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[34]), .Z(
        buf_in_last_level_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[34]), .Z(
        buf_in_last_level_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[35]), .Z(
        buf_in_last_level_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[35]), .Z(
        buf_in_last_level_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[35]), .Z(
        buf_in_last_level_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[35]), .Z(
        buf_in_last_level_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[36]), .Z(
        buf_in_last_level_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[36]), .Z(
        buf_in_last_level_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[36]), .Z(
        buf_in_last_level_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[36]), .Z(
        buf_in_last_level_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[37]), .Z(
        buf_in_last_level_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[37]), .Z(
        buf_in_last_level_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[37]), .Z(
        buf_in_last_level_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[37]), .Z(
        buf_in_last_level_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[38]), .Z(
        buf_in_last_level_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[38]), .Z(
        buf_in_last_level_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[38]), .Z(
        buf_in_last_level_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[38]), .Z(
        buf_in_last_level_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[39]), .Z(
        buf_in_last_level_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[39]), .Z(
        buf_in_last_level_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[39]), .Z(
        buf_in_last_level_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[39]), .Z(
        buf_in_last_level_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[40]), .Z(
        buf_in_last_level_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[40]), .Z(
        buf_in_last_level_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[40]), .Z(
        buf_in_last_level_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[40]), .Z(
        buf_in_last_level_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[41]), .Z(
        buf_in_last_level_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[41]), .Z(
        buf_in_last_level_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[41]), .Z(
        buf_in_last_level_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[41]), .Z(
        buf_in_last_level_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[42]), .Z(
        buf_in_last_level_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[42]), .Z(
        buf_in_last_level_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[42]), .Z(
        buf_in_last_level_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[42]), .Z(
        buf_in_last_level_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[43]), .Z(
        buf_in_last_level_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[43]), .Z(
        buf_in_last_level_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[43]), .Z(
        buf_in_last_level_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[43]), .Z(
        buf_in_last_level_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[44]), .Z(
        buf_in_last_level_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[44]), .Z(
        buf_in_last_level_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[44]), .Z(
        buf_in_last_level_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[44]), .Z(
        buf_in_last_level_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[45]), .Z(
        buf_in_last_level_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[45]), .Z(
        buf_in_last_level_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[45]), .Z(
        buf_in_last_level_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[45]), .Z(
        buf_in_last_level_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[46]), .Z(
        buf_in_last_level_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[46]), .Z(
        buf_in_last_level_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[46]), .Z(
        buf_in_last_level_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[46]), .Z(
        buf_in_last_level_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[47]), .Z(
        buf_in_last_level_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[47]), .Z(
        buf_in_last_level_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[47]), .Z(
        buf_in_last_level_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[47]), .Z(
        buf_in_last_level_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[48]), .Z(
        buf_in_last_level_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[48]), .Z(
        buf_in_last_level_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[48]), .Z(
        buf_in_last_level_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[48]), .Z(
        buf_in_last_level_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[49]), .Z(
        buf_in_last_level_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[49]), .Z(
        buf_in_last_level_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[49]), .Z(
        buf_in_last_level_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[49]), .Z(
        buf_in_last_level_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[50]), .Z(
        buf_in_last_level_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[50]), .Z(
        buf_in_last_level_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[50]), .Z(
        buf_in_last_level_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[50]), .Z(
        buf_in_last_level_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[51]), .Z(
        buf_in_last_level_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[51]), .Z(
        buf_in_last_level_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[51]), .Z(
        buf_in_last_level_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[51]), .Z(
        buf_in_last_level_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[52]), .Z(
        buf_in_last_level_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[52]), .Z(
        buf_in_last_level_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[52]), .Z(
        buf_in_last_level_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[52]), .Z(
        buf_in_last_level_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[53]), .Z(
        buf_in_last_level_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[53]), .Z(
        buf_in_last_level_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[53]), .Z(
        buf_in_last_level_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[53]), .Z(
        buf_in_last_level_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[54]), .Z(
        buf_in_last_level_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[54]), .Z(
        buf_in_last_level_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[54]), .Z(
        buf_in_last_level_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[54]), .Z(
        buf_in_last_level_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[55]), .Z(
        buf_in_last_level_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[55]), .Z(
        buf_in_last_level_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[55]), .Z(
        buf_in_last_level_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[55]), .Z(
        buf_in_last_level_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[56]), .Z(
        buf_in_last_level_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[56]), .Z(
        buf_in_last_level_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[56]), .Z(
        buf_in_last_level_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[56]), .Z(
        buf_in_last_level_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[57]), .Z(
        buf_in_last_level_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[57]), .Z(
        buf_in_last_level_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[57]), .Z(
        buf_in_last_level_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[57]), .Z(
        buf_in_last_level_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[58]), .Z(
        buf_in_last_level_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[58]), .Z(
        buf_in_last_level_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[58]), .Z(
        buf_in_last_level_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[58]), .Z(
        buf_in_last_level_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[59]), .Z(
        buf_in_last_level_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[59]), .Z(
        buf_in_last_level_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[59]), .Z(
        buf_in_last_level_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[59]), .Z(
        buf_in_last_level_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[60]), .Z(
        buf_in_last_level_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[60]), .Z(
        buf_in_last_level_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[60]), .Z(
        buf_in_last_level_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[60]), .Z(
        buf_in_last_level_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[61]), .Z(
        buf_in_last_level_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[61]), .Z(
        buf_in_last_level_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[61]), .Z(
        buf_in_last_level_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[61]), .Z(
        buf_in_last_level_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[62]), .Z(
        buf_in_last_level_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[62]), .Z(
        buf_in_last_level_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[62]), .Z(
        buf_in_last_level_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[62]), .Z(
        buf_in_last_level_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[63]), .Z(
        buf_in_last_level_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[63]), .Z(
        buf_in_last_level_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[63]), .Z(
        buf_in_last_level_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[63]), .Z(
        buf_in_last_level_3__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[64]), .Z(
        buf_in_last_level_0__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[64]), .Z(
        buf_in_last_level_1__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[64]), .Z(
        buf_in_last_level_2__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[64]), .Z(
        buf_in_last_level_3__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[65]), .Z(
        buf_in_last_level_0__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[65]), .Z(
        buf_in_last_level_1__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[65]), .Z(
        buf_in_last_level_2__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[65]), .Z(
        buf_in_last_level_3__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[66]), .Z(
        buf_in_last_level_0__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[66]), .Z(
        buf_in_last_level_1__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[66]), .Z(
        buf_in_last_level_2__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[66]), .Z(
        buf_in_last_level_3__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[67]), .Z(
        buf_in_last_level_0__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[67]), .Z(
        buf_in_last_level_1__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[67]), .Z(
        buf_in_last_level_2__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[67]), .Z(
        buf_in_last_level_3__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[68]), .Z(
        buf_in_last_level_0__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[68]), .Z(
        buf_in_last_level_1__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[68]), .Z(
        buf_in_last_level_2__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[68]), .Z(
        buf_in_last_level_3__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[69]), .Z(
        buf_in_last_level_0__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[69]), .Z(
        buf_in_last_level_1__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[69]), .Z(
        buf_in_last_level_2__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[69]), .Z(
        buf_in_last_level_3__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[70]), .Z(
        buf_in_last_level_0__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[70]), .Z(
        buf_in_last_level_1__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[70]), .Z(
        buf_in_last_level_2__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[70]), .Z(
        buf_in_last_level_3__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[71]), .Z(
        buf_in_last_level_0__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[71]), .Z(
        buf_in_last_level_1__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[71]), .Z(
        buf_in_last_level_2__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[71]), .Z(
        buf_in_last_level_3__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[72]), .Z(
        buf_in_last_level_0__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[72]), .Z(
        buf_in_last_level_1__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[72]), .Z(
        buf_in_last_level_2__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[72]), .Z(
        buf_in_last_level_3__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[73]), .Z(
        buf_in_last_level_0__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[73]), .Z(
        buf_in_last_level_1__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[73]), .Z(
        buf_in_last_level_2__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[73]), .Z(
        buf_in_last_level_3__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[74]), .Z(
        buf_in_last_level_0__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[74]), .Z(
        buf_in_last_level_1__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[74]), .Z(
        buf_in_last_level_2__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[74]), .Z(
        buf_in_last_level_3__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[75]), .Z(
        buf_in_last_level_0__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[75]), .Z(
        buf_in_last_level_1__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[75]), .Z(
        buf_in_last_level_2__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[75]), .Z(
        buf_in_last_level_3__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[76]), .Z(
        buf_in_last_level_0__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[76]), .Z(
        buf_in_last_level_1__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[76]), .Z(
        buf_in_last_level_2__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[76]), .Z(
        buf_in_last_level_3__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[77]), .Z(
        buf_in_last_level_0__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[77]), .Z(
        buf_in_last_level_1__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[77]), .Z(
        buf_in_last_level_2__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[77]), .Z(
        buf_in_last_level_3__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[78]), .Z(
        buf_in_last_level_0__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[78]), .Z(
        buf_in_last_level_1__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[78]), .Z(
        buf_in_last_level_2__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[78]), .Z(
        buf_in_last_level_3__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[79]), .Z(
        buf_in_last_level_0__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[79]), .Z(
        buf_in_last_level_1__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[79]), .Z(
        buf_in_last_level_2__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[79]), .Z(
        buf_in_last_level_3__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[80]), .Z(
        buf_in_last_level_0__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[80]), .Z(
        buf_in_last_level_1__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[80]), .Z(
        buf_in_last_level_2__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[80]), .Z(
        buf_in_last_level_3__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[81]), .Z(
        buf_in_last_level_0__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[81]), .Z(
        buf_in_last_level_1__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[81]), .Z(
        buf_in_last_level_2__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[81]), .Z(
        buf_in_last_level_3__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[82]), .Z(
        buf_in_last_level_0__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[82]), .Z(
        buf_in_last_level_1__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[82]), .Z(
        buf_in_last_level_2__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[82]), .Z(
        buf_in_last_level_3__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[83]), .Z(
        buf_in_last_level_0__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[83]), .Z(
        buf_in_last_level_1__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[83]), .Z(
        buf_in_last_level_2__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[83]), .Z(
        buf_in_last_level_3__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[84]), .Z(
        buf_in_last_level_0__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[84]), .Z(
        buf_in_last_level_1__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[84]), .Z(
        buf_in_last_level_2__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[84]), .Z(
        buf_in_last_level_3__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[85]), .Z(
        buf_in_last_level_0__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[85]), .Z(
        buf_in_last_level_1__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[85]), .Z(
        buf_in_last_level_2__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[85]), .Z(
        buf_in_last_level_3__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[86]), .Z(
        buf_in_last_level_0__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[86]), .Z(
        buf_in_last_level_1__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[86]), .Z(
        buf_in_last_level_2__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[86]), .Z(
        buf_in_last_level_3__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[87]), .Z(
        buf_in_last_level_0__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[87]), .Z(
        buf_in_last_level_1__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[87]), .Z(
        buf_in_last_level_2__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[87]), .Z(
        buf_in_last_level_3__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[88]), .Z(
        buf_in_last_level_0__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[88]), .Z(
        buf_in_last_level_1__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[88]), .Z(
        buf_in_last_level_2__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[88]), .Z(
        buf_in_last_level_3__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[89]), .Z(
        buf_in_last_level_0__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[89]), .Z(
        buf_in_last_level_1__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[89]), .Z(
        buf_in_last_level_2__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[89]), .Z(
        buf_in_last_level_3__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[90]), .Z(
        buf_in_last_level_0__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[90]), .Z(
        buf_in_last_level_1__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[90]), .Z(
        buf_in_last_level_2__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[90]), .Z(
        buf_in_last_level_3__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[91]), .Z(
        buf_in_last_level_0__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[91]), .Z(
        buf_in_last_level_1__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[91]), .Z(
        buf_in_last_level_2__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[91]), .Z(
        buf_in_last_level_3__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[92]), .Z(
        buf_in_last_level_0__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[92]), .Z(
        buf_in_last_level_1__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[92]), .Z(
        buf_in_last_level_2__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[92]), .Z(
        buf_in_last_level_3__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[93]), .Z(
        buf_in_last_level_0__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[93]), .Z(
        buf_in_last_level_1__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[93]), .Z(
        buf_in_last_level_2__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[93]), .Z(
        buf_in_last_level_3__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[94]), .Z(
        buf_in_last_level_0__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[94]), .Z(
        buf_in_last_level_1__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[94]), .Z(
        buf_in_last_level_2__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[94]), .Z(
        buf_in_last_level_3__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[95]), .Z(
        buf_in_last_level_0__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[95]), .Z(
        buf_in_last_level_1__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[95]), .Z(
        buf_in_last_level_2__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[95]), .Z(
        buf_in_last_level_3__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[96]), .Z(
        buf_in_last_level_0__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[96]), .Z(
        buf_in_last_level_1__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[96]), .Z(
        buf_in_last_level_2__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[96]), .Z(
        buf_in_last_level_3__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[97]), .Z(
        buf_in_last_level_0__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[97]), .Z(
        buf_in_last_level_1__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[97]), .Z(
        buf_in_last_level_2__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[97]), .Z(
        buf_in_last_level_3__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[98]), .Z(
        buf_in_last_level_0__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[98]), .Z(
        buf_in_last_level_1__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[98]), .Z(
        buf_in_last_level_2__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[98]), .Z(
        buf_in_last_level_3__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[99]), .Z(
        buf_in_last_level_0__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[99]), .Z(
        buf_in_last_level_1__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[99]), .Z(
        buf_in_last_level_2__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[99]), .Z(
        buf_in_last_level_3__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[100]), .Z(
        buf_in_last_level_0__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[100]), .Z(
        buf_in_last_level_1__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[100]), .Z(
        buf_in_last_level_2__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[100]), .Z(
        buf_in_last_level_3__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[101]), .Z(
        buf_in_last_level_0__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[101]), .Z(
        buf_in_last_level_1__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[101]), .Z(
        buf_in_last_level_2__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[101]), .Z(
        buf_in_last_level_3__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[102]), .Z(
        buf_in_last_level_0__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[102]), .Z(
        buf_in_last_level_1__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[102]), .Z(
        buf_in_last_level_2__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[102]), .Z(
        buf_in_last_level_3__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[103]), .Z(
        buf_in_last_level_0__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[103]), .Z(
        buf_in_last_level_1__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[103]), .Z(
        buf_in_last_level_2__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[103]), .Z(
        buf_in_last_level_3__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[104]), .Z(
        buf_in_last_level_0__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[104]), .Z(
        buf_in_last_level_1__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[104]), .Z(
        buf_in_last_level_2__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[104]), .Z(
        buf_in_last_level_3__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[105]), .Z(
        buf_in_last_level_0__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[105]), .Z(
        buf_in_last_level_1__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[105]), .Z(
        buf_in_last_level_2__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[105]), .Z(
        buf_in_last_level_3__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[106]), .Z(
        buf_in_last_level_0__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[106]), .Z(
        buf_in_last_level_1__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[106]), .Z(
        buf_in_last_level_2__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[106]), .Z(
        buf_in_last_level_3__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[107]), .Z(
        buf_in_last_level_0__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[107]), .Z(
        buf_in_last_level_1__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[107]), .Z(
        buf_in_last_level_2__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[107]), .Z(
        buf_in_last_level_3__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[108]), .Z(
        buf_in_last_level_0__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[108]), .Z(
        buf_in_last_level_1__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[108]), .Z(
        buf_in_last_level_2__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[108]), .Z(
        buf_in_last_level_3__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[109]), .Z(
        buf_in_last_level_0__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[109]), .Z(
        buf_in_last_level_1__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[109]), .Z(
        buf_in_last_level_2__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[109]), .Z(
        buf_in_last_level_3__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[110]), .Z(
        buf_in_last_level_0__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[110]), .Z(
        buf_in_last_level_1__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[110]), .Z(
        buf_in_last_level_2__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[110]), .Z(
        buf_in_last_level_3__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[111]), .Z(
        buf_in_last_level_0__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[111]), .Z(
        buf_in_last_level_1__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[111]), .Z(
        buf_in_last_level_2__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[111]), .Z(
        buf_in_last_level_3__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[112]), .Z(
        buf_in_last_level_0__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[112]), .Z(
        buf_in_last_level_1__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[112]), .Z(
        buf_in_last_level_2__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[112]), .Z(
        buf_in_last_level_3__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[113]), .Z(
        buf_in_last_level_0__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[113]), .Z(
        buf_in_last_level_1__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[113]), .Z(
        buf_in_last_level_2__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[113]), .Z(
        buf_in_last_level_3__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[114]), .Z(
        buf_in_last_level_0__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[114]), .Z(
        buf_in_last_level_1__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[114]), .Z(
        buf_in_last_level_2__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[114]), .Z(
        buf_in_last_level_3__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[115]), .Z(
        buf_in_last_level_0__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[115]), .Z(
        buf_in_last_level_1__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[115]), .Z(
        buf_in_last_level_2__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[115]), .Z(
        buf_in_last_level_3__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[116]), .Z(
        buf_in_last_level_0__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[116]), .Z(
        buf_in_last_level_1__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[116]), .Z(
        buf_in_last_level_2__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[116]), .Z(
        buf_in_last_level_3__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[117]), .Z(
        buf_in_last_level_0__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[117]), .Z(
        buf_in_last_level_1__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[117]), .Z(
        buf_in_last_level_2__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[117]), .Z(
        buf_in_last_level_3__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[118]), .Z(
        buf_in_last_level_0__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[118]), .Z(
        buf_in_last_level_1__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[118]), .Z(
        buf_in_last_level_2__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[118]), .Z(
        buf_in_last_level_3__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[119]), .Z(
        buf_in_last_level_0__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[119]), .Z(
        buf_in_last_level_1__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[119]), .Z(
        buf_in_last_level_2__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[119]), .Z(
        buf_in_last_level_3__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[120]), .Z(
        buf_in_last_level_0__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[120]), .Z(
        buf_in_last_level_1__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[120]), .Z(
        buf_in_last_level_2__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[120]), .Z(
        buf_in_last_level_3__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[121]), .Z(
        buf_in_last_level_0__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[121]), .Z(
        buf_in_last_level_1__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[121]), .Z(
        buf_in_last_level_2__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[121]), .Z(
        buf_in_last_level_3__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[122]), .Z(
        buf_in_last_level_0__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[122]), .Z(
        buf_in_last_level_1__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[122]), .Z(
        buf_in_last_level_2__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[122]), .Z(
        buf_in_last_level_3__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[123]), .Z(
        buf_in_last_level_0__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[123]), .Z(
        buf_in_last_level_1__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[123]), .Z(
        buf_in_last_level_2__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[123]), .Z(
        buf_in_last_level_3__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[124]), .Z(
        buf_in_last_level_0__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[124]), .Z(
        buf_in_last_level_1__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[124]), .Z(
        buf_in_last_level_2__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[124]), .Z(
        buf_in_last_level_3__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[125]), .Z(
        buf_in_last_level_0__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[125]), .Z(
        buf_in_last_level_1__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[125]), .Z(
        buf_in_last_level_2__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[125]), .Z(
        buf_in_last_level_3__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[126]), .Z(
        buf_in_last_level_0__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[126]), .Z(
        buf_in_last_level_1__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[126]), .Z(
        buf_in_last_level_2__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[126]), .Z(
        buf_in_last_level_3__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[127]), .Z(
        buf_in_last_level_0__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[127]), .Z(
        buf_in_last_level_1__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[127]), .Z(
        buf_in_last_level_2__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[127]), .Z(
        buf_in_last_level_3__i_data_o_buf[127]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(CLK), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(CLK), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(CLK), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(CLK), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(CLK), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(CLK), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(CLK), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(CLK), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[101]), .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[102]), .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[105]), .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[107]), .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[109]), .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[110]), .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[111]), .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[112]), .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[115]), .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[82]), .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[86]), .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[61]), .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[63]), .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[31]), .Z(N297) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[23]), .Z(N289) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[24]), .Z(N290) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[25]), .Z(N291) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[21]), .Z(N287) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[30]), .Z(N296) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[20]), .Z(N286) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[26]), .Z(N292) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[22]), .Z(N288) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[28]), .Z(N294) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[29]), .Z(N295) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[27]), .Z(N293) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[19]), .Z(N285) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[18]), .Z(N284) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[16]), .Z(N282) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[15]), .Z(N281) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[14]), .Z(N280) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[13]), .Z(N279) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[12]), .Z(N278) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[11]), .Z(N277) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[10]), .Z(N276) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[9]), .Z(N275) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[8]), .Z(N274) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[7]), .Z(N273) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[5]), .Z(N271) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[4]), .Z(N270) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[3]), .Z(N269) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[1]), .Z(N267) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[0]), .Z(N266) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[62]), .Z(N362) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[60]), .Z(N360) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[59]), .Z(N359) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[58]), .Z(N358) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[57]), .Z(N357) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[56]), .Z(N356) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[55]), .Z(N355) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[54]), .Z(N354) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[53]), .Z(N353) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[52]), .Z(N352) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[51]), .Z(N351) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[50]), .Z(N350) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[49]), .Z(N349) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[48]), .Z(N348) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[47]), .Z(N347) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[46]), .Z(N346) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[45]), .Z(N345) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[44]), .Z(N344) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[43]), .Z(N343) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[42]), .Z(N342) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[41]), .Z(N341) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[40]), .Z(N340) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[17]), .Z(N283) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[39]), .Z(N339) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[38]), .Z(N338) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[37]), .Z(N337) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[36]), .Z(N336) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[64]), .Z(N398) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[65]), .Z(N399) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[66]), .Z(N400) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[67]), .Z(N401) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[68]), .Z(N402) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[69]), .Z(N403) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[70]), .Z(N404) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[71]), .Z(N405) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[72]), .Z(N406) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[73]), .Z(N407) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[74]), .Z(N408) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[75]), .Z(N409) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[76]), .Z(N410) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[77]), .Z(N411) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[78]), .Z(N412) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[79]), .Z(N413) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[80]), .Z(N414) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[81]), .Z(N415) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[83]), .Z(N417) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[84]), .Z(N418) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[85]), .Z(N419) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[87]), .Z(N421) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[88]), .Z(N422) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[89]), .Z(N423) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[90]), .Z(N424) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[91]), .Z(N425) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[92]), .Z(N426) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[93]), .Z(N427) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[94]), .Z(N428) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[95]), .Z(N429) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[32]), .Z(N332) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[33]), .Z(N333) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[34]), .Z(N334) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[35]), .Z(N335) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        CLK, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input CLK, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;
  wire   [127:0] buf_in_last_level_0__i_data_o_buf;
  wire   [127:0] buf_in_last_level_1__i_data_o_buf;
  wire   [127:0] buf_in_last_level_2__i_data_o_buf;
  wire   [127:0] buf_in_last_level_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[0]), .Z(
        buf_in_last_level_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[0]), .Z(
        buf_in_last_level_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[0]), .Z(
        buf_in_last_level_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[0]), .Z(
        buf_in_last_level_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[1]), .Z(
        buf_in_last_level_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[1]), .Z(
        buf_in_last_level_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[1]), .Z(
        buf_in_last_level_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[1]), .Z(
        buf_in_last_level_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[2]), .Z(
        buf_in_last_level_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[2]), .Z(
        buf_in_last_level_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[2]), .Z(
        buf_in_last_level_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[2]), .Z(
        buf_in_last_level_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[3]), .Z(
        buf_in_last_level_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[3]), .Z(
        buf_in_last_level_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[3]), .Z(
        buf_in_last_level_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[3]), .Z(
        buf_in_last_level_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[4]), .Z(
        buf_in_last_level_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[4]), .Z(
        buf_in_last_level_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[4]), .Z(
        buf_in_last_level_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[4]), .Z(
        buf_in_last_level_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[5]), .Z(
        buf_in_last_level_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[5]), .Z(
        buf_in_last_level_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[5]), .Z(
        buf_in_last_level_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[5]), .Z(
        buf_in_last_level_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[6]), .Z(
        buf_in_last_level_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[6]), .Z(
        buf_in_last_level_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[6]), .Z(
        buf_in_last_level_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[6]), .Z(
        buf_in_last_level_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[7]), .Z(
        buf_in_last_level_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[7]), .Z(
        buf_in_last_level_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[7]), .Z(
        buf_in_last_level_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[7]), .Z(
        buf_in_last_level_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[8]), .Z(
        buf_in_last_level_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[8]), .Z(
        buf_in_last_level_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[8]), .Z(
        buf_in_last_level_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[8]), .Z(
        buf_in_last_level_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[9]), .Z(
        buf_in_last_level_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[9]), .Z(
        buf_in_last_level_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[9]), .Z(
        buf_in_last_level_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[9]), .Z(
        buf_in_last_level_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[10]), .Z(
        buf_in_last_level_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[10]), .Z(
        buf_in_last_level_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[10]), .Z(
        buf_in_last_level_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[10]), .Z(
        buf_in_last_level_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[11]), .Z(
        buf_in_last_level_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[11]), .Z(
        buf_in_last_level_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[11]), .Z(
        buf_in_last_level_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[11]), .Z(
        buf_in_last_level_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[12]), .Z(
        buf_in_last_level_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[12]), .Z(
        buf_in_last_level_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[12]), .Z(
        buf_in_last_level_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[12]), .Z(
        buf_in_last_level_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[13]), .Z(
        buf_in_last_level_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[13]), .Z(
        buf_in_last_level_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[13]), .Z(
        buf_in_last_level_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[13]), .Z(
        buf_in_last_level_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[14]), .Z(
        buf_in_last_level_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[14]), .Z(
        buf_in_last_level_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[14]), .Z(
        buf_in_last_level_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[14]), .Z(
        buf_in_last_level_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[15]), .Z(
        buf_in_last_level_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[15]), .Z(
        buf_in_last_level_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[15]), .Z(
        buf_in_last_level_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[15]), .Z(
        buf_in_last_level_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[16]), .Z(
        buf_in_last_level_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[16]), .Z(
        buf_in_last_level_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[16]), .Z(
        buf_in_last_level_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[16]), .Z(
        buf_in_last_level_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[17]), .Z(
        buf_in_last_level_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[17]), .Z(
        buf_in_last_level_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[17]), .Z(
        buf_in_last_level_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[17]), .Z(
        buf_in_last_level_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[18]), .Z(
        buf_in_last_level_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[18]), .Z(
        buf_in_last_level_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[18]), .Z(
        buf_in_last_level_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[18]), .Z(
        buf_in_last_level_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[19]), .Z(
        buf_in_last_level_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[19]), .Z(
        buf_in_last_level_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[19]), .Z(
        buf_in_last_level_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[19]), .Z(
        buf_in_last_level_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[20]), .Z(
        buf_in_last_level_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[20]), .Z(
        buf_in_last_level_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[20]), .Z(
        buf_in_last_level_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[20]), .Z(
        buf_in_last_level_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[21]), .Z(
        buf_in_last_level_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[21]), .Z(
        buf_in_last_level_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[21]), .Z(
        buf_in_last_level_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[21]), .Z(
        buf_in_last_level_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[22]), .Z(
        buf_in_last_level_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[22]), .Z(
        buf_in_last_level_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[22]), .Z(
        buf_in_last_level_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[22]), .Z(
        buf_in_last_level_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[23]), .Z(
        buf_in_last_level_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[23]), .Z(
        buf_in_last_level_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[23]), .Z(
        buf_in_last_level_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[23]), .Z(
        buf_in_last_level_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[24]), .Z(
        buf_in_last_level_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[24]), .Z(
        buf_in_last_level_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[24]), .Z(
        buf_in_last_level_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[24]), .Z(
        buf_in_last_level_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[25]), .Z(
        buf_in_last_level_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[25]), .Z(
        buf_in_last_level_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[25]), .Z(
        buf_in_last_level_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[25]), .Z(
        buf_in_last_level_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[26]), .Z(
        buf_in_last_level_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[26]), .Z(
        buf_in_last_level_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[26]), .Z(
        buf_in_last_level_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[26]), .Z(
        buf_in_last_level_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[27]), .Z(
        buf_in_last_level_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[27]), .Z(
        buf_in_last_level_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[27]), .Z(
        buf_in_last_level_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[27]), .Z(
        buf_in_last_level_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[28]), .Z(
        buf_in_last_level_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[28]), .Z(
        buf_in_last_level_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[28]), .Z(
        buf_in_last_level_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[28]), .Z(
        buf_in_last_level_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[29]), .Z(
        buf_in_last_level_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[29]), .Z(
        buf_in_last_level_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[29]), .Z(
        buf_in_last_level_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[29]), .Z(
        buf_in_last_level_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[30]), .Z(
        buf_in_last_level_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[30]), .Z(
        buf_in_last_level_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[30]), .Z(
        buf_in_last_level_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[30]), .Z(
        buf_in_last_level_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[31]), .Z(
        buf_in_last_level_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[31]), .Z(
        buf_in_last_level_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[31]), .Z(
        buf_in_last_level_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[31]), .Z(
        buf_in_last_level_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[32]), .Z(
        buf_in_last_level_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[32]), .Z(
        buf_in_last_level_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[32]), .Z(
        buf_in_last_level_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[32]), .Z(
        buf_in_last_level_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[33]), .Z(
        buf_in_last_level_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[33]), .Z(
        buf_in_last_level_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[33]), .Z(
        buf_in_last_level_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[33]), .Z(
        buf_in_last_level_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[34]), .Z(
        buf_in_last_level_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[34]), .Z(
        buf_in_last_level_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[34]), .Z(
        buf_in_last_level_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[34]), .Z(
        buf_in_last_level_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[35]), .Z(
        buf_in_last_level_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[35]), .Z(
        buf_in_last_level_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[35]), .Z(
        buf_in_last_level_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[35]), .Z(
        buf_in_last_level_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[36]), .Z(
        buf_in_last_level_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[36]), .Z(
        buf_in_last_level_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[36]), .Z(
        buf_in_last_level_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[36]), .Z(
        buf_in_last_level_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[37]), .Z(
        buf_in_last_level_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[37]), .Z(
        buf_in_last_level_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[37]), .Z(
        buf_in_last_level_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[37]), .Z(
        buf_in_last_level_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[38]), .Z(
        buf_in_last_level_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[38]), .Z(
        buf_in_last_level_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[38]), .Z(
        buf_in_last_level_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[38]), .Z(
        buf_in_last_level_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[39]), .Z(
        buf_in_last_level_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[39]), .Z(
        buf_in_last_level_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[39]), .Z(
        buf_in_last_level_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[39]), .Z(
        buf_in_last_level_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[40]), .Z(
        buf_in_last_level_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[40]), .Z(
        buf_in_last_level_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[40]), .Z(
        buf_in_last_level_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[40]), .Z(
        buf_in_last_level_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[41]), .Z(
        buf_in_last_level_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[41]), .Z(
        buf_in_last_level_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[41]), .Z(
        buf_in_last_level_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[41]), .Z(
        buf_in_last_level_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[42]), .Z(
        buf_in_last_level_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[42]), .Z(
        buf_in_last_level_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[42]), .Z(
        buf_in_last_level_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[42]), .Z(
        buf_in_last_level_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[43]), .Z(
        buf_in_last_level_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[43]), .Z(
        buf_in_last_level_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[43]), .Z(
        buf_in_last_level_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[43]), .Z(
        buf_in_last_level_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[44]), .Z(
        buf_in_last_level_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[44]), .Z(
        buf_in_last_level_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[44]), .Z(
        buf_in_last_level_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[44]), .Z(
        buf_in_last_level_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[45]), .Z(
        buf_in_last_level_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[45]), .Z(
        buf_in_last_level_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[45]), .Z(
        buf_in_last_level_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[45]), .Z(
        buf_in_last_level_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[46]), .Z(
        buf_in_last_level_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[46]), .Z(
        buf_in_last_level_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[46]), .Z(
        buf_in_last_level_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[46]), .Z(
        buf_in_last_level_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[47]), .Z(
        buf_in_last_level_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[47]), .Z(
        buf_in_last_level_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[47]), .Z(
        buf_in_last_level_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[47]), .Z(
        buf_in_last_level_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[48]), .Z(
        buf_in_last_level_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[48]), .Z(
        buf_in_last_level_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[48]), .Z(
        buf_in_last_level_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[48]), .Z(
        buf_in_last_level_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[49]), .Z(
        buf_in_last_level_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[49]), .Z(
        buf_in_last_level_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[49]), .Z(
        buf_in_last_level_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[49]), .Z(
        buf_in_last_level_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[50]), .Z(
        buf_in_last_level_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[50]), .Z(
        buf_in_last_level_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[50]), .Z(
        buf_in_last_level_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[50]), .Z(
        buf_in_last_level_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[51]), .Z(
        buf_in_last_level_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[51]), .Z(
        buf_in_last_level_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[51]), .Z(
        buf_in_last_level_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[51]), .Z(
        buf_in_last_level_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[52]), .Z(
        buf_in_last_level_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[52]), .Z(
        buf_in_last_level_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[52]), .Z(
        buf_in_last_level_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[52]), .Z(
        buf_in_last_level_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[53]), .Z(
        buf_in_last_level_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[53]), .Z(
        buf_in_last_level_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[53]), .Z(
        buf_in_last_level_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[53]), .Z(
        buf_in_last_level_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[54]), .Z(
        buf_in_last_level_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[54]), .Z(
        buf_in_last_level_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[54]), .Z(
        buf_in_last_level_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[54]), .Z(
        buf_in_last_level_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[55]), .Z(
        buf_in_last_level_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[55]), .Z(
        buf_in_last_level_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[55]), .Z(
        buf_in_last_level_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[55]), .Z(
        buf_in_last_level_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[56]), .Z(
        buf_in_last_level_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[56]), .Z(
        buf_in_last_level_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[56]), .Z(
        buf_in_last_level_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[56]), .Z(
        buf_in_last_level_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[57]), .Z(
        buf_in_last_level_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[57]), .Z(
        buf_in_last_level_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[57]), .Z(
        buf_in_last_level_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[57]), .Z(
        buf_in_last_level_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[58]), .Z(
        buf_in_last_level_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[58]), .Z(
        buf_in_last_level_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[58]), .Z(
        buf_in_last_level_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[58]), .Z(
        buf_in_last_level_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[59]), .Z(
        buf_in_last_level_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[59]), .Z(
        buf_in_last_level_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[59]), .Z(
        buf_in_last_level_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[59]), .Z(
        buf_in_last_level_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[60]), .Z(
        buf_in_last_level_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[60]), .Z(
        buf_in_last_level_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[60]), .Z(
        buf_in_last_level_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[60]), .Z(
        buf_in_last_level_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[61]), .Z(
        buf_in_last_level_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[61]), .Z(
        buf_in_last_level_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[61]), .Z(
        buf_in_last_level_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[61]), .Z(
        buf_in_last_level_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[62]), .Z(
        buf_in_last_level_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[62]), .Z(
        buf_in_last_level_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[62]), .Z(
        buf_in_last_level_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[62]), .Z(
        buf_in_last_level_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[63]), .Z(
        buf_in_last_level_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[63]), .Z(
        buf_in_last_level_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[63]), .Z(
        buf_in_last_level_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[63]), .Z(
        buf_in_last_level_3__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[64]), .Z(
        buf_in_last_level_0__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[64]), .Z(
        buf_in_last_level_1__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[64]), .Z(
        buf_in_last_level_2__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[64]), .Z(
        buf_in_last_level_3__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[65]), .Z(
        buf_in_last_level_0__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[65]), .Z(
        buf_in_last_level_1__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[65]), .Z(
        buf_in_last_level_2__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[65]), .Z(
        buf_in_last_level_3__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[66]), .Z(
        buf_in_last_level_0__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[66]), .Z(
        buf_in_last_level_1__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[66]), .Z(
        buf_in_last_level_2__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[66]), .Z(
        buf_in_last_level_3__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[67]), .Z(
        buf_in_last_level_0__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[67]), .Z(
        buf_in_last_level_1__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[67]), .Z(
        buf_in_last_level_2__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[67]), .Z(
        buf_in_last_level_3__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[68]), .Z(
        buf_in_last_level_0__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[68]), .Z(
        buf_in_last_level_1__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[68]), .Z(
        buf_in_last_level_2__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[68]), .Z(
        buf_in_last_level_3__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[69]), .Z(
        buf_in_last_level_0__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[69]), .Z(
        buf_in_last_level_1__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[69]), .Z(
        buf_in_last_level_2__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[69]), .Z(
        buf_in_last_level_3__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[70]), .Z(
        buf_in_last_level_0__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[70]), .Z(
        buf_in_last_level_1__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[70]), .Z(
        buf_in_last_level_2__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[70]), .Z(
        buf_in_last_level_3__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[71]), .Z(
        buf_in_last_level_0__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[71]), .Z(
        buf_in_last_level_1__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[71]), .Z(
        buf_in_last_level_2__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[71]), .Z(
        buf_in_last_level_3__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[72]), .Z(
        buf_in_last_level_0__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[72]), .Z(
        buf_in_last_level_1__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[72]), .Z(
        buf_in_last_level_2__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[72]), .Z(
        buf_in_last_level_3__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[73]), .Z(
        buf_in_last_level_0__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[73]), .Z(
        buf_in_last_level_1__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[73]), .Z(
        buf_in_last_level_2__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[73]), .Z(
        buf_in_last_level_3__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[74]), .Z(
        buf_in_last_level_0__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[74]), .Z(
        buf_in_last_level_1__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[74]), .Z(
        buf_in_last_level_2__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[74]), .Z(
        buf_in_last_level_3__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[75]), .Z(
        buf_in_last_level_0__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[75]), .Z(
        buf_in_last_level_1__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[75]), .Z(
        buf_in_last_level_2__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[75]), .Z(
        buf_in_last_level_3__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[76]), .Z(
        buf_in_last_level_0__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[76]), .Z(
        buf_in_last_level_1__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[76]), .Z(
        buf_in_last_level_2__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[76]), .Z(
        buf_in_last_level_3__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[77]), .Z(
        buf_in_last_level_0__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[77]), .Z(
        buf_in_last_level_1__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[77]), .Z(
        buf_in_last_level_2__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[77]), .Z(
        buf_in_last_level_3__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[78]), .Z(
        buf_in_last_level_0__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[78]), .Z(
        buf_in_last_level_1__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[78]), .Z(
        buf_in_last_level_2__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[78]), .Z(
        buf_in_last_level_3__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[79]), .Z(
        buf_in_last_level_0__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[79]), .Z(
        buf_in_last_level_1__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[79]), .Z(
        buf_in_last_level_2__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[79]), .Z(
        buf_in_last_level_3__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[80]), .Z(
        buf_in_last_level_0__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[80]), .Z(
        buf_in_last_level_1__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[80]), .Z(
        buf_in_last_level_2__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[80]), .Z(
        buf_in_last_level_3__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[81]), .Z(
        buf_in_last_level_0__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[81]), .Z(
        buf_in_last_level_1__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[81]), .Z(
        buf_in_last_level_2__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[81]), .Z(
        buf_in_last_level_3__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[82]), .Z(
        buf_in_last_level_0__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[82]), .Z(
        buf_in_last_level_1__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[82]), .Z(
        buf_in_last_level_2__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[82]), .Z(
        buf_in_last_level_3__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[83]), .Z(
        buf_in_last_level_0__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[83]), .Z(
        buf_in_last_level_1__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[83]), .Z(
        buf_in_last_level_2__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[83]), .Z(
        buf_in_last_level_3__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[84]), .Z(
        buf_in_last_level_0__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[84]), .Z(
        buf_in_last_level_1__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[84]), .Z(
        buf_in_last_level_2__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[84]), .Z(
        buf_in_last_level_3__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[85]), .Z(
        buf_in_last_level_0__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[85]), .Z(
        buf_in_last_level_1__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[85]), .Z(
        buf_in_last_level_2__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[85]), .Z(
        buf_in_last_level_3__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[86]), .Z(
        buf_in_last_level_0__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[86]), .Z(
        buf_in_last_level_1__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[86]), .Z(
        buf_in_last_level_2__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[86]), .Z(
        buf_in_last_level_3__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[87]), .Z(
        buf_in_last_level_0__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[87]), .Z(
        buf_in_last_level_1__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[87]), .Z(
        buf_in_last_level_2__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[87]), .Z(
        buf_in_last_level_3__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[88]), .Z(
        buf_in_last_level_0__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[88]), .Z(
        buf_in_last_level_1__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[88]), .Z(
        buf_in_last_level_2__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[88]), .Z(
        buf_in_last_level_3__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[89]), .Z(
        buf_in_last_level_0__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[89]), .Z(
        buf_in_last_level_1__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[89]), .Z(
        buf_in_last_level_2__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[89]), .Z(
        buf_in_last_level_3__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[90]), .Z(
        buf_in_last_level_0__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[90]), .Z(
        buf_in_last_level_1__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[90]), .Z(
        buf_in_last_level_2__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[90]), .Z(
        buf_in_last_level_3__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[91]), .Z(
        buf_in_last_level_0__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[91]), .Z(
        buf_in_last_level_1__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[91]), .Z(
        buf_in_last_level_2__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[91]), .Z(
        buf_in_last_level_3__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[92]), .Z(
        buf_in_last_level_0__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[92]), .Z(
        buf_in_last_level_1__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[92]), .Z(
        buf_in_last_level_2__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[92]), .Z(
        buf_in_last_level_3__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[93]), .Z(
        buf_in_last_level_0__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[93]), .Z(
        buf_in_last_level_1__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[93]), .Z(
        buf_in_last_level_2__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[93]), .Z(
        buf_in_last_level_3__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[94]), .Z(
        buf_in_last_level_0__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[94]), .Z(
        buf_in_last_level_1__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[94]), .Z(
        buf_in_last_level_2__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[94]), .Z(
        buf_in_last_level_3__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[95]), .Z(
        buf_in_last_level_0__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[95]), .Z(
        buf_in_last_level_1__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[95]), .Z(
        buf_in_last_level_2__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[95]), .Z(
        buf_in_last_level_3__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[96]), .Z(
        buf_in_last_level_0__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[96]), .Z(
        buf_in_last_level_1__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[96]), .Z(
        buf_in_last_level_2__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[96]), .Z(
        buf_in_last_level_3__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[97]), .Z(
        buf_in_last_level_0__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[97]), .Z(
        buf_in_last_level_1__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[97]), .Z(
        buf_in_last_level_2__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[97]), .Z(
        buf_in_last_level_3__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[98]), .Z(
        buf_in_last_level_0__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[98]), .Z(
        buf_in_last_level_1__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[98]), .Z(
        buf_in_last_level_2__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[98]), .Z(
        buf_in_last_level_3__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[99]), .Z(
        buf_in_last_level_0__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[99]), .Z(
        buf_in_last_level_1__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[99]), .Z(
        buf_in_last_level_2__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[99]), .Z(
        buf_in_last_level_3__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[100]), .Z(
        buf_in_last_level_0__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[100]), .Z(
        buf_in_last_level_1__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[100]), .Z(
        buf_in_last_level_2__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[100]), .Z(
        buf_in_last_level_3__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[101]), .Z(
        buf_in_last_level_0__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[101]), .Z(
        buf_in_last_level_1__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[101]), .Z(
        buf_in_last_level_2__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[101]), .Z(
        buf_in_last_level_3__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[102]), .Z(
        buf_in_last_level_0__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[102]), .Z(
        buf_in_last_level_1__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[102]), .Z(
        buf_in_last_level_2__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[102]), .Z(
        buf_in_last_level_3__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[103]), .Z(
        buf_in_last_level_0__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[103]), .Z(
        buf_in_last_level_1__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[103]), .Z(
        buf_in_last_level_2__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[103]), .Z(
        buf_in_last_level_3__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[104]), .Z(
        buf_in_last_level_0__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[104]), .Z(
        buf_in_last_level_1__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[104]), .Z(
        buf_in_last_level_2__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[104]), .Z(
        buf_in_last_level_3__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[105]), .Z(
        buf_in_last_level_0__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[105]), .Z(
        buf_in_last_level_1__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[105]), .Z(
        buf_in_last_level_2__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[105]), .Z(
        buf_in_last_level_3__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[106]), .Z(
        buf_in_last_level_0__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[106]), .Z(
        buf_in_last_level_1__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[106]), .Z(
        buf_in_last_level_2__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[106]), .Z(
        buf_in_last_level_3__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[107]), .Z(
        buf_in_last_level_0__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[107]), .Z(
        buf_in_last_level_1__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[107]), .Z(
        buf_in_last_level_2__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[107]), .Z(
        buf_in_last_level_3__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[108]), .Z(
        buf_in_last_level_0__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[108]), .Z(
        buf_in_last_level_1__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[108]), .Z(
        buf_in_last_level_2__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[108]), .Z(
        buf_in_last_level_3__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[109]), .Z(
        buf_in_last_level_0__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[109]), .Z(
        buf_in_last_level_1__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[109]), .Z(
        buf_in_last_level_2__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[109]), .Z(
        buf_in_last_level_3__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[110]), .Z(
        buf_in_last_level_0__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[110]), .Z(
        buf_in_last_level_1__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[110]), .Z(
        buf_in_last_level_2__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[110]), .Z(
        buf_in_last_level_3__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[111]), .Z(
        buf_in_last_level_0__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[111]), .Z(
        buf_in_last_level_1__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[111]), .Z(
        buf_in_last_level_2__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[111]), .Z(
        buf_in_last_level_3__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[112]), .Z(
        buf_in_last_level_0__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[112]), .Z(
        buf_in_last_level_1__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[112]), .Z(
        buf_in_last_level_2__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[112]), .Z(
        buf_in_last_level_3__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[113]), .Z(
        buf_in_last_level_0__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[113]), .Z(
        buf_in_last_level_1__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[113]), .Z(
        buf_in_last_level_2__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[113]), .Z(
        buf_in_last_level_3__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[114]), .Z(
        buf_in_last_level_0__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[114]), .Z(
        buf_in_last_level_1__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[114]), .Z(
        buf_in_last_level_2__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[114]), .Z(
        buf_in_last_level_3__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[115]), .Z(
        buf_in_last_level_0__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[115]), .Z(
        buf_in_last_level_1__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[115]), .Z(
        buf_in_last_level_2__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[115]), .Z(
        buf_in_last_level_3__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[116]), .Z(
        buf_in_last_level_0__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[116]), .Z(
        buf_in_last_level_1__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[116]), .Z(
        buf_in_last_level_2__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[116]), .Z(
        buf_in_last_level_3__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[117]), .Z(
        buf_in_last_level_0__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[117]), .Z(
        buf_in_last_level_1__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[117]), .Z(
        buf_in_last_level_2__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[117]), .Z(
        buf_in_last_level_3__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[118]), .Z(
        buf_in_last_level_0__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[118]), .Z(
        buf_in_last_level_1__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[118]), .Z(
        buf_in_last_level_2__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[118]), .Z(
        buf_in_last_level_3__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[119]), .Z(
        buf_in_last_level_0__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[119]), .Z(
        buf_in_last_level_1__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[119]), .Z(
        buf_in_last_level_2__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[119]), .Z(
        buf_in_last_level_3__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[120]), .Z(
        buf_in_last_level_0__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[120]), .Z(
        buf_in_last_level_1__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[120]), .Z(
        buf_in_last_level_2__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[120]), .Z(
        buf_in_last_level_3__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[121]), .Z(
        buf_in_last_level_0__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[121]), .Z(
        buf_in_last_level_1__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[121]), .Z(
        buf_in_last_level_2__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[121]), .Z(
        buf_in_last_level_3__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[122]), .Z(
        buf_in_last_level_0__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[122]), .Z(
        buf_in_last_level_1__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[122]), .Z(
        buf_in_last_level_2__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[122]), .Z(
        buf_in_last_level_3__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[123]), .Z(
        buf_in_last_level_0__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[123]), .Z(
        buf_in_last_level_1__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[123]), .Z(
        buf_in_last_level_2__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[123]), .Z(
        buf_in_last_level_3__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[124]), .Z(
        buf_in_last_level_0__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[124]), .Z(
        buf_in_last_level_1__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[124]), .Z(
        buf_in_last_level_2__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[124]), .Z(
        buf_in_last_level_3__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[125]), .Z(
        buf_in_last_level_0__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[125]), .Z(
        buf_in_last_level_1__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[125]), .Z(
        buf_in_last_level_2__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[125]), .Z(
        buf_in_last_level_3__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[126]), .Z(
        buf_in_last_level_0__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[126]), .Z(
        buf_in_last_level_1__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[126]), .Z(
        buf_in_last_level_2__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[126]), .Z(
        buf_in_last_level_3__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[127]), .Z(
        buf_in_last_level_0__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[127]), .Z(
        buf_in_last_level_1__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[127]), .Z(
        buf_in_last_level_2__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[127]), .Z(
        buf_in_last_level_3__i_data_o_buf[127]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(CLK), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(CLK), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(CLK), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(CLK), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(CLK), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(CLK), .Q(o_valid[7]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(CLK), .Q(o_valid[3]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(CLK), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[101]), .Z(N469) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[102]), .Z(N470) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[105]), .Z(N473) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[107]), .Z(N475) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[109]), .Z(N477) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[110]), .Z(N478) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[111]), .Z(N479) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[112]), .Z(N480) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[115]), .Z(N483) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[82]), .Z(N416) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[86]), .Z(N420) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[61]), .Z(N361) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[63]), .Z(N363) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[31]), .Z(N297) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[30]), .Z(N296) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[29]), .Z(N295) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[28]), .Z(N294) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[27]), .Z(N293) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[26]), .Z(N292) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[25]), .Z(N291) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[24]), .Z(N290) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[23]), .Z(N289) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[22]), .Z(N288) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[21]), .Z(N287) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[20]), .Z(N286) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[18]), .Z(N284) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[17]), .Z(N283) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[16]), .Z(N282) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[15]), .Z(N281) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[14]), .Z(N280) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[13]), .Z(N279) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[12]), .Z(N278) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[11]), .Z(N277) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[10]), .Z(N276) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[9]), .Z(N275) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[8]), .Z(N274) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[7]), .Z(N273) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[5]), .Z(N271) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[4]), .Z(N270) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[3]), .Z(N269) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[1]), .Z(N267) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[0]), .Z(N266) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[62]), .Z(N362) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[60]), .Z(N360) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[59]), .Z(N359) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[58]), .Z(N358) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[57]), .Z(N357) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[56]), .Z(N356) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[55]), .Z(N355) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[54]), .Z(N354) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[53]), .Z(N353) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[52]), .Z(N352) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[51]), .Z(N351) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[50]), .Z(N350) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[49]), .Z(N349) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[48]), .Z(N348) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[47]), .Z(N347) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[46]), .Z(N346) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[45]), .Z(N345) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[44]), .Z(N344) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[43]), .Z(N343) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[42]), .Z(N342) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[41]), .Z(N341) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[40]), .Z(N340) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[39]), .Z(N339) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[38]), .Z(N338) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[37]), .Z(N337) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[19]), .Z(N285) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[89]), .Z(N423) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[88]), .Z(N422) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[87]), .Z(N421) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[85]), .Z(N419) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[84]), .Z(N418) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[83]), .Z(N417) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[81]), .Z(N415) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[80]), .Z(N414) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[79]), .Z(N413) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[78]), .Z(N412) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[77]), .Z(N411) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[76]), .Z(N410) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[75]), .Z(N409) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[74]), .Z(N408) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[73]), .Z(N407) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[72]), .Z(N406) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[71]), .Z(N405) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[70]), .Z(N404) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[69]), .Z(N403) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[68]), .Z(N402) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[67]), .Z(N401) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[66]), .Z(N400) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[65]), .Z(N399) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[64]), .Z(N398) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[36]), .Z(N336) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[34]), .Z(N334) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[33]), .Z(N333) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[32]), .Z(N332) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[95]), .Z(N429) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[94]), .Z(N428) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[93]), .Z(N427) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[92]), .Z(N426) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[35]), .Z(N335) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[91]), .Z(N425) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[90]), .Z(N424) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        CLK, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input CLK, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;
  wire   [127:0] buf_in_last_level_0__i_data_o_buf;
  wire   [127:0] buf_in_last_level_1__i_data_o_buf;
  wire   [127:0] buf_in_last_level_2__i_data_o_buf;
  wire   [127:0] buf_in_last_level_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[0]), .Z(
        buf_in_last_level_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[0]), .Z(
        buf_in_last_level_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[0]), .Z(
        buf_in_last_level_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[0]), .Z(
        buf_in_last_level_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[1]), .Z(
        buf_in_last_level_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[1]), .Z(
        buf_in_last_level_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[1]), .Z(
        buf_in_last_level_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[1]), .Z(
        buf_in_last_level_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[2]), .Z(
        buf_in_last_level_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[2]), .Z(
        buf_in_last_level_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[2]), .Z(
        buf_in_last_level_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[2]), .Z(
        buf_in_last_level_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[3]), .Z(
        buf_in_last_level_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[3]), .Z(
        buf_in_last_level_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[3]), .Z(
        buf_in_last_level_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[3]), .Z(
        buf_in_last_level_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[4]), .Z(
        buf_in_last_level_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[4]), .Z(
        buf_in_last_level_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[4]), .Z(
        buf_in_last_level_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[4]), .Z(
        buf_in_last_level_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[5]), .Z(
        buf_in_last_level_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[5]), .Z(
        buf_in_last_level_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[5]), .Z(
        buf_in_last_level_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[5]), .Z(
        buf_in_last_level_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[6]), .Z(
        buf_in_last_level_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[6]), .Z(
        buf_in_last_level_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[6]), .Z(
        buf_in_last_level_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[6]), .Z(
        buf_in_last_level_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[7]), .Z(
        buf_in_last_level_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[7]), .Z(
        buf_in_last_level_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[7]), .Z(
        buf_in_last_level_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[7]), .Z(
        buf_in_last_level_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[8]), .Z(
        buf_in_last_level_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[8]), .Z(
        buf_in_last_level_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[8]), .Z(
        buf_in_last_level_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[8]), .Z(
        buf_in_last_level_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[9]), .Z(
        buf_in_last_level_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[9]), .Z(
        buf_in_last_level_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[9]), .Z(
        buf_in_last_level_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[9]), .Z(
        buf_in_last_level_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[10]), .Z(
        buf_in_last_level_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[10]), .Z(
        buf_in_last_level_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[10]), .Z(
        buf_in_last_level_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[10]), .Z(
        buf_in_last_level_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[11]), .Z(
        buf_in_last_level_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[11]), .Z(
        buf_in_last_level_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[11]), .Z(
        buf_in_last_level_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[11]), .Z(
        buf_in_last_level_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[12]), .Z(
        buf_in_last_level_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[12]), .Z(
        buf_in_last_level_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[12]), .Z(
        buf_in_last_level_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[12]), .Z(
        buf_in_last_level_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[13]), .Z(
        buf_in_last_level_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[13]), .Z(
        buf_in_last_level_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[13]), .Z(
        buf_in_last_level_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[13]), .Z(
        buf_in_last_level_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[14]), .Z(
        buf_in_last_level_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[14]), .Z(
        buf_in_last_level_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[14]), .Z(
        buf_in_last_level_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[14]), .Z(
        buf_in_last_level_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[15]), .Z(
        buf_in_last_level_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[15]), .Z(
        buf_in_last_level_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[15]), .Z(
        buf_in_last_level_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[15]), .Z(
        buf_in_last_level_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[16]), .Z(
        buf_in_last_level_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[16]), .Z(
        buf_in_last_level_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[16]), .Z(
        buf_in_last_level_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[16]), .Z(
        buf_in_last_level_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[17]), .Z(
        buf_in_last_level_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[17]), .Z(
        buf_in_last_level_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[17]), .Z(
        buf_in_last_level_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[17]), .Z(
        buf_in_last_level_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[18]), .Z(
        buf_in_last_level_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[18]), .Z(
        buf_in_last_level_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[18]), .Z(
        buf_in_last_level_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[18]), .Z(
        buf_in_last_level_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[19]), .Z(
        buf_in_last_level_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[19]), .Z(
        buf_in_last_level_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[19]), .Z(
        buf_in_last_level_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[19]), .Z(
        buf_in_last_level_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[20]), .Z(
        buf_in_last_level_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[20]), .Z(
        buf_in_last_level_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[20]), .Z(
        buf_in_last_level_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[20]), .Z(
        buf_in_last_level_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[21]), .Z(
        buf_in_last_level_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[21]), .Z(
        buf_in_last_level_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[21]), .Z(
        buf_in_last_level_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[21]), .Z(
        buf_in_last_level_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[22]), .Z(
        buf_in_last_level_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[22]), .Z(
        buf_in_last_level_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[22]), .Z(
        buf_in_last_level_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[22]), .Z(
        buf_in_last_level_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[23]), .Z(
        buf_in_last_level_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[23]), .Z(
        buf_in_last_level_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[23]), .Z(
        buf_in_last_level_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[23]), .Z(
        buf_in_last_level_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[24]), .Z(
        buf_in_last_level_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[24]), .Z(
        buf_in_last_level_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[24]), .Z(
        buf_in_last_level_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[24]), .Z(
        buf_in_last_level_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[25]), .Z(
        buf_in_last_level_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[25]), .Z(
        buf_in_last_level_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[25]), .Z(
        buf_in_last_level_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[25]), .Z(
        buf_in_last_level_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[26]), .Z(
        buf_in_last_level_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[26]), .Z(
        buf_in_last_level_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[26]), .Z(
        buf_in_last_level_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[26]), .Z(
        buf_in_last_level_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[27]), .Z(
        buf_in_last_level_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[27]), .Z(
        buf_in_last_level_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[27]), .Z(
        buf_in_last_level_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[27]), .Z(
        buf_in_last_level_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[28]), .Z(
        buf_in_last_level_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[28]), .Z(
        buf_in_last_level_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[28]), .Z(
        buf_in_last_level_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[28]), .Z(
        buf_in_last_level_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[29]), .Z(
        buf_in_last_level_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[29]), .Z(
        buf_in_last_level_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[29]), .Z(
        buf_in_last_level_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[29]), .Z(
        buf_in_last_level_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[30]), .Z(
        buf_in_last_level_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[30]), .Z(
        buf_in_last_level_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[30]), .Z(
        buf_in_last_level_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[30]), .Z(
        buf_in_last_level_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[31]), .Z(
        buf_in_last_level_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[31]), .Z(
        buf_in_last_level_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[31]), .Z(
        buf_in_last_level_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[31]), .Z(
        buf_in_last_level_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[32]), .Z(
        buf_in_last_level_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[32]), .Z(
        buf_in_last_level_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[32]), .Z(
        buf_in_last_level_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[32]), .Z(
        buf_in_last_level_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[33]), .Z(
        buf_in_last_level_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[33]), .Z(
        buf_in_last_level_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[33]), .Z(
        buf_in_last_level_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[33]), .Z(
        buf_in_last_level_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[34]), .Z(
        buf_in_last_level_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[34]), .Z(
        buf_in_last_level_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[34]), .Z(
        buf_in_last_level_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[34]), .Z(
        buf_in_last_level_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[35]), .Z(
        buf_in_last_level_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[35]), .Z(
        buf_in_last_level_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[35]), .Z(
        buf_in_last_level_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[35]), .Z(
        buf_in_last_level_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[36]), .Z(
        buf_in_last_level_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[36]), .Z(
        buf_in_last_level_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[36]), .Z(
        buf_in_last_level_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[36]), .Z(
        buf_in_last_level_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[37]), .Z(
        buf_in_last_level_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[37]), .Z(
        buf_in_last_level_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[37]), .Z(
        buf_in_last_level_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[37]), .Z(
        buf_in_last_level_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[38]), .Z(
        buf_in_last_level_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[38]), .Z(
        buf_in_last_level_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[38]), .Z(
        buf_in_last_level_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[38]), .Z(
        buf_in_last_level_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[39]), .Z(
        buf_in_last_level_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[39]), .Z(
        buf_in_last_level_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[39]), .Z(
        buf_in_last_level_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[39]), .Z(
        buf_in_last_level_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[40]), .Z(
        buf_in_last_level_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[40]), .Z(
        buf_in_last_level_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[40]), .Z(
        buf_in_last_level_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[40]), .Z(
        buf_in_last_level_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[41]), .Z(
        buf_in_last_level_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[41]), .Z(
        buf_in_last_level_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[41]), .Z(
        buf_in_last_level_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[41]), .Z(
        buf_in_last_level_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[42]), .Z(
        buf_in_last_level_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[42]), .Z(
        buf_in_last_level_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[42]), .Z(
        buf_in_last_level_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[42]), .Z(
        buf_in_last_level_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[43]), .Z(
        buf_in_last_level_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[43]), .Z(
        buf_in_last_level_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[43]), .Z(
        buf_in_last_level_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[43]), .Z(
        buf_in_last_level_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[44]), .Z(
        buf_in_last_level_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[44]), .Z(
        buf_in_last_level_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[44]), .Z(
        buf_in_last_level_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[44]), .Z(
        buf_in_last_level_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[45]), .Z(
        buf_in_last_level_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[45]), .Z(
        buf_in_last_level_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[45]), .Z(
        buf_in_last_level_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[45]), .Z(
        buf_in_last_level_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[46]), .Z(
        buf_in_last_level_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[46]), .Z(
        buf_in_last_level_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[46]), .Z(
        buf_in_last_level_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[46]), .Z(
        buf_in_last_level_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[47]), .Z(
        buf_in_last_level_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[47]), .Z(
        buf_in_last_level_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[47]), .Z(
        buf_in_last_level_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[47]), .Z(
        buf_in_last_level_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[48]), .Z(
        buf_in_last_level_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[48]), .Z(
        buf_in_last_level_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[48]), .Z(
        buf_in_last_level_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[48]), .Z(
        buf_in_last_level_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[49]), .Z(
        buf_in_last_level_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[49]), .Z(
        buf_in_last_level_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[49]), .Z(
        buf_in_last_level_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[49]), .Z(
        buf_in_last_level_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[50]), .Z(
        buf_in_last_level_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[50]), .Z(
        buf_in_last_level_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[50]), .Z(
        buf_in_last_level_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[50]), .Z(
        buf_in_last_level_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[51]), .Z(
        buf_in_last_level_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[51]), .Z(
        buf_in_last_level_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[51]), .Z(
        buf_in_last_level_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[51]), .Z(
        buf_in_last_level_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[52]), .Z(
        buf_in_last_level_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[52]), .Z(
        buf_in_last_level_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[52]), .Z(
        buf_in_last_level_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[52]), .Z(
        buf_in_last_level_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[53]), .Z(
        buf_in_last_level_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[53]), .Z(
        buf_in_last_level_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[53]), .Z(
        buf_in_last_level_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[53]), .Z(
        buf_in_last_level_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[54]), .Z(
        buf_in_last_level_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[54]), .Z(
        buf_in_last_level_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[54]), .Z(
        buf_in_last_level_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[54]), .Z(
        buf_in_last_level_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[55]), .Z(
        buf_in_last_level_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[55]), .Z(
        buf_in_last_level_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[55]), .Z(
        buf_in_last_level_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[55]), .Z(
        buf_in_last_level_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[56]), .Z(
        buf_in_last_level_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[56]), .Z(
        buf_in_last_level_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[56]), .Z(
        buf_in_last_level_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[56]), .Z(
        buf_in_last_level_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[57]), .Z(
        buf_in_last_level_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[57]), .Z(
        buf_in_last_level_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[57]), .Z(
        buf_in_last_level_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[57]), .Z(
        buf_in_last_level_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[58]), .Z(
        buf_in_last_level_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[58]), .Z(
        buf_in_last_level_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[58]), .Z(
        buf_in_last_level_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[58]), .Z(
        buf_in_last_level_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[59]), .Z(
        buf_in_last_level_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[59]), .Z(
        buf_in_last_level_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[59]), .Z(
        buf_in_last_level_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[59]), .Z(
        buf_in_last_level_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[60]), .Z(
        buf_in_last_level_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[60]), .Z(
        buf_in_last_level_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[60]), .Z(
        buf_in_last_level_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[60]), .Z(
        buf_in_last_level_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[61]), .Z(
        buf_in_last_level_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[61]), .Z(
        buf_in_last_level_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[61]), .Z(
        buf_in_last_level_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[61]), .Z(
        buf_in_last_level_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[62]), .Z(
        buf_in_last_level_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[62]), .Z(
        buf_in_last_level_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[62]), .Z(
        buf_in_last_level_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[62]), .Z(
        buf_in_last_level_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[63]), .Z(
        buf_in_last_level_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[63]), .Z(
        buf_in_last_level_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[63]), .Z(
        buf_in_last_level_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[63]), .Z(
        buf_in_last_level_3__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[64]), .Z(
        buf_in_last_level_0__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[64]), .Z(
        buf_in_last_level_1__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[64]), .Z(
        buf_in_last_level_2__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[64]), .Z(
        buf_in_last_level_3__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[65]), .Z(
        buf_in_last_level_0__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[65]), .Z(
        buf_in_last_level_1__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[65]), .Z(
        buf_in_last_level_2__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[65]), .Z(
        buf_in_last_level_3__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[66]), .Z(
        buf_in_last_level_0__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[66]), .Z(
        buf_in_last_level_1__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[66]), .Z(
        buf_in_last_level_2__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[66]), .Z(
        buf_in_last_level_3__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[67]), .Z(
        buf_in_last_level_0__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[67]), .Z(
        buf_in_last_level_1__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[67]), .Z(
        buf_in_last_level_2__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[67]), .Z(
        buf_in_last_level_3__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[68]), .Z(
        buf_in_last_level_0__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[68]), .Z(
        buf_in_last_level_1__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[68]), .Z(
        buf_in_last_level_2__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[68]), .Z(
        buf_in_last_level_3__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[69]), .Z(
        buf_in_last_level_0__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[69]), .Z(
        buf_in_last_level_1__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[69]), .Z(
        buf_in_last_level_2__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[69]), .Z(
        buf_in_last_level_3__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[70]), .Z(
        buf_in_last_level_0__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[70]), .Z(
        buf_in_last_level_1__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[70]), .Z(
        buf_in_last_level_2__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[70]), .Z(
        buf_in_last_level_3__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[71]), .Z(
        buf_in_last_level_0__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[71]), .Z(
        buf_in_last_level_1__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[71]), .Z(
        buf_in_last_level_2__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[71]), .Z(
        buf_in_last_level_3__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[72]), .Z(
        buf_in_last_level_0__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[72]), .Z(
        buf_in_last_level_1__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[72]), .Z(
        buf_in_last_level_2__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[72]), .Z(
        buf_in_last_level_3__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[73]), .Z(
        buf_in_last_level_0__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[73]), .Z(
        buf_in_last_level_1__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[73]), .Z(
        buf_in_last_level_2__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[73]), .Z(
        buf_in_last_level_3__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[74]), .Z(
        buf_in_last_level_0__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[74]), .Z(
        buf_in_last_level_1__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[74]), .Z(
        buf_in_last_level_2__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[74]), .Z(
        buf_in_last_level_3__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[75]), .Z(
        buf_in_last_level_0__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[75]), .Z(
        buf_in_last_level_1__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[75]), .Z(
        buf_in_last_level_2__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[75]), .Z(
        buf_in_last_level_3__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[76]), .Z(
        buf_in_last_level_0__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[76]), .Z(
        buf_in_last_level_1__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[76]), .Z(
        buf_in_last_level_2__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[76]), .Z(
        buf_in_last_level_3__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[77]), .Z(
        buf_in_last_level_0__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[77]), .Z(
        buf_in_last_level_1__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[77]), .Z(
        buf_in_last_level_2__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[77]), .Z(
        buf_in_last_level_3__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[78]), .Z(
        buf_in_last_level_0__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[78]), .Z(
        buf_in_last_level_1__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[78]), .Z(
        buf_in_last_level_2__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[78]), .Z(
        buf_in_last_level_3__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[79]), .Z(
        buf_in_last_level_0__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[79]), .Z(
        buf_in_last_level_1__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[79]), .Z(
        buf_in_last_level_2__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[79]), .Z(
        buf_in_last_level_3__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[80]), .Z(
        buf_in_last_level_0__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[80]), .Z(
        buf_in_last_level_1__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[80]), .Z(
        buf_in_last_level_2__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[80]), .Z(
        buf_in_last_level_3__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[81]), .Z(
        buf_in_last_level_0__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[81]), .Z(
        buf_in_last_level_1__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[81]), .Z(
        buf_in_last_level_2__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[81]), .Z(
        buf_in_last_level_3__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[82]), .Z(
        buf_in_last_level_0__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[82]), .Z(
        buf_in_last_level_1__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[82]), .Z(
        buf_in_last_level_2__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[82]), .Z(
        buf_in_last_level_3__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[83]), .Z(
        buf_in_last_level_0__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[83]), .Z(
        buf_in_last_level_1__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[83]), .Z(
        buf_in_last_level_2__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[83]), .Z(
        buf_in_last_level_3__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[84]), .Z(
        buf_in_last_level_0__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[84]), .Z(
        buf_in_last_level_1__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[84]), .Z(
        buf_in_last_level_2__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[84]), .Z(
        buf_in_last_level_3__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[85]), .Z(
        buf_in_last_level_0__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[85]), .Z(
        buf_in_last_level_1__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[85]), .Z(
        buf_in_last_level_2__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[85]), .Z(
        buf_in_last_level_3__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[86]), .Z(
        buf_in_last_level_0__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[86]), .Z(
        buf_in_last_level_1__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[86]), .Z(
        buf_in_last_level_2__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[86]), .Z(
        buf_in_last_level_3__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[87]), .Z(
        buf_in_last_level_0__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[87]), .Z(
        buf_in_last_level_1__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[87]), .Z(
        buf_in_last_level_2__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[87]), .Z(
        buf_in_last_level_3__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[88]), .Z(
        buf_in_last_level_0__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[88]), .Z(
        buf_in_last_level_1__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[88]), .Z(
        buf_in_last_level_2__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[88]), .Z(
        buf_in_last_level_3__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[89]), .Z(
        buf_in_last_level_0__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[89]), .Z(
        buf_in_last_level_1__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[89]), .Z(
        buf_in_last_level_2__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[89]), .Z(
        buf_in_last_level_3__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[90]), .Z(
        buf_in_last_level_0__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[90]), .Z(
        buf_in_last_level_1__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[90]), .Z(
        buf_in_last_level_2__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[90]), .Z(
        buf_in_last_level_3__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[91]), .Z(
        buf_in_last_level_0__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[91]), .Z(
        buf_in_last_level_1__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[91]), .Z(
        buf_in_last_level_2__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[91]), .Z(
        buf_in_last_level_3__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[92]), .Z(
        buf_in_last_level_0__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[92]), .Z(
        buf_in_last_level_1__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[92]), .Z(
        buf_in_last_level_2__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[92]), .Z(
        buf_in_last_level_3__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[93]), .Z(
        buf_in_last_level_0__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[93]), .Z(
        buf_in_last_level_1__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[93]), .Z(
        buf_in_last_level_2__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[93]), .Z(
        buf_in_last_level_3__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[94]), .Z(
        buf_in_last_level_0__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[94]), .Z(
        buf_in_last_level_1__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[94]), .Z(
        buf_in_last_level_2__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[94]), .Z(
        buf_in_last_level_3__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[95]), .Z(
        buf_in_last_level_0__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[95]), .Z(
        buf_in_last_level_1__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[95]), .Z(
        buf_in_last_level_2__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[95]), .Z(
        buf_in_last_level_3__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[96]), .Z(
        buf_in_last_level_0__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[96]), .Z(
        buf_in_last_level_1__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[96]), .Z(
        buf_in_last_level_2__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[96]), .Z(
        buf_in_last_level_3__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[97]), .Z(
        buf_in_last_level_0__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[97]), .Z(
        buf_in_last_level_1__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[97]), .Z(
        buf_in_last_level_2__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[97]), .Z(
        buf_in_last_level_3__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[98]), .Z(
        buf_in_last_level_0__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[98]), .Z(
        buf_in_last_level_1__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[98]), .Z(
        buf_in_last_level_2__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[98]), .Z(
        buf_in_last_level_3__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[99]), .Z(
        buf_in_last_level_0__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[99]), .Z(
        buf_in_last_level_1__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[99]), .Z(
        buf_in_last_level_2__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[99]), .Z(
        buf_in_last_level_3__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[100]), .Z(
        buf_in_last_level_0__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[100]), .Z(
        buf_in_last_level_1__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[100]), .Z(
        buf_in_last_level_2__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[100]), .Z(
        buf_in_last_level_3__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[101]), .Z(
        buf_in_last_level_0__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[101]), .Z(
        buf_in_last_level_1__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[101]), .Z(
        buf_in_last_level_2__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[101]), .Z(
        buf_in_last_level_3__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[102]), .Z(
        buf_in_last_level_0__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[102]), .Z(
        buf_in_last_level_1__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[102]), .Z(
        buf_in_last_level_2__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[102]), .Z(
        buf_in_last_level_3__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[103]), .Z(
        buf_in_last_level_0__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[103]), .Z(
        buf_in_last_level_1__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[103]), .Z(
        buf_in_last_level_2__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[103]), .Z(
        buf_in_last_level_3__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[104]), .Z(
        buf_in_last_level_0__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[104]), .Z(
        buf_in_last_level_1__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[104]), .Z(
        buf_in_last_level_2__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[104]), .Z(
        buf_in_last_level_3__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[105]), .Z(
        buf_in_last_level_0__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[105]), .Z(
        buf_in_last_level_1__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[105]), .Z(
        buf_in_last_level_2__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[105]), .Z(
        buf_in_last_level_3__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[106]), .Z(
        buf_in_last_level_0__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[106]), .Z(
        buf_in_last_level_1__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[106]), .Z(
        buf_in_last_level_2__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[106]), .Z(
        buf_in_last_level_3__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[107]), .Z(
        buf_in_last_level_0__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[107]), .Z(
        buf_in_last_level_1__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[107]), .Z(
        buf_in_last_level_2__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[107]), .Z(
        buf_in_last_level_3__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[108]), .Z(
        buf_in_last_level_0__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[108]), .Z(
        buf_in_last_level_1__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[108]), .Z(
        buf_in_last_level_2__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[108]), .Z(
        buf_in_last_level_3__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[109]), .Z(
        buf_in_last_level_0__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[109]), .Z(
        buf_in_last_level_1__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[109]), .Z(
        buf_in_last_level_2__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[109]), .Z(
        buf_in_last_level_3__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[110]), .Z(
        buf_in_last_level_0__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[110]), .Z(
        buf_in_last_level_1__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[110]), .Z(
        buf_in_last_level_2__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[110]), .Z(
        buf_in_last_level_3__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[111]), .Z(
        buf_in_last_level_0__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[111]), .Z(
        buf_in_last_level_1__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[111]), .Z(
        buf_in_last_level_2__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[111]), .Z(
        buf_in_last_level_3__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[112]), .Z(
        buf_in_last_level_0__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[112]), .Z(
        buf_in_last_level_1__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[112]), .Z(
        buf_in_last_level_2__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[112]), .Z(
        buf_in_last_level_3__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[113]), .Z(
        buf_in_last_level_0__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[113]), .Z(
        buf_in_last_level_1__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[113]), .Z(
        buf_in_last_level_2__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[113]), .Z(
        buf_in_last_level_3__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[114]), .Z(
        buf_in_last_level_0__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[114]), .Z(
        buf_in_last_level_1__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[114]), .Z(
        buf_in_last_level_2__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[114]), .Z(
        buf_in_last_level_3__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[115]), .Z(
        buf_in_last_level_0__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[115]), .Z(
        buf_in_last_level_1__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[115]), .Z(
        buf_in_last_level_2__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[115]), .Z(
        buf_in_last_level_3__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[116]), .Z(
        buf_in_last_level_0__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[116]), .Z(
        buf_in_last_level_1__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[116]), .Z(
        buf_in_last_level_2__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[116]), .Z(
        buf_in_last_level_3__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[117]), .Z(
        buf_in_last_level_0__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[117]), .Z(
        buf_in_last_level_1__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[117]), .Z(
        buf_in_last_level_2__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[117]), .Z(
        buf_in_last_level_3__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[118]), .Z(
        buf_in_last_level_0__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[118]), .Z(
        buf_in_last_level_1__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[118]), .Z(
        buf_in_last_level_2__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[118]), .Z(
        buf_in_last_level_3__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[119]), .Z(
        buf_in_last_level_0__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[119]), .Z(
        buf_in_last_level_1__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[119]), .Z(
        buf_in_last_level_2__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[119]), .Z(
        buf_in_last_level_3__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[120]), .Z(
        buf_in_last_level_0__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[120]), .Z(
        buf_in_last_level_1__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[120]), .Z(
        buf_in_last_level_2__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[120]), .Z(
        buf_in_last_level_3__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[121]), .Z(
        buf_in_last_level_0__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[121]), .Z(
        buf_in_last_level_1__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[121]), .Z(
        buf_in_last_level_2__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[121]), .Z(
        buf_in_last_level_3__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[122]), .Z(
        buf_in_last_level_0__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[122]), .Z(
        buf_in_last_level_1__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[122]), .Z(
        buf_in_last_level_2__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[122]), .Z(
        buf_in_last_level_3__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[123]), .Z(
        buf_in_last_level_0__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[123]), .Z(
        buf_in_last_level_1__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[123]), .Z(
        buf_in_last_level_2__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[123]), .Z(
        buf_in_last_level_3__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[124]), .Z(
        buf_in_last_level_0__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[124]), .Z(
        buf_in_last_level_1__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[124]), .Z(
        buf_in_last_level_2__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[124]), .Z(
        buf_in_last_level_3__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[125]), .Z(
        buf_in_last_level_0__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[125]), .Z(
        buf_in_last_level_1__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[125]), .Z(
        buf_in_last_level_2__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[125]), .Z(
        buf_in_last_level_3__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[126]), .Z(
        buf_in_last_level_0__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[126]), .Z(
        buf_in_last_level_1__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[126]), .Z(
        buf_in_last_level_2__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[126]), .Z(
        buf_in_last_level_3__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[127]), .Z(
        buf_in_last_level_0__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[127]), .Z(
        buf_in_last_level_1__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[127]), .Z(
        buf_in_last_level_2__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[127]), .Z(
        buf_in_last_level_3__i_data_o_buf[127]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(CLK), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(CLK), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(CLK), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(CLK), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(CLK), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(CLK), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(CLK), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(CLK), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[101]), .Z(N469) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[102]), .Z(N470) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[105]), .Z(N473) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[107]), .Z(N475) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[109]), .Z(N477) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[110]), .Z(N478) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[111]), .Z(N479) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[112]), .Z(N480) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[115]), .Z(N483) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[82]), .Z(N416) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[86]), .Z(N420) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[61]), .Z(N361) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[63]), .Z(N363) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[31]), .Z(N297) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[30]), .Z(N296) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[29]), .Z(N295) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[28]), .Z(N294) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[27]), .Z(N293) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[26]), .Z(N292) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[25]), .Z(N291) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[24]), .Z(N290) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[23]), .Z(N289) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[22]), .Z(N288) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[21]), .Z(N287) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[20]), .Z(N286) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[37]), .Z(N337) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[38]), .Z(N338) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[39]), .Z(N339) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[40]), .Z(N340) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[41]), .Z(N341) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[42]), .Z(N342) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[43]), .Z(N343) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[44]), .Z(N344) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[45]), .Z(N345) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[46]), .Z(N346) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[47]), .Z(N347) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[48]), .Z(N348) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[49]), .Z(N349) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[50]), .Z(N350) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[51]), .Z(N351) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[52]), .Z(N352) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[53]), .Z(N353) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[54]), .Z(N354) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[55]), .Z(N355) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[56]), .Z(N356) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[57]), .Z(N357) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[58]), .Z(N358) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[59]), .Z(N359) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[60]), .Z(N360) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[62]), .Z(N362) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[0]), .Z(N266) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[1]), .Z(N267) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[3]), .Z(N269) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[4]), .Z(N270) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[5]), .Z(N271) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[7]), .Z(N273) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[8]), .Z(N274) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[9]), .Z(N275) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[10]), .Z(N276) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[11]), .Z(N277) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[12]), .Z(N278) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[13]), .Z(N279) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[14]), .Z(N280) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[15]), .Z(N281) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[16]), .Z(N282) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[17]), .Z(N283) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[18]), .Z(N284) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[19]), .Z(N285) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[36]), .Z(N336) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[35]), .Z(N335) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[34]), .Z(N334) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[65]), .Z(N399) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[66]), .Z(N400) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[67]), .Z(N401) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[64]), .Z(N398) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[69]), .Z(N403) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[70]), .Z(N404) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[71]), .Z(N405) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[72]), .Z(N406) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[73]), .Z(N407) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[74]), .Z(N408) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[75]), .Z(N409) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[76]), .Z(N410) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[77]), .Z(N411) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[78]), .Z(N412) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[79]), .Z(N413) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[80]), .Z(N414) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[81]), .Z(N415) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[83]), .Z(N417) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[84]), .Z(N418) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[85]), .Z(N419) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[89]), .Z(N423) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[68]), .Z(N402) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[32]), .Z(N332) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[33]), .Z(N333) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[91]), .Z(N425) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[92]), .Z(N426) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[95]), .Z(N429) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[93]), .Z(N427) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[90]), .Z(N424) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[88]), .Z(N422) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[87]), .Z(N421) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[94]), .Z(N428) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        CLK, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input CLK, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;
  wire   [127:0] buf_in_last_level_0__i_data_o_buf;
  wire   [127:0] buf_in_last_level_1__i_data_o_buf;
  wire   [127:0] buf_in_last_level_2__i_data_o_buf;
  wire   [127:0] buf_in_last_level_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[0]), .Z(
        buf_in_last_level_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[0]), .Z(
        buf_in_last_level_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[0]), .Z(
        buf_in_last_level_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[0]), .Z(
        buf_in_last_level_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[1]), .Z(
        buf_in_last_level_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[1]), .Z(
        buf_in_last_level_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[1]), .Z(
        buf_in_last_level_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[1]), .Z(
        buf_in_last_level_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[2]), .Z(
        buf_in_last_level_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[2]), .Z(
        buf_in_last_level_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[2]), .Z(
        buf_in_last_level_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[2]), .Z(
        buf_in_last_level_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[3]), .Z(
        buf_in_last_level_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[3]), .Z(
        buf_in_last_level_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[3]), .Z(
        buf_in_last_level_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[3]), .Z(
        buf_in_last_level_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[4]), .Z(
        buf_in_last_level_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[4]), .Z(
        buf_in_last_level_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[4]), .Z(
        buf_in_last_level_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[4]), .Z(
        buf_in_last_level_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[5]), .Z(
        buf_in_last_level_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[5]), .Z(
        buf_in_last_level_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[5]), .Z(
        buf_in_last_level_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[5]), .Z(
        buf_in_last_level_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[6]), .Z(
        buf_in_last_level_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[6]), .Z(
        buf_in_last_level_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[6]), .Z(
        buf_in_last_level_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[6]), .Z(
        buf_in_last_level_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[7]), .Z(
        buf_in_last_level_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[7]), .Z(
        buf_in_last_level_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[7]), .Z(
        buf_in_last_level_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[7]), .Z(
        buf_in_last_level_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[8]), .Z(
        buf_in_last_level_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[8]), .Z(
        buf_in_last_level_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[8]), .Z(
        buf_in_last_level_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[8]), .Z(
        buf_in_last_level_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[9]), .Z(
        buf_in_last_level_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[9]), .Z(
        buf_in_last_level_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[9]), .Z(
        buf_in_last_level_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[9]), .Z(
        buf_in_last_level_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[10]), .Z(
        buf_in_last_level_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[10]), .Z(
        buf_in_last_level_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[10]), .Z(
        buf_in_last_level_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[10]), .Z(
        buf_in_last_level_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[11]), .Z(
        buf_in_last_level_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[11]), .Z(
        buf_in_last_level_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[11]), .Z(
        buf_in_last_level_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[11]), .Z(
        buf_in_last_level_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[12]), .Z(
        buf_in_last_level_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[12]), .Z(
        buf_in_last_level_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[12]), .Z(
        buf_in_last_level_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[12]), .Z(
        buf_in_last_level_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[13]), .Z(
        buf_in_last_level_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[13]), .Z(
        buf_in_last_level_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[13]), .Z(
        buf_in_last_level_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[13]), .Z(
        buf_in_last_level_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[14]), .Z(
        buf_in_last_level_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[14]), .Z(
        buf_in_last_level_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[14]), .Z(
        buf_in_last_level_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[14]), .Z(
        buf_in_last_level_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[15]), .Z(
        buf_in_last_level_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[15]), .Z(
        buf_in_last_level_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[15]), .Z(
        buf_in_last_level_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[15]), .Z(
        buf_in_last_level_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[16]), .Z(
        buf_in_last_level_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[16]), .Z(
        buf_in_last_level_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[16]), .Z(
        buf_in_last_level_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[16]), .Z(
        buf_in_last_level_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[17]), .Z(
        buf_in_last_level_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[17]), .Z(
        buf_in_last_level_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[17]), .Z(
        buf_in_last_level_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[17]), .Z(
        buf_in_last_level_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[18]), .Z(
        buf_in_last_level_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[18]), .Z(
        buf_in_last_level_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[18]), .Z(
        buf_in_last_level_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[18]), .Z(
        buf_in_last_level_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[19]), .Z(
        buf_in_last_level_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[19]), .Z(
        buf_in_last_level_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[19]), .Z(
        buf_in_last_level_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[19]), .Z(
        buf_in_last_level_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[20]), .Z(
        buf_in_last_level_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[20]), .Z(
        buf_in_last_level_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[20]), .Z(
        buf_in_last_level_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[20]), .Z(
        buf_in_last_level_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[21]), .Z(
        buf_in_last_level_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[21]), .Z(
        buf_in_last_level_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[21]), .Z(
        buf_in_last_level_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[21]), .Z(
        buf_in_last_level_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[22]), .Z(
        buf_in_last_level_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[22]), .Z(
        buf_in_last_level_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[22]), .Z(
        buf_in_last_level_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[22]), .Z(
        buf_in_last_level_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[23]), .Z(
        buf_in_last_level_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[23]), .Z(
        buf_in_last_level_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[23]), .Z(
        buf_in_last_level_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[23]), .Z(
        buf_in_last_level_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[24]), .Z(
        buf_in_last_level_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[24]), .Z(
        buf_in_last_level_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[24]), .Z(
        buf_in_last_level_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[24]), .Z(
        buf_in_last_level_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[25]), .Z(
        buf_in_last_level_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[25]), .Z(
        buf_in_last_level_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[25]), .Z(
        buf_in_last_level_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[25]), .Z(
        buf_in_last_level_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[26]), .Z(
        buf_in_last_level_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[26]), .Z(
        buf_in_last_level_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[26]), .Z(
        buf_in_last_level_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[26]), .Z(
        buf_in_last_level_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[27]), .Z(
        buf_in_last_level_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[27]), .Z(
        buf_in_last_level_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[27]), .Z(
        buf_in_last_level_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[27]), .Z(
        buf_in_last_level_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[28]), .Z(
        buf_in_last_level_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[28]), .Z(
        buf_in_last_level_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[28]), .Z(
        buf_in_last_level_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[28]), .Z(
        buf_in_last_level_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[29]), .Z(
        buf_in_last_level_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[29]), .Z(
        buf_in_last_level_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[29]), .Z(
        buf_in_last_level_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[29]), .Z(
        buf_in_last_level_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[30]), .Z(
        buf_in_last_level_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[30]), .Z(
        buf_in_last_level_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[30]), .Z(
        buf_in_last_level_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[30]), .Z(
        buf_in_last_level_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[31]), .Z(
        buf_in_last_level_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[31]), .Z(
        buf_in_last_level_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[31]), .Z(
        buf_in_last_level_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[31]), .Z(
        buf_in_last_level_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[32]), .Z(
        buf_in_last_level_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[32]), .Z(
        buf_in_last_level_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[32]), .Z(
        buf_in_last_level_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[32]), .Z(
        buf_in_last_level_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[33]), .Z(
        buf_in_last_level_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[33]), .Z(
        buf_in_last_level_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[33]), .Z(
        buf_in_last_level_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[33]), .Z(
        buf_in_last_level_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[34]), .Z(
        buf_in_last_level_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[34]), .Z(
        buf_in_last_level_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[34]), .Z(
        buf_in_last_level_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[34]), .Z(
        buf_in_last_level_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[35]), .Z(
        buf_in_last_level_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[35]), .Z(
        buf_in_last_level_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[35]), .Z(
        buf_in_last_level_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[35]), .Z(
        buf_in_last_level_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[36]), .Z(
        buf_in_last_level_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[36]), .Z(
        buf_in_last_level_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[36]), .Z(
        buf_in_last_level_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[36]), .Z(
        buf_in_last_level_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[37]), .Z(
        buf_in_last_level_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[37]), .Z(
        buf_in_last_level_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[37]), .Z(
        buf_in_last_level_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[37]), .Z(
        buf_in_last_level_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[38]), .Z(
        buf_in_last_level_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[38]), .Z(
        buf_in_last_level_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[38]), .Z(
        buf_in_last_level_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[38]), .Z(
        buf_in_last_level_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[39]), .Z(
        buf_in_last_level_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[39]), .Z(
        buf_in_last_level_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[39]), .Z(
        buf_in_last_level_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[39]), .Z(
        buf_in_last_level_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[40]), .Z(
        buf_in_last_level_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[40]), .Z(
        buf_in_last_level_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[40]), .Z(
        buf_in_last_level_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[40]), .Z(
        buf_in_last_level_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[41]), .Z(
        buf_in_last_level_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[41]), .Z(
        buf_in_last_level_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[41]), .Z(
        buf_in_last_level_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[41]), .Z(
        buf_in_last_level_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[42]), .Z(
        buf_in_last_level_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[42]), .Z(
        buf_in_last_level_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[42]), .Z(
        buf_in_last_level_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[42]), .Z(
        buf_in_last_level_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[43]), .Z(
        buf_in_last_level_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[43]), .Z(
        buf_in_last_level_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[43]), .Z(
        buf_in_last_level_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[43]), .Z(
        buf_in_last_level_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[44]), .Z(
        buf_in_last_level_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[44]), .Z(
        buf_in_last_level_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[44]), .Z(
        buf_in_last_level_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[44]), .Z(
        buf_in_last_level_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[45]), .Z(
        buf_in_last_level_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[45]), .Z(
        buf_in_last_level_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[45]), .Z(
        buf_in_last_level_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[45]), .Z(
        buf_in_last_level_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[46]), .Z(
        buf_in_last_level_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[46]), .Z(
        buf_in_last_level_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[46]), .Z(
        buf_in_last_level_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[46]), .Z(
        buf_in_last_level_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[47]), .Z(
        buf_in_last_level_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[47]), .Z(
        buf_in_last_level_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[47]), .Z(
        buf_in_last_level_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[47]), .Z(
        buf_in_last_level_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[48]), .Z(
        buf_in_last_level_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[48]), .Z(
        buf_in_last_level_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[48]), .Z(
        buf_in_last_level_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[48]), .Z(
        buf_in_last_level_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[49]), .Z(
        buf_in_last_level_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[49]), .Z(
        buf_in_last_level_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[49]), .Z(
        buf_in_last_level_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[49]), .Z(
        buf_in_last_level_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[50]), .Z(
        buf_in_last_level_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[50]), .Z(
        buf_in_last_level_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[50]), .Z(
        buf_in_last_level_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[50]), .Z(
        buf_in_last_level_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[51]), .Z(
        buf_in_last_level_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[51]), .Z(
        buf_in_last_level_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[51]), .Z(
        buf_in_last_level_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[51]), .Z(
        buf_in_last_level_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[52]), .Z(
        buf_in_last_level_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[52]), .Z(
        buf_in_last_level_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[52]), .Z(
        buf_in_last_level_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[52]), .Z(
        buf_in_last_level_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[53]), .Z(
        buf_in_last_level_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[53]), .Z(
        buf_in_last_level_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[53]), .Z(
        buf_in_last_level_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[53]), .Z(
        buf_in_last_level_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[54]), .Z(
        buf_in_last_level_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[54]), .Z(
        buf_in_last_level_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[54]), .Z(
        buf_in_last_level_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[54]), .Z(
        buf_in_last_level_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[55]), .Z(
        buf_in_last_level_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[55]), .Z(
        buf_in_last_level_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[55]), .Z(
        buf_in_last_level_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[55]), .Z(
        buf_in_last_level_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[56]), .Z(
        buf_in_last_level_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[56]), .Z(
        buf_in_last_level_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[56]), .Z(
        buf_in_last_level_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[56]), .Z(
        buf_in_last_level_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[57]), .Z(
        buf_in_last_level_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[57]), .Z(
        buf_in_last_level_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[57]), .Z(
        buf_in_last_level_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[57]), .Z(
        buf_in_last_level_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[58]), .Z(
        buf_in_last_level_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[58]), .Z(
        buf_in_last_level_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[58]), .Z(
        buf_in_last_level_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[58]), .Z(
        buf_in_last_level_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[59]), .Z(
        buf_in_last_level_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[59]), .Z(
        buf_in_last_level_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[59]), .Z(
        buf_in_last_level_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[59]), .Z(
        buf_in_last_level_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[60]), .Z(
        buf_in_last_level_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[60]), .Z(
        buf_in_last_level_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[60]), .Z(
        buf_in_last_level_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[60]), .Z(
        buf_in_last_level_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[61]), .Z(
        buf_in_last_level_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[61]), .Z(
        buf_in_last_level_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[61]), .Z(
        buf_in_last_level_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[61]), .Z(
        buf_in_last_level_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[62]), .Z(
        buf_in_last_level_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[62]), .Z(
        buf_in_last_level_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[62]), .Z(
        buf_in_last_level_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[62]), .Z(
        buf_in_last_level_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[63]), .Z(
        buf_in_last_level_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[63]), .Z(
        buf_in_last_level_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[63]), .Z(
        buf_in_last_level_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[63]), .Z(
        buf_in_last_level_3__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[64]), .Z(
        buf_in_last_level_0__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[64]), .Z(
        buf_in_last_level_1__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[64]), .Z(
        buf_in_last_level_2__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[64]), .Z(
        buf_in_last_level_3__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[65]), .Z(
        buf_in_last_level_0__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[65]), .Z(
        buf_in_last_level_1__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[65]), .Z(
        buf_in_last_level_2__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[65]), .Z(
        buf_in_last_level_3__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[66]), .Z(
        buf_in_last_level_0__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[66]), .Z(
        buf_in_last_level_1__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[66]), .Z(
        buf_in_last_level_2__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[66]), .Z(
        buf_in_last_level_3__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[67]), .Z(
        buf_in_last_level_0__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[67]), .Z(
        buf_in_last_level_1__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[67]), .Z(
        buf_in_last_level_2__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[67]), .Z(
        buf_in_last_level_3__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[68]), .Z(
        buf_in_last_level_0__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[68]), .Z(
        buf_in_last_level_1__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[68]), .Z(
        buf_in_last_level_2__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[68]), .Z(
        buf_in_last_level_3__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[69]), .Z(
        buf_in_last_level_0__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[69]), .Z(
        buf_in_last_level_1__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[69]), .Z(
        buf_in_last_level_2__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[69]), .Z(
        buf_in_last_level_3__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[70]), .Z(
        buf_in_last_level_0__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[70]), .Z(
        buf_in_last_level_1__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[70]), .Z(
        buf_in_last_level_2__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[70]), .Z(
        buf_in_last_level_3__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[71]), .Z(
        buf_in_last_level_0__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[71]), .Z(
        buf_in_last_level_1__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[71]), .Z(
        buf_in_last_level_2__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[71]), .Z(
        buf_in_last_level_3__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[72]), .Z(
        buf_in_last_level_0__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[72]), .Z(
        buf_in_last_level_1__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[72]), .Z(
        buf_in_last_level_2__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[72]), .Z(
        buf_in_last_level_3__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[73]), .Z(
        buf_in_last_level_0__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[73]), .Z(
        buf_in_last_level_1__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[73]), .Z(
        buf_in_last_level_2__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[73]), .Z(
        buf_in_last_level_3__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[74]), .Z(
        buf_in_last_level_0__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[74]), .Z(
        buf_in_last_level_1__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[74]), .Z(
        buf_in_last_level_2__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[74]), .Z(
        buf_in_last_level_3__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[75]), .Z(
        buf_in_last_level_0__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[75]), .Z(
        buf_in_last_level_1__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[75]), .Z(
        buf_in_last_level_2__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[75]), .Z(
        buf_in_last_level_3__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[76]), .Z(
        buf_in_last_level_0__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[76]), .Z(
        buf_in_last_level_1__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[76]), .Z(
        buf_in_last_level_2__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[76]), .Z(
        buf_in_last_level_3__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[77]), .Z(
        buf_in_last_level_0__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[77]), .Z(
        buf_in_last_level_1__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[77]), .Z(
        buf_in_last_level_2__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[77]), .Z(
        buf_in_last_level_3__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[78]), .Z(
        buf_in_last_level_0__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[78]), .Z(
        buf_in_last_level_1__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[78]), .Z(
        buf_in_last_level_2__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[78]), .Z(
        buf_in_last_level_3__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[79]), .Z(
        buf_in_last_level_0__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[79]), .Z(
        buf_in_last_level_1__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[79]), .Z(
        buf_in_last_level_2__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[79]), .Z(
        buf_in_last_level_3__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[80]), .Z(
        buf_in_last_level_0__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[80]), .Z(
        buf_in_last_level_1__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[80]), .Z(
        buf_in_last_level_2__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[80]), .Z(
        buf_in_last_level_3__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[81]), .Z(
        buf_in_last_level_0__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[81]), .Z(
        buf_in_last_level_1__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[81]), .Z(
        buf_in_last_level_2__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[81]), .Z(
        buf_in_last_level_3__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[82]), .Z(
        buf_in_last_level_0__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[82]), .Z(
        buf_in_last_level_1__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[82]), .Z(
        buf_in_last_level_2__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[82]), .Z(
        buf_in_last_level_3__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[83]), .Z(
        buf_in_last_level_0__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[83]), .Z(
        buf_in_last_level_1__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[83]), .Z(
        buf_in_last_level_2__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[83]), .Z(
        buf_in_last_level_3__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[84]), .Z(
        buf_in_last_level_0__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[84]), .Z(
        buf_in_last_level_1__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[84]), .Z(
        buf_in_last_level_2__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[84]), .Z(
        buf_in_last_level_3__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[85]), .Z(
        buf_in_last_level_0__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[85]), .Z(
        buf_in_last_level_1__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[85]), .Z(
        buf_in_last_level_2__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[85]), .Z(
        buf_in_last_level_3__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[86]), .Z(
        buf_in_last_level_0__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[86]), .Z(
        buf_in_last_level_1__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[86]), .Z(
        buf_in_last_level_2__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[86]), .Z(
        buf_in_last_level_3__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[87]), .Z(
        buf_in_last_level_0__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[87]), .Z(
        buf_in_last_level_1__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[87]), .Z(
        buf_in_last_level_2__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[87]), .Z(
        buf_in_last_level_3__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[88]), .Z(
        buf_in_last_level_0__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[88]), .Z(
        buf_in_last_level_1__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[88]), .Z(
        buf_in_last_level_2__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[88]), .Z(
        buf_in_last_level_3__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[89]), .Z(
        buf_in_last_level_0__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[89]), .Z(
        buf_in_last_level_1__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[89]), .Z(
        buf_in_last_level_2__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[89]), .Z(
        buf_in_last_level_3__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[90]), .Z(
        buf_in_last_level_0__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[90]), .Z(
        buf_in_last_level_1__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[90]), .Z(
        buf_in_last_level_2__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[90]), .Z(
        buf_in_last_level_3__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[91]), .Z(
        buf_in_last_level_0__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[91]), .Z(
        buf_in_last_level_1__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[91]), .Z(
        buf_in_last_level_2__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[91]), .Z(
        buf_in_last_level_3__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[92]), .Z(
        buf_in_last_level_0__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[92]), .Z(
        buf_in_last_level_1__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[92]), .Z(
        buf_in_last_level_2__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[92]), .Z(
        buf_in_last_level_3__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[93]), .Z(
        buf_in_last_level_0__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[93]), .Z(
        buf_in_last_level_1__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[93]), .Z(
        buf_in_last_level_2__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[93]), .Z(
        buf_in_last_level_3__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[94]), .Z(
        buf_in_last_level_0__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[94]), .Z(
        buf_in_last_level_1__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[94]), .Z(
        buf_in_last_level_2__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[94]), .Z(
        buf_in_last_level_3__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[95]), .Z(
        buf_in_last_level_0__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[95]), .Z(
        buf_in_last_level_1__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[95]), .Z(
        buf_in_last_level_2__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[95]), .Z(
        buf_in_last_level_3__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[96]), .Z(
        buf_in_last_level_0__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[96]), .Z(
        buf_in_last_level_1__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[96]), .Z(
        buf_in_last_level_2__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[96]), .Z(
        buf_in_last_level_3__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[97]), .Z(
        buf_in_last_level_0__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[97]), .Z(
        buf_in_last_level_1__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[97]), .Z(
        buf_in_last_level_2__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[97]), .Z(
        buf_in_last_level_3__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[98]), .Z(
        buf_in_last_level_0__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[98]), .Z(
        buf_in_last_level_1__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[98]), .Z(
        buf_in_last_level_2__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[98]), .Z(
        buf_in_last_level_3__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[99]), .Z(
        buf_in_last_level_0__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[99]), .Z(
        buf_in_last_level_1__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[99]), .Z(
        buf_in_last_level_2__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[99]), .Z(
        buf_in_last_level_3__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[100]), .Z(
        buf_in_last_level_0__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[100]), .Z(
        buf_in_last_level_1__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[100]), .Z(
        buf_in_last_level_2__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[100]), .Z(
        buf_in_last_level_3__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[101]), .Z(
        buf_in_last_level_0__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[101]), .Z(
        buf_in_last_level_1__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[101]), .Z(
        buf_in_last_level_2__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[101]), .Z(
        buf_in_last_level_3__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[102]), .Z(
        buf_in_last_level_0__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[102]), .Z(
        buf_in_last_level_1__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[102]), .Z(
        buf_in_last_level_2__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[102]), .Z(
        buf_in_last_level_3__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[103]), .Z(
        buf_in_last_level_0__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[103]), .Z(
        buf_in_last_level_1__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[103]), .Z(
        buf_in_last_level_2__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[103]), .Z(
        buf_in_last_level_3__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[104]), .Z(
        buf_in_last_level_0__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[104]), .Z(
        buf_in_last_level_1__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[104]), .Z(
        buf_in_last_level_2__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[104]), .Z(
        buf_in_last_level_3__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[105]), .Z(
        buf_in_last_level_0__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[105]), .Z(
        buf_in_last_level_1__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[105]), .Z(
        buf_in_last_level_2__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[105]), .Z(
        buf_in_last_level_3__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[106]), .Z(
        buf_in_last_level_0__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[106]), .Z(
        buf_in_last_level_1__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[106]), .Z(
        buf_in_last_level_2__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[106]), .Z(
        buf_in_last_level_3__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[107]), .Z(
        buf_in_last_level_0__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[107]), .Z(
        buf_in_last_level_1__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[107]), .Z(
        buf_in_last_level_2__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[107]), .Z(
        buf_in_last_level_3__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[108]), .Z(
        buf_in_last_level_0__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[108]), .Z(
        buf_in_last_level_1__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[108]), .Z(
        buf_in_last_level_2__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[108]), .Z(
        buf_in_last_level_3__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[109]), .Z(
        buf_in_last_level_0__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[109]), .Z(
        buf_in_last_level_1__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[109]), .Z(
        buf_in_last_level_2__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[109]), .Z(
        buf_in_last_level_3__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[110]), .Z(
        buf_in_last_level_0__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[110]), .Z(
        buf_in_last_level_1__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[110]), .Z(
        buf_in_last_level_2__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[110]), .Z(
        buf_in_last_level_3__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[111]), .Z(
        buf_in_last_level_0__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[111]), .Z(
        buf_in_last_level_1__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[111]), .Z(
        buf_in_last_level_2__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[111]), .Z(
        buf_in_last_level_3__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[112]), .Z(
        buf_in_last_level_0__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[112]), .Z(
        buf_in_last_level_1__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[112]), .Z(
        buf_in_last_level_2__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[112]), .Z(
        buf_in_last_level_3__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[113]), .Z(
        buf_in_last_level_0__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[113]), .Z(
        buf_in_last_level_1__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[113]), .Z(
        buf_in_last_level_2__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[113]), .Z(
        buf_in_last_level_3__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[114]), .Z(
        buf_in_last_level_0__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[114]), .Z(
        buf_in_last_level_1__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[114]), .Z(
        buf_in_last_level_2__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[114]), .Z(
        buf_in_last_level_3__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[115]), .Z(
        buf_in_last_level_0__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[115]), .Z(
        buf_in_last_level_1__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[115]), .Z(
        buf_in_last_level_2__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[115]), .Z(
        buf_in_last_level_3__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[116]), .Z(
        buf_in_last_level_0__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[116]), .Z(
        buf_in_last_level_1__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[116]), .Z(
        buf_in_last_level_2__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[116]), .Z(
        buf_in_last_level_3__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[117]), .Z(
        buf_in_last_level_0__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[117]), .Z(
        buf_in_last_level_1__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[117]), .Z(
        buf_in_last_level_2__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[117]), .Z(
        buf_in_last_level_3__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[118]), .Z(
        buf_in_last_level_0__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[118]), .Z(
        buf_in_last_level_1__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[118]), .Z(
        buf_in_last_level_2__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[118]), .Z(
        buf_in_last_level_3__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[119]), .Z(
        buf_in_last_level_0__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[119]), .Z(
        buf_in_last_level_1__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[119]), .Z(
        buf_in_last_level_2__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[119]), .Z(
        buf_in_last_level_3__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[120]), .Z(
        buf_in_last_level_0__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[120]), .Z(
        buf_in_last_level_1__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[120]), .Z(
        buf_in_last_level_2__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[120]), .Z(
        buf_in_last_level_3__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[121]), .Z(
        buf_in_last_level_0__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[121]), .Z(
        buf_in_last_level_1__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[121]), .Z(
        buf_in_last_level_2__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[121]), .Z(
        buf_in_last_level_3__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[122]), .Z(
        buf_in_last_level_0__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[122]), .Z(
        buf_in_last_level_1__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[122]), .Z(
        buf_in_last_level_2__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[122]), .Z(
        buf_in_last_level_3__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[123]), .Z(
        buf_in_last_level_0__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[123]), .Z(
        buf_in_last_level_1__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[123]), .Z(
        buf_in_last_level_2__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[123]), .Z(
        buf_in_last_level_3__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[124]), .Z(
        buf_in_last_level_0__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[124]), .Z(
        buf_in_last_level_1__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[124]), .Z(
        buf_in_last_level_2__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[124]), .Z(
        buf_in_last_level_3__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[125]), .Z(
        buf_in_last_level_0__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[125]), .Z(
        buf_in_last_level_1__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[125]), .Z(
        buf_in_last_level_2__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[125]), .Z(
        buf_in_last_level_3__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[126]), .Z(
        buf_in_last_level_0__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[126]), .Z(
        buf_in_last_level_1__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[126]), .Z(
        buf_in_last_level_2__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[126]), .Z(
        buf_in_last_level_3__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[127]), .Z(
        buf_in_last_level_0__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[127]), .Z(
        buf_in_last_level_1__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[127]), .Z(
        buf_in_last_level_2__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[127]), .Z(
        buf_in_last_level_3__i_data_o_buf[127]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(CLK), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(CLK), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(CLK), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(CLK), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(CLK), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(CLK), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(CLK), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(CLK), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[101]), .Z(N469) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[102]), .Z(N470) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[105]), .Z(N473) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[107]), .Z(N475) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[109]), .Z(N477) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[110]), .Z(N478) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[111]), .Z(N479) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[112]), .Z(N480) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[115]), .Z(N483) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[82]), .Z(N416) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[86]), .Z(N420) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[61]), .Z(N361) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[63]), .Z(N363) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[30]), .Z(N296) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[22]), .Z(N288) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[21]), .Z(N287) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[20]), .Z(N286) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[23]), .Z(N289) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[24]), .Z(N290) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[25]), .Z(N291) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[26]), .Z(N292) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[27]), .Z(N293) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[28]), .Z(N294) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[29]), .Z(N295) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[31]), .Z(N297) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[37]), .Z(N337) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[19]), .Z(N285) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[18]), .Z(N284) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[17]), .Z(N283) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[16]), .Z(N282) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[15]), .Z(N281) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[14]), .Z(N280) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[13]), .Z(N279) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[12]), .Z(N278) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[11]), .Z(N277) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[10]), .Z(N276) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[9]), .Z(N275) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[8]), .Z(N274) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[7]), .Z(N273) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[5]), .Z(N271) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[4]), .Z(N270) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[3]), .Z(N269) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[1]), .Z(N267) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[0]), .Z(N266) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[62]), .Z(N362) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[60]), .Z(N360) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[59]), .Z(N359) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[57]), .Z(N357) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[56]), .Z(N356) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[55]), .Z(N355) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[54]), .Z(N354) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[53]), .Z(N353) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[52]), .Z(N352) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[51]), .Z(N351) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[50]), .Z(N350) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[49]), .Z(N349) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[48]), .Z(N348) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[47]), .Z(N347) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[46]), .Z(N346) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[45]), .Z(N345) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[44]), .Z(N344) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[43]), .Z(N343) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[42]), .Z(N342) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[41]), .Z(N341) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[40]), .Z(N340) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[39]), .Z(N339) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[38]), .Z(N338) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[58]), .Z(N358) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[64]), .Z(N398) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[65]), .Z(N399) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[66]), .Z(N400) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[67]), .Z(N401) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[68]), .Z(N402) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[69]), .Z(N403) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[70]), .Z(N404) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[71]), .Z(N405) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[72]), .Z(N406) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[73]), .Z(N407) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[74]), .Z(N408) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[75]), .Z(N409) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[76]), .Z(N410) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[77]), .Z(N411) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[78]), .Z(N412) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[79]), .Z(N413) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[80]), .Z(N414) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[81]), .Z(N415) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[83]), .Z(N417) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[84]), .Z(N418) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[85]), .Z(N419) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[87]), .Z(N421) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[88]), .Z(N422) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[89]), .Z(N423) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[90]), .Z(N424) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[91]), .Z(N425) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[92]), .Z(N426) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[93]), .Z(N427) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[94]), .Z(N428) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[95]), .Z(N429) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[32]), .Z(N332) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[33]), .Z(N333) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[34]), .Z(N334) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[35]), .Z(N335) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[36]), .Z(N336) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        CLK, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input CLK, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;
  wire   [127:0] buf_in_last_level_0__i_data_o_buf;
  wire   [127:0] buf_in_last_level_1__i_data_o_buf;
  wire   [127:0] buf_in_last_level_2__i_data_o_buf;
  wire   [127:0] buf_in_last_level_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[0]), .Z(
        buf_in_last_level_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[0]), .Z(
        buf_in_last_level_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[0]), .Z(
        buf_in_last_level_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[0]), .Z(
        buf_in_last_level_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[1]), .Z(
        buf_in_last_level_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[1]), .Z(
        buf_in_last_level_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[1]), .Z(
        buf_in_last_level_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[1]), .Z(
        buf_in_last_level_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[2]), .Z(
        buf_in_last_level_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[2]), .Z(
        buf_in_last_level_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[2]), .Z(
        buf_in_last_level_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[2]), .Z(
        buf_in_last_level_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[3]), .Z(
        buf_in_last_level_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[3]), .Z(
        buf_in_last_level_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[3]), .Z(
        buf_in_last_level_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[3]), .Z(
        buf_in_last_level_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[4]), .Z(
        buf_in_last_level_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[4]), .Z(
        buf_in_last_level_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[4]), .Z(
        buf_in_last_level_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[4]), .Z(
        buf_in_last_level_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[5]), .Z(
        buf_in_last_level_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[5]), .Z(
        buf_in_last_level_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[5]), .Z(
        buf_in_last_level_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[5]), .Z(
        buf_in_last_level_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[6]), .Z(
        buf_in_last_level_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[6]), .Z(
        buf_in_last_level_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[6]), .Z(
        buf_in_last_level_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[6]), .Z(
        buf_in_last_level_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[7]), .Z(
        buf_in_last_level_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[7]), .Z(
        buf_in_last_level_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[7]), .Z(
        buf_in_last_level_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[7]), .Z(
        buf_in_last_level_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[8]), .Z(
        buf_in_last_level_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[8]), .Z(
        buf_in_last_level_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[8]), .Z(
        buf_in_last_level_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[8]), .Z(
        buf_in_last_level_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[9]), .Z(
        buf_in_last_level_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[9]), .Z(
        buf_in_last_level_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[9]), .Z(
        buf_in_last_level_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[9]), .Z(
        buf_in_last_level_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[10]), .Z(
        buf_in_last_level_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[10]), .Z(
        buf_in_last_level_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[10]), .Z(
        buf_in_last_level_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[10]), .Z(
        buf_in_last_level_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[11]), .Z(
        buf_in_last_level_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[11]), .Z(
        buf_in_last_level_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[11]), .Z(
        buf_in_last_level_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[11]), .Z(
        buf_in_last_level_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[12]), .Z(
        buf_in_last_level_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[12]), .Z(
        buf_in_last_level_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[12]), .Z(
        buf_in_last_level_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[12]), .Z(
        buf_in_last_level_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[13]), .Z(
        buf_in_last_level_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[13]), .Z(
        buf_in_last_level_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[13]), .Z(
        buf_in_last_level_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[13]), .Z(
        buf_in_last_level_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[14]), .Z(
        buf_in_last_level_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[14]), .Z(
        buf_in_last_level_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[14]), .Z(
        buf_in_last_level_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[14]), .Z(
        buf_in_last_level_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[15]), .Z(
        buf_in_last_level_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[15]), .Z(
        buf_in_last_level_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[15]), .Z(
        buf_in_last_level_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[15]), .Z(
        buf_in_last_level_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[16]), .Z(
        buf_in_last_level_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[16]), .Z(
        buf_in_last_level_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[16]), .Z(
        buf_in_last_level_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[16]), .Z(
        buf_in_last_level_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[17]), .Z(
        buf_in_last_level_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[17]), .Z(
        buf_in_last_level_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[17]), .Z(
        buf_in_last_level_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[17]), .Z(
        buf_in_last_level_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[18]), .Z(
        buf_in_last_level_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[18]), .Z(
        buf_in_last_level_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[18]), .Z(
        buf_in_last_level_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[18]), .Z(
        buf_in_last_level_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[19]), .Z(
        buf_in_last_level_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[19]), .Z(
        buf_in_last_level_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[19]), .Z(
        buf_in_last_level_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[19]), .Z(
        buf_in_last_level_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[20]), .Z(
        buf_in_last_level_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[20]), .Z(
        buf_in_last_level_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[20]), .Z(
        buf_in_last_level_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[20]), .Z(
        buf_in_last_level_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[21]), .Z(
        buf_in_last_level_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[21]), .Z(
        buf_in_last_level_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[21]), .Z(
        buf_in_last_level_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[21]), .Z(
        buf_in_last_level_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[22]), .Z(
        buf_in_last_level_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[22]), .Z(
        buf_in_last_level_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[22]), .Z(
        buf_in_last_level_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[22]), .Z(
        buf_in_last_level_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[23]), .Z(
        buf_in_last_level_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[23]), .Z(
        buf_in_last_level_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[23]), .Z(
        buf_in_last_level_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[23]), .Z(
        buf_in_last_level_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[24]), .Z(
        buf_in_last_level_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[24]), .Z(
        buf_in_last_level_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[24]), .Z(
        buf_in_last_level_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[24]), .Z(
        buf_in_last_level_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[25]), .Z(
        buf_in_last_level_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[25]), .Z(
        buf_in_last_level_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[25]), .Z(
        buf_in_last_level_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[25]), .Z(
        buf_in_last_level_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[26]), .Z(
        buf_in_last_level_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[26]), .Z(
        buf_in_last_level_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[26]), .Z(
        buf_in_last_level_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[26]), .Z(
        buf_in_last_level_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[27]), .Z(
        buf_in_last_level_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[27]), .Z(
        buf_in_last_level_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[27]), .Z(
        buf_in_last_level_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[27]), .Z(
        buf_in_last_level_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[28]), .Z(
        buf_in_last_level_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[28]), .Z(
        buf_in_last_level_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[28]), .Z(
        buf_in_last_level_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[28]), .Z(
        buf_in_last_level_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[29]), .Z(
        buf_in_last_level_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[29]), .Z(
        buf_in_last_level_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[29]), .Z(
        buf_in_last_level_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[29]), .Z(
        buf_in_last_level_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[30]), .Z(
        buf_in_last_level_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[30]), .Z(
        buf_in_last_level_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[30]), .Z(
        buf_in_last_level_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[30]), .Z(
        buf_in_last_level_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[31]), .Z(
        buf_in_last_level_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[31]), .Z(
        buf_in_last_level_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[31]), .Z(
        buf_in_last_level_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[31]), .Z(
        buf_in_last_level_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[32]), .Z(
        buf_in_last_level_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[32]), .Z(
        buf_in_last_level_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[32]), .Z(
        buf_in_last_level_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[32]), .Z(
        buf_in_last_level_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[33]), .Z(
        buf_in_last_level_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[33]), .Z(
        buf_in_last_level_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[33]), .Z(
        buf_in_last_level_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[33]), .Z(
        buf_in_last_level_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[34]), .Z(
        buf_in_last_level_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[34]), .Z(
        buf_in_last_level_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[34]), .Z(
        buf_in_last_level_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[34]), .Z(
        buf_in_last_level_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[35]), .Z(
        buf_in_last_level_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[35]), .Z(
        buf_in_last_level_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[35]), .Z(
        buf_in_last_level_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[35]), .Z(
        buf_in_last_level_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[36]), .Z(
        buf_in_last_level_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[36]), .Z(
        buf_in_last_level_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[36]), .Z(
        buf_in_last_level_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[36]), .Z(
        buf_in_last_level_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[37]), .Z(
        buf_in_last_level_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[37]), .Z(
        buf_in_last_level_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[37]), .Z(
        buf_in_last_level_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[37]), .Z(
        buf_in_last_level_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[38]), .Z(
        buf_in_last_level_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[38]), .Z(
        buf_in_last_level_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[38]), .Z(
        buf_in_last_level_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[38]), .Z(
        buf_in_last_level_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[39]), .Z(
        buf_in_last_level_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[39]), .Z(
        buf_in_last_level_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[39]), .Z(
        buf_in_last_level_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[39]), .Z(
        buf_in_last_level_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[40]), .Z(
        buf_in_last_level_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[40]), .Z(
        buf_in_last_level_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[40]), .Z(
        buf_in_last_level_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[40]), .Z(
        buf_in_last_level_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[41]), .Z(
        buf_in_last_level_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[41]), .Z(
        buf_in_last_level_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[41]), .Z(
        buf_in_last_level_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[41]), .Z(
        buf_in_last_level_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[42]), .Z(
        buf_in_last_level_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[42]), .Z(
        buf_in_last_level_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[42]), .Z(
        buf_in_last_level_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[42]), .Z(
        buf_in_last_level_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[43]), .Z(
        buf_in_last_level_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[43]), .Z(
        buf_in_last_level_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[43]), .Z(
        buf_in_last_level_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[43]), .Z(
        buf_in_last_level_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[44]), .Z(
        buf_in_last_level_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[44]), .Z(
        buf_in_last_level_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[44]), .Z(
        buf_in_last_level_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[44]), .Z(
        buf_in_last_level_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[45]), .Z(
        buf_in_last_level_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[45]), .Z(
        buf_in_last_level_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[45]), .Z(
        buf_in_last_level_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[45]), .Z(
        buf_in_last_level_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[46]), .Z(
        buf_in_last_level_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[46]), .Z(
        buf_in_last_level_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[46]), .Z(
        buf_in_last_level_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[46]), .Z(
        buf_in_last_level_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[47]), .Z(
        buf_in_last_level_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[47]), .Z(
        buf_in_last_level_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[47]), .Z(
        buf_in_last_level_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[47]), .Z(
        buf_in_last_level_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[48]), .Z(
        buf_in_last_level_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[48]), .Z(
        buf_in_last_level_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[48]), .Z(
        buf_in_last_level_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[48]), .Z(
        buf_in_last_level_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[49]), .Z(
        buf_in_last_level_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[49]), .Z(
        buf_in_last_level_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[49]), .Z(
        buf_in_last_level_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[49]), .Z(
        buf_in_last_level_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[50]), .Z(
        buf_in_last_level_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[50]), .Z(
        buf_in_last_level_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[50]), .Z(
        buf_in_last_level_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[50]), .Z(
        buf_in_last_level_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[51]), .Z(
        buf_in_last_level_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[51]), .Z(
        buf_in_last_level_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[51]), .Z(
        buf_in_last_level_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[51]), .Z(
        buf_in_last_level_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[52]), .Z(
        buf_in_last_level_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[52]), .Z(
        buf_in_last_level_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[52]), .Z(
        buf_in_last_level_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[52]), .Z(
        buf_in_last_level_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[53]), .Z(
        buf_in_last_level_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[53]), .Z(
        buf_in_last_level_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[53]), .Z(
        buf_in_last_level_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[53]), .Z(
        buf_in_last_level_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[54]), .Z(
        buf_in_last_level_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[54]), .Z(
        buf_in_last_level_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[54]), .Z(
        buf_in_last_level_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[54]), .Z(
        buf_in_last_level_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[55]), .Z(
        buf_in_last_level_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[55]), .Z(
        buf_in_last_level_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[55]), .Z(
        buf_in_last_level_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[55]), .Z(
        buf_in_last_level_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[56]), .Z(
        buf_in_last_level_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[56]), .Z(
        buf_in_last_level_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[56]), .Z(
        buf_in_last_level_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[56]), .Z(
        buf_in_last_level_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[57]), .Z(
        buf_in_last_level_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[57]), .Z(
        buf_in_last_level_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[57]), .Z(
        buf_in_last_level_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[57]), .Z(
        buf_in_last_level_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[58]), .Z(
        buf_in_last_level_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[58]), .Z(
        buf_in_last_level_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[58]), .Z(
        buf_in_last_level_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[58]), .Z(
        buf_in_last_level_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[59]), .Z(
        buf_in_last_level_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[59]), .Z(
        buf_in_last_level_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[59]), .Z(
        buf_in_last_level_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[59]), .Z(
        buf_in_last_level_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[60]), .Z(
        buf_in_last_level_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[60]), .Z(
        buf_in_last_level_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[60]), .Z(
        buf_in_last_level_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[60]), .Z(
        buf_in_last_level_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[61]), .Z(
        buf_in_last_level_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[61]), .Z(
        buf_in_last_level_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[61]), .Z(
        buf_in_last_level_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[61]), .Z(
        buf_in_last_level_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[62]), .Z(
        buf_in_last_level_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[62]), .Z(
        buf_in_last_level_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[62]), .Z(
        buf_in_last_level_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[62]), .Z(
        buf_in_last_level_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[63]), .Z(
        buf_in_last_level_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[63]), .Z(
        buf_in_last_level_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[63]), .Z(
        buf_in_last_level_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[63]), .Z(
        buf_in_last_level_3__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[64]), .Z(
        buf_in_last_level_0__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[64]), .Z(
        buf_in_last_level_1__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[64]), .Z(
        buf_in_last_level_2__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[64]), .Z(
        buf_in_last_level_3__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[65]), .Z(
        buf_in_last_level_0__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[65]), .Z(
        buf_in_last_level_1__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[65]), .Z(
        buf_in_last_level_2__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[65]), .Z(
        buf_in_last_level_3__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[66]), .Z(
        buf_in_last_level_0__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[66]), .Z(
        buf_in_last_level_1__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[66]), .Z(
        buf_in_last_level_2__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[66]), .Z(
        buf_in_last_level_3__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[67]), .Z(
        buf_in_last_level_0__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[67]), .Z(
        buf_in_last_level_1__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[67]), .Z(
        buf_in_last_level_2__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[67]), .Z(
        buf_in_last_level_3__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[68]), .Z(
        buf_in_last_level_0__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[68]), .Z(
        buf_in_last_level_1__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[68]), .Z(
        buf_in_last_level_2__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[68]), .Z(
        buf_in_last_level_3__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[69]), .Z(
        buf_in_last_level_0__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[69]), .Z(
        buf_in_last_level_1__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[69]), .Z(
        buf_in_last_level_2__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[69]), .Z(
        buf_in_last_level_3__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[70]), .Z(
        buf_in_last_level_0__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[70]), .Z(
        buf_in_last_level_1__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[70]), .Z(
        buf_in_last_level_2__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[70]), .Z(
        buf_in_last_level_3__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[71]), .Z(
        buf_in_last_level_0__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[71]), .Z(
        buf_in_last_level_1__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[71]), .Z(
        buf_in_last_level_2__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[71]), .Z(
        buf_in_last_level_3__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[72]), .Z(
        buf_in_last_level_0__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[72]), .Z(
        buf_in_last_level_1__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[72]), .Z(
        buf_in_last_level_2__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[72]), .Z(
        buf_in_last_level_3__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[73]), .Z(
        buf_in_last_level_0__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[73]), .Z(
        buf_in_last_level_1__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[73]), .Z(
        buf_in_last_level_2__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[73]), .Z(
        buf_in_last_level_3__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[74]), .Z(
        buf_in_last_level_0__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[74]), .Z(
        buf_in_last_level_1__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[74]), .Z(
        buf_in_last_level_2__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[74]), .Z(
        buf_in_last_level_3__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[75]), .Z(
        buf_in_last_level_0__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[75]), .Z(
        buf_in_last_level_1__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[75]), .Z(
        buf_in_last_level_2__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[75]), .Z(
        buf_in_last_level_3__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[76]), .Z(
        buf_in_last_level_0__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[76]), .Z(
        buf_in_last_level_1__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[76]), .Z(
        buf_in_last_level_2__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[76]), .Z(
        buf_in_last_level_3__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[77]), .Z(
        buf_in_last_level_0__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[77]), .Z(
        buf_in_last_level_1__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[77]), .Z(
        buf_in_last_level_2__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[77]), .Z(
        buf_in_last_level_3__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[78]), .Z(
        buf_in_last_level_0__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[78]), .Z(
        buf_in_last_level_1__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[78]), .Z(
        buf_in_last_level_2__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[78]), .Z(
        buf_in_last_level_3__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[79]), .Z(
        buf_in_last_level_0__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[79]), .Z(
        buf_in_last_level_1__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[79]), .Z(
        buf_in_last_level_2__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[79]), .Z(
        buf_in_last_level_3__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[80]), .Z(
        buf_in_last_level_0__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[80]), .Z(
        buf_in_last_level_1__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[80]), .Z(
        buf_in_last_level_2__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[80]), .Z(
        buf_in_last_level_3__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[81]), .Z(
        buf_in_last_level_0__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[81]), .Z(
        buf_in_last_level_1__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[81]), .Z(
        buf_in_last_level_2__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[81]), .Z(
        buf_in_last_level_3__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[82]), .Z(
        buf_in_last_level_0__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[82]), .Z(
        buf_in_last_level_1__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[82]), .Z(
        buf_in_last_level_2__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[82]), .Z(
        buf_in_last_level_3__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[83]), .Z(
        buf_in_last_level_0__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[83]), .Z(
        buf_in_last_level_1__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[83]), .Z(
        buf_in_last_level_2__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[83]), .Z(
        buf_in_last_level_3__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[84]), .Z(
        buf_in_last_level_0__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[84]), .Z(
        buf_in_last_level_1__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[84]), .Z(
        buf_in_last_level_2__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[84]), .Z(
        buf_in_last_level_3__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[85]), .Z(
        buf_in_last_level_0__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[85]), .Z(
        buf_in_last_level_1__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[85]), .Z(
        buf_in_last_level_2__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[85]), .Z(
        buf_in_last_level_3__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[86]), .Z(
        buf_in_last_level_0__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[86]), .Z(
        buf_in_last_level_1__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[86]), .Z(
        buf_in_last_level_2__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[86]), .Z(
        buf_in_last_level_3__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[87]), .Z(
        buf_in_last_level_0__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[87]), .Z(
        buf_in_last_level_1__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[87]), .Z(
        buf_in_last_level_2__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[87]), .Z(
        buf_in_last_level_3__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[88]), .Z(
        buf_in_last_level_0__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[88]), .Z(
        buf_in_last_level_1__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[88]), .Z(
        buf_in_last_level_2__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[88]), .Z(
        buf_in_last_level_3__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[89]), .Z(
        buf_in_last_level_0__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[89]), .Z(
        buf_in_last_level_1__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[89]), .Z(
        buf_in_last_level_2__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[89]), .Z(
        buf_in_last_level_3__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[90]), .Z(
        buf_in_last_level_0__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[90]), .Z(
        buf_in_last_level_1__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[90]), .Z(
        buf_in_last_level_2__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[90]), .Z(
        buf_in_last_level_3__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[91]), .Z(
        buf_in_last_level_0__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[91]), .Z(
        buf_in_last_level_1__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[91]), .Z(
        buf_in_last_level_2__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[91]), .Z(
        buf_in_last_level_3__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[92]), .Z(
        buf_in_last_level_0__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[92]), .Z(
        buf_in_last_level_1__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[92]), .Z(
        buf_in_last_level_2__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[92]), .Z(
        buf_in_last_level_3__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[93]), .Z(
        buf_in_last_level_0__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[93]), .Z(
        buf_in_last_level_1__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[93]), .Z(
        buf_in_last_level_2__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[93]), .Z(
        buf_in_last_level_3__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[94]), .Z(
        buf_in_last_level_0__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[94]), .Z(
        buf_in_last_level_1__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[94]), .Z(
        buf_in_last_level_2__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[94]), .Z(
        buf_in_last_level_3__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[95]), .Z(
        buf_in_last_level_0__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[95]), .Z(
        buf_in_last_level_1__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[95]), .Z(
        buf_in_last_level_2__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[95]), .Z(
        buf_in_last_level_3__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[96]), .Z(
        buf_in_last_level_0__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[96]), .Z(
        buf_in_last_level_1__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[96]), .Z(
        buf_in_last_level_2__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[96]), .Z(
        buf_in_last_level_3__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[97]), .Z(
        buf_in_last_level_0__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[97]), .Z(
        buf_in_last_level_1__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[97]), .Z(
        buf_in_last_level_2__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[97]), .Z(
        buf_in_last_level_3__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[98]), .Z(
        buf_in_last_level_0__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[98]), .Z(
        buf_in_last_level_1__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[98]), .Z(
        buf_in_last_level_2__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[98]), .Z(
        buf_in_last_level_3__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[99]), .Z(
        buf_in_last_level_0__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[99]), .Z(
        buf_in_last_level_1__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[99]), .Z(
        buf_in_last_level_2__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[99]), .Z(
        buf_in_last_level_3__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[100]), .Z(
        buf_in_last_level_0__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[100]), .Z(
        buf_in_last_level_1__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[100]), .Z(
        buf_in_last_level_2__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[100]), .Z(
        buf_in_last_level_3__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[101]), .Z(
        buf_in_last_level_0__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[101]), .Z(
        buf_in_last_level_1__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[101]), .Z(
        buf_in_last_level_2__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[101]), .Z(
        buf_in_last_level_3__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[102]), .Z(
        buf_in_last_level_0__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[102]), .Z(
        buf_in_last_level_1__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[102]), .Z(
        buf_in_last_level_2__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[102]), .Z(
        buf_in_last_level_3__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[103]), .Z(
        buf_in_last_level_0__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[103]), .Z(
        buf_in_last_level_1__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[103]), .Z(
        buf_in_last_level_2__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[103]), .Z(
        buf_in_last_level_3__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[104]), .Z(
        buf_in_last_level_0__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[104]), .Z(
        buf_in_last_level_1__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[104]), .Z(
        buf_in_last_level_2__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[104]), .Z(
        buf_in_last_level_3__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[105]), .Z(
        buf_in_last_level_0__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[105]), .Z(
        buf_in_last_level_1__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[105]), .Z(
        buf_in_last_level_2__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[105]), .Z(
        buf_in_last_level_3__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[106]), .Z(
        buf_in_last_level_0__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[106]), .Z(
        buf_in_last_level_1__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[106]), .Z(
        buf_in_last_level_2__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[106]), .Z(
        buf_in_last_level_3__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[107]), .Z(
        buf_in_last_level_0__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[107]), .Z(
        buf_in_last_level_1__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[107]), .Z(
        buf_in_last_level_2__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[107]), .Z(
        buf_in_last_level_3__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[108]), .Z(
        buf_in_last_level_0__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[108]), .Z(
        buf_in_last_level_1__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[108]), .Z(
        buf_in_last_level_2__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[108]), .Z(
        buf_in_last_level_3__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[109]), .Z(
        buf_in_last_level_0__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[109]), .Z(
        buf_in_last_level_1__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[109]), .Z(
        buf_in_last_level_2__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[109]), .Z(
        buf_in_last_level_3__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[110]), .Z(
        buf_in_last_level_0__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[110]), .Z(
        buf_in_last_level_1__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[110]), .Z(
        buf_in_last_level_2__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[110]), .Z(
        buf_in_last_level_3__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[111]), .Z(
        buf_in_last_level_0__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[111]), .Z(
        buf_in_last_level_1__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[111]), .Z(
        buf_in_last_level_2__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[111]), .Z(
        buf_in_last_level_3__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[112]), .Z(
        buf_in_last_level_0__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[112]), .Z(
        buf_in_last_level_1__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[112]), .Z(
        buf_in_last_level_2__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[112]), .Z(
        buf_in_last_level_3__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[113]), .Z(
        buf_in_last_level_0__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[113]), .Z(
        buf_in_last_level_1__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[113]), .Z(
        buf_in_last_level_2__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[113]), .Z(
        buf_in_last_level_3__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[114]), .Z(
        buf_in_last_level_0__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[114]), .Z(
        buf_in_last_level_1__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[114]), .Z(
        buf_in_last_level_2__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[114]), .Z(
        buf_in_last_level_3__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[115]), .Z(
        buf_in_last_level_0__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[115]), .Z(
        buf_in_last_level_1__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[115]), .Z(
        buf_in_last_level_2__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[115]), .Z(
        buf_in_last_level_3__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[116]), .Z(
        buf_in_last_level_0__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[116]), .Z(
        buf_in_last_level_1__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[116]), .Z(
        buf_in_last_level_2__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[116]), .Z(
        buf_in_last_level_3__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[117]), .Z(
        buf_in_last_level_0__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[117]), .Z(
        buf_in_last_level_1__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[117]), .Z(
        buf_in_last_level_2__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[117]), .Z(
        buf_in_last_level_3__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[118]), .Z(
        buf_in_last_level_0__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[118]), .Z(
        buf_in_last_level_1__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[118]), .Z(
        buf_in_last_level_2__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[118]), .Z(
        buf_in_last_level_3__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[119]), .Z(
        buf_in_last_level_0__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[119]), .Z(
        buf_in_last_level_1__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[119]), .Z(
        buf_in_last_level_2__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[119]), .Z(
        buf_in_last_level_3__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[120]), .Z(
        buf_in_last_level_0__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[120]), .Z(
        buf_in_last_level_1__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[120]), .Z(
        buf_in_last_level_2__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[120]), .Z(
        buf_in_last_level_3__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[121]), .Z(
        buf_in_last_level_0__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[121]), .Z(
        buf_in_last_level_1__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[121]), .Z(
        buf_in_last_level_2__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[121]), .Z(
        buf_in_last_level_3__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[122]), .Z(
        buf_in_last_level_0__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[122]), .Z(
        buf_in_last_level_1__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[122]), .Z(
        buf_in_last_level_2__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[122]), .Z(
        buf_in_last_level_3__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[123]), .Z(
        buf_in_last_level_0__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[123]), .Z(
        buf_in_last_level_1__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[123]), .Z(
        buf_in_last_level_2__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[123]), .Z(
        buf_in_last_level_3__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[124]), .Z(
        buf_in_last_level_0__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[124]), .Z(
        buf_in_last_level_1__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[124]), .Z(
        buf_in_last_level_2__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[124]), .Z(
        buf_in_last_level_3__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[125]), .Z(
        buf_in_last_level_0__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[125]), .Z(
        buf_in_last_level_1__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[125]), .Z(
        buf_in_last_level_2__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[125]), .Z(
        buf_in_last_level_3__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[126]), .Z(
        buf_in_last_level_0__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[126]), .Z(
        buf_in_last_level_1__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[126]), .Z(
        buf_in_last_level_2__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[126]), .Z(
        buf_in_last_level_3__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[127]), .Z(
        buf_in_last_level_0__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[127]), .Z(
        buf_in_last_level_1__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[127]), .Z(
        buf_in_last_level_2__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[127]), .Z(
        buf_in_last_level_3__i_data_o_buf[127]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(CLK), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(CLK), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(CLK), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(CLK), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(CLK), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(CLK), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(CLK), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(CLK), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[101]), .Z(N469) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[102]), .Z(N470) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[105]), .Z(N473) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[107]), .Z(N475) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[109]), .Z(N477) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[110]), .Z(N478) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[111]), .Z(N479) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[112]), .Z(N480) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[115]), .Z(N483) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[82]), .Z(N416) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[86]), .Z(N420) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[61]), .Z(N361) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[63]), .Z(N363) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[22]), .Z(N288) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[23]), .Z(N289) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[24]), .Z(N290) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[25]), .Z(N291) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[26]), .Z(N292) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[27]), .Z(N293) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[28]), .Z(N294) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[30]), .Z(N296) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[31]), .Z(N297) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[29]), .Z(N295) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[21]), .Z(N287) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[20]), .Z(N286) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[19]), .Z(N285) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[18]), .Z(N284) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[17]), .Z(N283) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[16]), .Z(N282) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[15]), .Z(N281) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[14]), .Z(N280) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[13]), .Z(N279) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[12]), .Z(N278) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[11]), .Z(N277) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[10]), .Z(N276) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[9]), .Z(N275) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[8]), .Z(N274) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[7]), .Z(N273) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[5]), .Z(N271) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[4]), .Z(N270) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[3]), .Z(N269) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[1]), .Z(N267) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[0]), .Z(N266) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[54]), .Z(N354) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[51]), .Z(N351) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[50]), .Z(N350) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[38]), .Z(N338) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[49]), .Z(N349) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[48]), .Z(N348) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[47]), .Z(N347) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[46]), .Z(N346) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[45]), .Z(N345) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[44]), .Z(N344) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[43]), .Z(N343) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[42]), .Z(N342) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[41]), .Z(N341) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[39]), .Z(N339) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[57]), .Z(N357) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[37]), .Z(N337) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[58]), .Z(N358) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[59]), .Z(N359) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[55]), .Z(N355) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[56]), .Z(N356) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[53]), .Z(N353) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[62]), .Z(N362) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[40]), .Z(N340) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[52]), .Z(N352) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[60]), .Z(N360) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[36]), .Z(N336) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[35]), .Z(N335) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[34]), .Z(N334) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[33]), .Z(N333) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[32]), .Z(N332) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[83]), .Z(N417) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[84]), .Z(N418) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[85]), .Z(N419) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[87]), .Z(N421) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[88]), .Z(N422) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[89]), .Z(N423) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[90]), .Z(N424) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[91]), .Z(N425) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[92]), .Z(N426) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[94]), .Z(N428) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[95]), .Z(N429) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[93]), .Z(N427) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[65]), .Z(N399) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[66]), .Z(N400) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[67]), .Z(N401) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[68]), .Z(N402) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[69]), .Z(N403) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[70]), .Z(N404) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[71]), .Z(N405) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[72]), .Z(N406) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[73]), .Z(N407) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[74]), .Z(N408) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[75]), .Z(N409) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[76]), .Z(N410) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[77]), .Z(N411) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[78]), .Z(N412) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[79]), .Z(N413) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[80]), .Z(N414) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[81]), .Z(N415) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[64]), .Z(N398) );
endmodule



    module wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        CLK, rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en );
  input [0:0] i_valid;
  input [31:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input CLK, rst, i_en;
  wire   wire_tree_level_0__i_valid_latch_0_, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N101, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N167, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N233, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N299, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N365, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N431, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N497, n1;
  wire   [31:0] wire_tree_level_0__i_data_latch;
  wire   [63:0] wire_tree_level_1__i_data_latch;
  wire   [1:0] wire_tree_level_1__i_valid_latch;
  wire   [127:0] wire_tree_level_2__i_data_latch;
  wire   [3:0] wire_tree_level_2__i_valid_latch;
  wire   [127:0] buf_in_last_level_0__i_data_o_buf;
  wire   [127:0] buf_in_last_level_1__i_data_o_buf;
  wire   [127:0] buf_in_last_level_2__i_data_o_buf;
  wire   [127:0] buf_in_last_level_3__i_data_o_buf;

  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[0]), .Z(
        buf_in_last_level_0__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[0]), .Z(
        buf_in_last_level_1__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[0]), .Z(
        buf_in_last_level_2__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_0__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[0]), .Z(
        buf_in_last_level_3__i_data_o_buf[0]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[1]), .Z(
        buf_in_last_level_0__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[1]), .Z(
        buf_in_last_level_1__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[1]), .Z(
        buf_in_last_level_2__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_1__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[1]), .Z(
        buf_in_last_level_3__i_data_o_buf[1]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[2]), .Z(
        buf_in_last_level_0__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[2]), .Z(
        buf_in_last_level_1__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[2]), .Z(
        buf_in_last_level_2__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_2__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[2]), .Z(
        buf_in_last_level_3__i_data_o_buf[2]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[3]), .Z(
        buf_in_last_level_0__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[3]), .Z(
        buf_in_last_level_1__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[3]), .Z(
        buf_in_last_level_2__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_3__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[3]), .Z(
        buf_in_last_level_3__i_data_o_buf[3]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[4]), .Z(
        buf_in_last_level_0__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[4]), .Z(
        buf_in_last_level_1__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[4]), .Z(
        buf_in_last_level_2__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_4__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[4]), .Z(
        buf_in_last_level_3__i_data_o_buf[4]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[5]), .Z(
        buf_in_last_level_0__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[5]), .Z(
        buf_in_last_level_1__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[5]), .Z(
        buf_in_last_level_2__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_5__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[5]), .Z(
        buf_in_last_level_3__i_data_o_buf[5]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[6]), .Z(
        buf_in_last_level_0__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[6]), .Z(
        buf_in_last_level_1__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[6]), .Z(
        buf_in_last_level_2__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_6__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[6]), .Z(
        buf_in_last_level_3__i_data_o_buf[6]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[7]), .Z(
        buf_in_last_level_0__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[7]), .Z(
        buf_in_last_level_1__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[7]), .Z(
        buf_in_last_level_2__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_7__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[7]), .Z(
        buf_in_last_level_3__i_data_o_buf[7]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[8]), .Z(
        buf_in_last_level_0__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[8]), .Z(
        buf_in_last_level_1__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[8]), .Z(
        buf_in_last_level_2__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_8__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[8]), .Z(
        buf_in_last_level_3__i_data_o_buf[8]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[9]), .Z(
        buf_in_last_level_0__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[9]), .Z(
        buf_in_last_level_1__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[9]), .Z(
        buf_in_last_level_2__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_9__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[9]), .Z(
        buf_in_last_level_3__i_data_o_buf[9]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[10]), .Z(
        buf_in_last_level_0__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[10]), .Z(
        buf_in_last_level_1__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[10]), .Z(
        buf_in_last_level_2__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_10__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[10]), .Z(
        buf_in_last_level_3__i_data_o_buf[10]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[11]), .Z(
        buf_in_last_level_0__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[11]), .Z(
        buf_in_last_level_1__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[11]), .Z(
        buf_in_last_level_2__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_11__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[11]), .Z(
        buf_in_last_level_3__i_data_o_buf[11]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[12]), .Z(
        buf_in_last_level_0__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[12]), .Z(
        buf_in_last_level_1__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[12]), .Z(
        buf_in_last_level_2__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_12__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[12]), .Z(
        buf_in_last_level_3__i_data_o_buf[12]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[13]), .Z(
        buf_in_last_level_0__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[13]), .Z(
        buf_in_last_level_1__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[13]), .Z(
        buf_in_last_level_2__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_13__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[13]), .Z(
        buf_in_last_level_3__i_data_o_buf[13]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[14]), .Z(
        buf_in_last_level_0__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[14]), .Z(
        buf_in_last_level_1__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[14]), .Z(
        buf_in_last_level_2__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_14__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[14]), .Z(
        buf_in_last_level_3__i_data_o_buf[14]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[15]), .Z(
        buf_in_last_level_0__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[15]), .Z(
        buf_in_last_level_1__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[15]), .Z(
        buf_in_last_level_2__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_15__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[15]), .Z(
        buf_in_last_level_3__i_data_o_buf[15]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[16]), .Z(
        buf_in_last_level_0__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[16]), .Z(
        buf_in_last_level_1__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[16]), .Z(
        buf_in_last_level_2__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_16__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[16]), .Z(
        buf_in_last_level_3__i_data_o_buf[16]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[17]), .Z(
        buf_in_last_level_0__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[17]), .Z(
        buf_in_last_level_1__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[17]), .Z(
        buf_in_last_level_2__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_17__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[17]), .Z(
        buf_in_last_level_3__i_data_o_buf[17]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[18]), .Z(
        buf_in_last_level_0__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[18]), .Z(
        buf_in_last_level_1__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[18]), .Z(
        buf_in_last_level_2__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_18__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[18]), .Z(
        buf_in_last_level_3__i_data_o_buf[18]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[19]), .Z(
        buf_in_last_level_0__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[19]), .Z(
        buf_in_last_level_1__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[19]), .Z(
        buf_in_last_level_2__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_19__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[19]), .Z(
        buf_in_last_level_3__i_data_o_buf[19]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[20]), .Z(
        buf_in_last_level_0__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[20]), .Z(
        buf_in_last_level_1__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[20]), .Z(
        buf_in_last_level_2__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_20__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[20]), .Z(
        buf_in_last_level_3__i_data_o_buf[20]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[21]), .Z(
        buf_in_last_level_0__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[21]), .Z(
        buf_in_last_level_1__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[21]), .Z(
        buf_in_last_level_2__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_21__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[21]), .Z(
        buf_in_last_level_3__i_data_o_buf[21]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[22]), .Z(
        buf_in_last_level_0__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[22]), .Z(
        buf_in_last_level_1__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[22]), .Z(
        buf_in_last_level_2__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_22__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[22]), .Z(
        buf_in_last_level_3__i_data_o_buf[22]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[23]), .Z(
        buf_in_last_level_0__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[23]), .Z(
        buf_in_last_level_1__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[23]), .Z(
        buf_in_last_level_2__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_23__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[23]), .Z(
        buf_in_last_level_3__i_data_o_buf[23]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[24]), .Z(
        buf_in_last_level_0__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[24]), .Z(
        buf_in_last_level_1__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[24]), .Z(
        buf_in_last_level_2__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_24__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[24]), .Z(
        buf_in_last_level_3__i_data_o_buf[24]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[25]), .Z(
        buf_in_last_level_0__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[25]), .Z(
        buf_in_last_level_1__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[25]), .Z(
        buf_in_last_level_2__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_25__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[25]), .Z(
        buf_in_last_level_3__i_data_o_buf[25]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[26]), .Z(
        buf_in_last_level_0__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[26]), .Z(
        buf_in_last_level_1__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[26]), .Z(
        buf_in_last_level_2__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_26__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[26]), .Z(
        buf_in_last_level_3__i_data_o_buf[26]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[27]), .Z(
        buf_in_last_level_0__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[27]), .Z(
        buf_in_last_level_1__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[27]), .Z(
        buf_in_last_level_2__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_27__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[27]), .Z(
        buf_in_last_level_3__i_data_o_buf[27]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[28]), .Z(
        buf_in_last_level_0__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[28]), .Z(
        buf_in_last_level_1__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[28]), .Z(
        buf_in_last_level_2__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_28__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[28]), .Z(
        buf_in_last_level_3__i_data_o_buf[28]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[29]), .Z(
        buf_in_last_level_0__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[29]), .Z(
        buf_in_last_level_1__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[29]), .Z(
        buf_in_last_level_2__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_29__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[29]), .Z(
        buf_in_last_level_3__i_data_o_buf[29]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[30]), .Z(
        buf_in_last_level_0__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[30]), .Z(
        buf_in_last_level_1__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[30]), .Z(
        buf_in_last_level_2__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_30__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[30]), .Z(
        buf_in_last_level_3__i_data_o_buf[30]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[31]), .Z(
        buf_in_last_level_0__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[31]), .Z(
        buf_in_last_level_1__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[31]), .Z(
        buf_in_last_level_2__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_31__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[31]), .Z(
        buf_in_last_level_3__i_data_o_buf[31]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[32]), .Z(
        buf_in_last_level_0__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[32]), .Z(
        buf_in_last_level_1__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[32]), .Z(
        buf_in_last_level_2__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_32__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[32]), .Z(
        buf_in_last_level_3__i_data_o_buf[32]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[33]), .Z(
        buf_in_last_level_0__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[33]), .Z(
        buf_in_last_level_1__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[33]), .Z(
        buf_in_last_level_2__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_33__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[33]), .Z(
        buf_in_last_level_3__i_data_o_buf[33]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[34]), .Z(
        buf_in_last_level_0__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[34]), .Z(
        buf_in_last_level_1__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[34]), .Z(
        buf_in_last_level_2__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_34__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[34]), .Z(
        buf_in_last_level_3__i_data_o_buf[34]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[35]), .Z(
        buf_in_last_level_0__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[35]), .Z(
        buf_in_last_level_1__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[35]), .Z(
        buf_in_last_level_2__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_35__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[35]), .Z(
        buf_in_last_level_3__i_data_o_buf[35]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[36]), .Z(
        buf_in_last_level_0__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[36]), .Z(
        buf_in_last_level_1__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[36]), .Z(
        buf_in_last_level_2__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_36__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[36]), .Z(
        buf_in_last_level_3__i_data_o_buf[36]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[37]), .Z(
        buf_in_last_level_0__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[37]), .Z(
        buf_in_last_level_1__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[37]), .Z(
        buf_in_last_level_2__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_37__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[37]), .Z(
        buf_in_last_level_3__i_data_o_buf[37]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[38]), .Z(
        buf_in_last_level_0__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[38]), .Z(
        buf_in_last_level_1__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[38]), .Z(
        buf_in_last_level_2__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_38__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[38]), .Z(
        buf_in_last_level_3__i_data_o_buf[38]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[39]), .Z(
        buf_in_last_level_0__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[39]), .Z(
        buf_in_last_level_1__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[39]), .Z(
        buf_in_last_level_2__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_39__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[39]), .Z(
        buf_in_last_level_3__i_data_o_buf[39]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[40]), .Z(
        buf_in_last_level_0__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[40]), .Z(
        buf_in_last_level_1__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[40]), .Z(
        buf_in_last_level_2__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_40__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[40]), .Z(
        buf_in_last_level_3__i_data_o_buf[40]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[41]), .Z(
        buf_in_last_level_0__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[41]), .Z(
        buf_in_last_level_1__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[41]), .Z(
        buf_in_last_level_2__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_41__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[41]), .Z(
        buf_in_last_level_3__i_data_o_buf[41]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[42]), .Z(
        buf_in_last_level_0__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[42]), .Z(
        buf_in_last_level_1__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[42]), .Z(
        buf_in_last_level_2__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_42__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[42]), .Z(
        buf_in_last_level_3__i_data_o_buf[42]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[43]), .Z(
        buf_in_last_level_0__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[43]), .Z(
        buf_in_last_level_1__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[43]), .Z(
        buf_in_last_level_2__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_43__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[43]), .Z(
        buf_in_last_level_3__i_data_o_buf[43]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[44]), .Z(
        buf_in_last_level_0__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[44]), .Z(
        buf_in_last_level_1__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[44]), .Z(
        buf_in_last_level_2__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_44__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[44]), .Z(
        buf_in_last_level_3__i_data_o_buf[44]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[45]), .Z(
        buf_in_last_level_0__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[45]), .Z(
        buf_in_last_level_1__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[45]), .Z(
        buf_in_last_level_2__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_45__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[45]), .Z(
        buf_in_last_level_3__i_data_o_buf[45]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[46]), .Z(
        buf_in_last_level_0__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[46]), .Z(
        buf_in_last_level_1__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[46]), .Z(
        buf_in_last_level_2__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_46__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[46]), .Z(
        buf_in_last_level_3__i_data_o_buf[46]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[47]), .Z(
        buf_in_last_level_0__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[47]), .Z(
        buf_in_last_level_1__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[47]), .Z(
        buf_in_last_level_2__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_47__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[47]), .Z(
        buf_in_last_level_3__i_data_o_buf[47]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[48]), .Z(
        buf_in_last_level_0__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[48]), .Z(
        buf_in_last_level_1__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[48]), .Z(
        buf_in_last_level_2__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_48__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[48]), .Z(
        buf_in_last_level_3__i_data_o_buf[48]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[49]), .Z(
        buf_in_last_level_0__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[49]), .Z(
        buf_in_last_level_1__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[49]), .Z(
        buf_in_last_level_2__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_49__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[49]), .Z(
        buf_in_last_level_3__i_data_o_buf[49]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[50]), .Z(
        buf_in_last_level_0__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[50]), .Z(
        buf_in_last_level_1__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[50]), .Z(
        buf_in_last_level_2__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_50__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[50]), .Z(
        buf_in_last_level_3__i_data_o_buf[50]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[51]), .Z(
        buf_in_last_level_0__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[51]), .Z(
        buf_in_last_level_1__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[51]), .Z(
        buf_in_last_level_2__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_51__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[51]), .Z(
        buf_in_last_level_3__i_data_o_buf[51]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[52]), .Z(
        buf_in_last_level_0__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[52]), .Z(
        buf_in_last_level_1__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[52]), .Z(
        buf_in_last_level_2__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_52__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[52]), .Z(
        buf_in_last_level_3__i_data_o_buf[52]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[53]), .Z(
        buf_in_last_level_0__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[53]), .Z(
        buf_in_last_level_1__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[53]), .Z(
        buf_in_last_level_2__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_53__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[53]), .Z(
        buf_in_last_level_3__i_data_o_buf[53]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[54]), .Z(
        buf_in_last_level_0__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[54]), .Z(
        buf_in_last_level_1__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[54]), .Z(
        buf_in_last_level_2__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_54__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[54]), .Z(
        buf_in_last_level_3__i_data_o_buf[54]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[55]), .Z(
        buf_in_last_level_0__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[55]), .Z(
        buf_in_last_level_1__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[55]), .Z(
        buf_in_last_level_2__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_55__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[55]), .Z(
        buf_in_last_level_3__i_data_o_buf[55]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[56]), .Z(
        buf_in_last_level_0__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[56]), .Z(
        buf_in_last_level_1__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[56]), .Z(
        buf_in_last_level_2__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_56__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[56]), .Z(
        buf_in_last_level_3__i_data_o_buf[56]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[57]), .Z(
        buf_in_last_level_0__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[57]), .Z(
        buf_in_last_level_1__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[57]), .Z(
        buf_in_last_level_2__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_57__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[57]), .Z(
        buf_in_last_level_3__i_data_o_buf[57]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[58]), .Z(
        buf_in_last_level_0__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[58]), .Z(
        buf_in_last_level_1__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[58]), .Z(
        buf_in_last_level_2__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_58__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[58]), .Z(
        buf_in_last_level_3__i_data_o_buf[58]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[59]), .Z(
        buf_in_last_level_0__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[59]), .Z(
        buf_in_last_level_1__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[59]), .Z(
        buf_in_last_level_2__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_59__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[59]), .Z(
        buf_in_last_level_3__i_data_o_buf[59]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[60]), .Z(
        buf_in_last_level_0__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[60]), .Z(
        buf_in_last_level_1__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[60]), .Z(
        buf_in_last_level_2__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_60__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[60]), .Z(
        buf_in_last_level_3__i_data_o_buf[60]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[61]), .Z(
        buf_in_last_level_0__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[61]), .Z(
        buf_in_last_level_1__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[61]), .Z(
        buf_in_last_level_2__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_61__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[61]), .Z(
        buf_in_last_level_3__i_data_o_buf[61]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[62]), .Z(
        buf_in_last_level_0__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[62]), .Z(
        buf_in_last_level_1__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[62]), .Z(
        buf_in_last_level_2__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_62__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[62]), .Z(
        buf_in_last_level_3__i_data_o_buf[62]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[63]), .Z(
        buf_in_last_level_0__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[63]), .Z(
        buf_in_last_level_1__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[63]), .Z(
        buf_in_last_level_2__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_63__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[63]), .Z(
        buf_in_last_level_3__i_data_o_buf[63]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[64]), .Z(
        buf_in_last_level_0__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[64]), .Z(
        buf_in_last_level_1__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[64]), .Z(
        buf_in_last_level_2__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_64__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[64]), .Z(
        buf_in_last_level_3__i_data_o_buf[64]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[65]), .Z(
        buf_in_last_level_0__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[65]), .Z(
        buf_in_last_level_1__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[65]), .Z(
        buf_in_last_level_2__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_65__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[65]), .Z(
        buf_in_last_level_3__i_data_o_buf[65]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[66]), .Z(
        buf_in_last_level_0__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[66]), .Z(
        buf_in_last_level_1__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[66]), .Z(
        buf_in_last_level_2__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_66__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[66]), .Z(
        buf_in_last_level_3__i_data_o_buf[66]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[67]), .Z(
        buf_in_last_level_0__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[67]), .Z(
        buf_in_last_level_1__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[67]), .Z(
        buf_in_last_level_2__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_67__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[67]), .Z(
        buf_in_last_level_3__i_data_o_buf[67]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[68]), .Z(
        buf_in_last_level_0__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[68]), .Z(
        buf_in_last_level_1__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[68]), .Z(
        buf_in_last_level_2__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_68__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[68]), .Z(
        buf_in_last_level_3__i_data_o_buf[68]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[69]), .Z(
        buf_in_last_level_0__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[69]), .Z(
        buf_in_last_level_1__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[69]), .Z(
        buf_in_last_level_2__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_69__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[69]), .Z(
        buf_in_last_level_3__i_data_o_buf[69]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[70]), .Z(
        buf_in_last_level_0__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[70]), .Z(
        buf_in_last_level_1__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[70]), .Z(
        buf_in_last_level_2__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_70__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[70]), .Z(
        buf_in_last_level_3__i_data_o_buf[70]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[71]), .Z(
        buf_in_last_level_0__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[71]), .Z(
        buf_in_last_level_1__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[71]), .Z(
        buf_in_last_level_2__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_71__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[71]), .Z(
        buf_in_last_level_3__i_data_o_buf[71]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[72]), .Z(
        buf_in_last_level_0__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[72]), .Z(
        buf_in_last_level_1__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[72]), .Z(
        buf_in_last_level_2__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_72__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[72]), .Z(
        buf_in_last_level_3__i_data_o_buf[72]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[73]), .Z(
        buf_in_last_level_0__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[73]), .Z(
        buf_in_last_level_1__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[73]), .Z(
        buf_in_last_level_2__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_73__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[73]), .Z(
        buf_in_last_level_3__i_data_o_buf[73]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[74]), .Z(
        buf_in_last_level_0__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[74]), .Z(
        buf_in_last_level_1__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[74]), .Z(
        buf_in_last_level_2__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_74__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[74]), .Z(
        buf_in_last_level_3__i_data_o_buf[74]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[75]), .Z(
        buf_in_last_level_0__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[75]), .Z(
        buf_in_last_level_1__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[75]), .Z(
        buf_in_last_level_2__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_75__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[75]), .Z(
        buf_in_last_level_3__i_data_o_buf[75]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[76]), .Z(
        buf_in_last_level_0__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[76]), .Z(
        buf_in_last_level_1__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[76]), .Z(
        buf_in_last_level_2__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_76__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[76]), .Z(
        buf_in_last_level_3__i_data_o_buf[76]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[77]), .Z(
        buf_in_last_level_0__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[77]), .Z(
        buf_in_last_level_1__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[77]), .Z(
        buf_in_last_level_2__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_77__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[77]), .Z(
        buf_in_last_level_3__i_data_o_buf[77]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[78]), .Z(
        buf_in_last_level_0__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[78]), .Z(
        buf_in_last_level_1__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[78]), .Z(
        buf_in_last_level_2__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_78__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[78]), .Z(
        buf_in_last_level_3__i_data_o_buf[78]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[79]), .Z(
        buf_in_last_level_0__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[79]), .Z(
        buf_in_last_level_1__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[79]), .Z(
        buf_in_last_level_2__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_79__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[79]), .Z(
        buf_in_last_level_3__i_data_o_buf[79]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[80]), .Z(
        buf_in_last_level_0__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[80]), .Z(
        buf_in_last_level_1__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[80]), .Z(
        buf_in_last_level_2__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_80__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[80]), .Z(
        buf_in_last_level_3__i_data_o_buf[80]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[81]), .Z(
        buf_in_last_level_0__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[81]), .Z(
        buf_in_last_level_1__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[81]), .Z(
        buf_in_last_level_2__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_81__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[81]), .Z(
        buf_in_last_level_3__i_data_o_buf[81]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[82]), .Z(
        buf_in_last_level_0__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[82]), .Z(
        buf_in_last_level_1__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[82]), .Z(
        buf_in_last_level_2__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_82__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[82]), .Z(
        buf_in_last_level_3__i_data_o_buf[82]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[83]), .Z(
        buf_in_last_level_0__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[83]), .Z(
        buf_in_last_level_1__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[83]), .Z(
        buf_in_last_level_2__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_83__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[83]), .Z(
        buf_in_last_level_3__i_data_o_buf[83]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[84]), .Z(
        buf_in_last_level_0__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[84]), .Z(
        buf_in_last_level_1__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[84]), .Z(
        buf_in_last_level_2__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_84__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[84]), .Z(
        buf_in_last_level_3__i_data_o_buf[84]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[85]), .Z(
        buf_in_last_level_0__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[85]), .Z(
        buf_in_last_level_1__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[85]), .Z(
        buf_in_last_level_2__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_85__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[85]), .Z(
        buf_in_last_level_3__i_data_o_buf[85]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[86]), .Z(
        buf_in_last_level_0__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[86]), .Z(
        buf_in_last_level_1__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[86]), .Z(
        buf_in_last_level_2__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_86__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[86]), .Z(
        buf_in_last_level_3__i_data_o_buf[86]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[87]), .Z(
        buf_in_last_level_0__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[87]), .Z(
        buf_in_last_level_1__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[87]), .Z(
        buf_in_last_level_2__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_87__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[87]), .Z(
        buf_in_last_level_3__i_data_o_buf[87]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[88]), .Z(
        buf_in_last_level_0__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[88]), .Z(
        buf_in_last_level_1__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[88]), .Z(
        buf_in_last_level_2__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_88__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[88]), .Z(
        buf_in_last_level_3__i_data_o_buf[88]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[89]), .Z(
        buf_in_last_level_0__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[89]), .Z(
        buf_in_last_level_1__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[89]), .Z(
        buf_in_last_level_2__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_89__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[89]), .Z(
        buf_in_last_level_3__i_data_o_buf[89]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[90]), .Z(
        buf_in_last_level_0__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[90]), .Z(
        buf_in_last_level_1__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[90]), .Z(
        buf_in_last_level_2__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_90__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[90]), .Z(
        buf_in_last_level_3__i_data_o_buf[90]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[91]), .Z(
        buf_in_last_level_0__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[91]), .Z(
        buf_in_last_level_1__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[91]), .Z(
        buf_in_last_level_2__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_91__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[91]), .Z(
        buf_in_last_level_3__i_data_o_buf[91]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[92]), .Z(
        buf_in_last_level_0__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[92]), .Z(
        buf_in_last_level_1__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[92]), .Z(
        buf_in_last_level_2__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_92__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[92]), .Z(
        buf_in_last_level_3__i_data_o_buf[92]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[93]), .Z(
        buf_in_last_level_0__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[93]), .Z(
        buf_in_last_level_1__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[93]), .Z(
        buf_in_last_level_2__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_93__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[93]), .Z(
        buf_in_last_level_3__i_data_o_buf[93]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[94]), .Z(
        buf_in_last_level_0__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[94]), .Z(
        buf_in_last_level_1__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[94]), .Z(
        buf_in_last_level_2__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_94__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[94]), .Z(
        buf_in_last_level_3__i_data_o_buf[94]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[95]), .Z(
        buf_in_last_level_0__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[95]), .Z(
        buf_in_last_level_1__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[95]), .Z(
        buf_in_last_level_2__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_95__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[95]), .Z(
        buf_in_last_level_3__i_data_o_buf[95]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[96]), .Z(
        buf_in_last_level_0__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[96]), .Z(
        buf_in_last_level_1__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[96]), .Z(
        buf_in_last_level_2__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_96__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[96]), .Z(
        buf_in_last_level_3__i_data_o_buf[96]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[97]), .Z(
        buf_in_last_level_0__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[97]), .Z(
        buf_in_last_level_1__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[97]), .Z(
        buf_in_last_level_2__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_97__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[97]), .Z(
        buf_in_last_level_3__i_data_o_buf[97]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[98]), .Z(
        buf_in_last_level_0__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[98]), .Z(
        buf_in_last_level_1__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[98]), .Z(
        buf_in_last_level_2__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_98__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[98]), .Z(
        buf_in_last_level_3__i_data_o_buf[98]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[99]), .Z(
        buf_in_last_level_0__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[99]), .Z(
        buf_in_last_level_1__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[99]), .Z(
        buf_in_last_level_2__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_99__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[99]), .Z(
        buf_in_last_level_3__i_data_o_buf[99]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[100]), .Z(
        buf_in_last_level_0__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[100]), .Z(
        buf_in_last_level_1__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[100]), .Z(
        buf_in_last_level_2__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_100__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[100]), .Z(
        buf_in_last_level_3__i_data_o_buf[100]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[101]), .Z(
        buf_in_last_level_0__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[101]), .Z(
        buf_in_last_level_1__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[101]), .Z(
        buf_in_last_level_2__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_101__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[101]), .Z(
        buf_in_last_level_3__i_data_o_buf[101]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[102]), .Z(
        buf_in_last_level_0__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[102]), .Z(
        buf_in_last_level_1__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[102]), .Z(
        buf_in_last_level_2__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_102__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[102]), .Z(
        buf_in_last_level_3__i_data_o_buf[102]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[103]), .Z(
        buf_in_last_level_0__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[103]), .Z(
        buf_in_last_level_1__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[103]), .Z(
        buf_in_last_level_2__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_103__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[103]), .Z(
        buf_in_last_level_3__i_data_o_buf[103]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[104]), .Z(
        buf_in_last_level_0__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[104]), .Z(
        buf_in_last_level_1__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[104]), .Z(
        buf_in_last_level_2__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_104__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[104]), .Z(
        buf_in_last_level_3__i_data_o_buf[104]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[105]), .Z(
        buf_in_last_level_0__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[105]), .Z(
        buf_in_last_level_1__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[105]), .Z(
        buf_in_last_level_2__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_105__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[105]), .Z(
        buf_in_last_level_3__i_data_o_buf[105]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[106]), .Z(
        buf_in_last_level_0__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[106]), .Z(
        buf_in_last_level_1__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[106]), .Z(
        buf_in_last_level_2__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_106__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[106]), .Z(
        buf_in_last_level_3__i_data_o_buf[106]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[107]), .Z(
        buf_in_last_level_0__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[107]), .Z(
        buf_in_last_level_1__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[107]), .Z(
        buf_in_last_level_2__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_107__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[107]), .Z(
        buf_in_last_level_3__i_data_o_buf[107]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[108]), .Z(
        buf_in_last_level_0__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[108]), .Z(
        buf_in_last_level_1__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[108]), .Z(
        buf_in_last_level_2__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_108__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[108]), .Z(
        buf_in_last_level_3__i_data_o_buf[108]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[109]), .Z(
        buf_in_last_level_0__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[109]), .Z(
        buf_in_last_level_1__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[109]), .Z(
        buf_in_last_level_2__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_109__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[109]), .Z(
        buf_in_last_level_3__i_data_o_buf[109]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[110]), .Z(
        buf_in_last_level_0__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[110]), .Z(
        buf_in_last_level_1__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[110]), .Z(
        buf_in_last_level_2__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_110__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[110]), .Z(
        buf_in_last_level_3__i_data_o_buf[110]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[111]), .Z(
        buf_in_last_level_0__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[111]), .Z(
        buf_in_last_level_1__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[111]), .Z(
        buf_in_last_level_2__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_111__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[111]), .Z(
        buf_in_last_level_3__i_data_o_buf[111]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[112]), .Z(
        buf_in_last_level_0__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[112]), .Z(
        buf_in_last_level_1__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[112]), .Z(
        buf_in_last_level_2__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_112__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[112]), .Z(
        buf_in_last_level_3__i_data_o_buf[112]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[113]), .Z(
        buf_in_last_level_0__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[113]), .Z(
        buf_in_last_level_1__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[113]), .Z(
        buf_in_last_level_2__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_113__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[113]), .Z(
        buf_in_last_level_3__i_data_o_buf[113]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[114]), .Z(
        buf_in_last_level_0__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[114]), .Z(
        buf_in_last_level_1__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[114]), .Z(
        buf_in_last_level_2__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_114__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[114]), .Z(
        buf_in_last_level_3__i_data_o_buf[114]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[115]), .Z(
        buf_in_last_level_0__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[115]), .Z(
        buf_in_last_level_1__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[115]), .Z(
        buf_in_last_level_2__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_115__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[115]), .Z(
        buf_in_last_level_3__i_data_o_buf[115]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[116]), .Z(
        buf_in_last_level_0__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[116]), .Z(
        buf_in_last_level_1__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[116]), .Z(
        buf_in_last_level_2__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_116__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[116]), .Z(
        buf_in_last_level_3__i_data_o_buf[116]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[117]), .Z(
        buf_in_last_level_0__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[117]), .Z(
        buf_in_last_level_1__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[117]), .Z(
        buf_in_last_level_2__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_117__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[117]), .Z(
        buf_in_last_level_3__i_data_o_buf[117]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[118]), .Z(
        buf_in_last_level_0__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[118]), .Z(
        buf_in_last_level_1__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[118]), .Z(
        buf_in_last_level_2__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_118__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[118]), .Z(
        buf_in_last_level_3__i_data_o_buf[118]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[119]), .Z(
        buf_in_last_level_0__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[119]), .Z(
        buf_in_last_level_1__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[119]), .Z(
        buf_in_last_level_2__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_119__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[119]), .Z(
        buf_in_last_level_3__i_data_o_buf[119]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[120]), .Z(
        buf_in_last_level_0__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[120]), .Z(
        buf_in_last_level_1__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[120]), .Z(
        buf_in_last_level_2__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_120__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[120]), .Z(
        buf_in_last_level_3__i_data_o_buf[120]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[121]), .Z(
        buf_in_last_level_0__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[121]), .Z(
        buf_in_last_level_1__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[121]), .Z(
        buf_in_last_level_2__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_121__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[121]), .Z(
        buf_in_last_level_3__i_data_o_buf[121]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[122]), .Z(
        buf_in_last_level_0__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[122]), .Z(
        buf_in_last_level_1__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[122]), .Z(
        buf_in_last_level_2__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_122__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[122]), .Z(
        buf_in_last_level_3__i_data_o_buf[122]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[123]), .Z(
        buf_in_last_level_0__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[123]), .Z(
        buf_in_last_level_1__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[123]), .Z(
        buf_in_last_level_2__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_123__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[123]), .Z(
        buf_in_last_level_3__i_data_o_buf[123]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[124]), .Z(
        buf_in_last_level_0__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[124]), .Z(
        buf_in_last_level_1__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[124]), .Z(
        buf_in_last_level_2__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_124__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[124]), .Z(
        buf_in_last_level_3__i_data_o_buf[124]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[125]), .Z(
        buf_in_last_level_0__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[125]), .Z(
        buf_in_last_level_1__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[125]), .Z(
        buf_in_last_level_2__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_125__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[125]), .Z(
        buf_in_last_level_3__i_data_o_buf[125]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[126]), .Z(
        buf_in_last_level_0__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[126]), .Z(
        buf_in_last_level_1__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[126]), .Z(
        buf_in_last_level_2__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_126__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[126]), .Z(
        buf_in_last_level_3__i_data_o_buf[126]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__UI_BUF_o_data_bus_first ( 
        .I(wire_tree_level_2__i_data_latch[127]), .Z(
        buf_in_last_level_0__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_0__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_0__i_data_o_buf[127]), .Z(
        buf_in_last_level_1__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_1__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_1__i_data_o_buf[127]), .Z(
        buf_in_last_level_2__i_data_o_buf[127]) );
  BUFFD0BWP30P140LVT UI_buf_in_last_level_assign_127__buf_levelS_2__UI_BUF_o_data_bus_stage_after ( 
        .I(buf_in_last_level_2__i_data_o_buf[127]), .Z(
        buf_in_last_level_3__i_data_o_buf[127]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_valid_latch_reg_0_ ( .D(N35), .CP(CLK), .Q(wire_tree_level_0__i_valid_latch_0_) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_31_ ( .D(N34), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_30_ ( .D(N33), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_29_ ( .D(N32), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_28_ ( .D(N31), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_27_ ( .D(N30), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_26_ ( .D(N29), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_25_ ( .D(N28), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_24_ ( .D(N27), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_23_ ( .D(N26), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_22_ ( .D(N25), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_21_ ( .D(N24), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_20_ ( .D(N23), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_19_ ( .D(N22), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_18_ ( .D(N21), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_17_ ( .D(N20), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_16_ ( .D(N19), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_15_ ( .D(N18), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_14_ ( .D(N17), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_13_ ( .D(N16), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_12_ ( .D(N15), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_11_ ( .D(N14), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_10_ ( .D(N13), .CP(CLK), .Q(wire_tree_level_0__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_9_ ( .D(N12), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_8_ ( .D(N11), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_7_ ( .D(N10), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_6_ ( .D(N9), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_5_ ( .D(N8), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_4_ ( .D(N7), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_3_ ( .D(N6), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_2_ ( .D(N5), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_1_ ( .D(N4), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_0__i_data_latch_reg_0_ ( .D(N3), .CP(CLK), 
        .Q(wire_tree_level_0__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_63_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_62_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_61_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_60_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_59_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_58_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_57_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_56_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_55_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_54_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_53_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_52_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_51_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_50_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_49_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_48_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_47_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_46_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_45_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_44_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_43_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_42_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_41_ ( .D(N77), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_40_ ( .D(N76), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_39_ ( .D(N75), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_38_ ( .D(N74), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_37_ ( .D(N73), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_36_ ( .D(N72), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_35_ ( .D(N71), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_34_ ( .D(N70), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_33_ ( .D(N69), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_32_ ( .D(N68), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_31_ ( .D(N99), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_30_ ( .D(N98), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_29_ ( .D(N97), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_28_ ( .D(N96), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_27_ ( .D(N95), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_26_ ( .D(N94), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_25_ ( .D(N93), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_24_ ( .D(N92), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_23_ ( .D(N91), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_22_ ( .D(N90), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_21_ ( .D(N89), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_20_ ( .D(N88), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_19_ ( .D(N87), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_18_ ( .D(N86), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_17_ ( .D(N85), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_16_ ( .D(N84), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_15_ ( .D(N83), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_14_ ( .D(N82), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_13_ ( .D(N81), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_12_ ( .D(N80), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_11_ ( .D(N79), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_10_ ( .D(N78), .CP(CLK), .Q(wire_tree_level_1__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_9_ ( .D(N77), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_8_ ( .D(N76), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_7_ ( .D(N75), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_6_ ( .D(N74), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_5_ ( .D(N73), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_4_ ( .D(N72), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_3_ ( .D(N71), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_2_ ( .D(N70), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_1_ ( .D(N69), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_data_latch_reg_0_ ( .D(N68), .CP(CLK), 
        .Q(wire_tree_level_1__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_1_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_1__i_valid_latch_reg_0_ ( .D(N101), .CP(
        CLK), .Q(wire_tree_level_1__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_63_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[63]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_62_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[62]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_61_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[61]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_60_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[60]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_59_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[59]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_58_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[58]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_57_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[57]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_56_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[56]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_55_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[55]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_54_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[54]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_53_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[53]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_52_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[52]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_51_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[51]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_50_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[50]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_49_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[49]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_48_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[48]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_47_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[47]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_46_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[46]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_45_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[45]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_44_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[44]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_43_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[43]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_42_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[42]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_41_ ( .D(N143), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[41]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_40_ ( .D(N142), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[40]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_39_ ( .D(N141), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[39]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_38_ ( .D(N140), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[38]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_37_ ( .D(N139), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[37]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_36_ ( .D(N138), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[36]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_35_ ( .D(N137), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[35]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_34_ ( .D(N136), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[34]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_33_ ( .D(N135), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[33]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_32_ ( .D(N134), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[32]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_31_ ( .D(N165), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[31]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_30_ ( .D(N164), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[30]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_29_ ( .D(N163), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[29]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_28_ ( .D(N162), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[28]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_27_ ( .D(N161), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[27]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_26_ ( .D(N160), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[26]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_25_ ( .D(N159), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[25]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_24_ ( .D(N158), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[24]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_23_ ( .D(N157), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[23]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_22_ ( .D(N156), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[22]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_21_ ( .D(N155), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[21]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_20_ ( .D(N154), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[20]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_19_ ( .D(N153), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[19]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_18_ ( .D(N152), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[18]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_17_ ( .D(N151), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[17]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_16_ ( .D(N150), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[16]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_15_ ( .D(N149), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[15]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_14_ ( .D(N148), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[14]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_13_ ( .D(N147), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[13]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_12_ ( .D(N146), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[12]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_11_ ( .D(N145), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[11]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_10_ ( .D(N144), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[10]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_9_ ( .D(N143), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[9]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_8_ ( .D(N142), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[8]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_7_ ( .D(N141), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[7]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_6_ ( .D(N140), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[6]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_5_ ( .D(N139), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[5]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_4_ ( .D(N138), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[4]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_3_ ( .D(N137), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_2_ ( .D(N136), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[2]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_1_ ( .D(N135), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_0_ ( .D(N134), .CP(CLK), .Q(wire_tree_level_2__i_data_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_1_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[1]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_0_ ( .D(N167), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[0]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_127_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[127]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_126_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[126]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_125_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[125]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_124_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[124]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_123_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[123]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_122_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[122]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_121_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[121]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_120_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[120]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_119_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[119]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_118_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[118]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_117_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[117]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_116_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[116]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_115_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[115]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_114_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[114]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_113_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[113]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_112_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[112]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_111_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[111]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_110_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[110]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_109_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[109]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_108_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[108]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_107_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[107]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_106_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[106]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_105_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[105]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_104_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[104]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_103_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[103]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_102_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[102]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_101_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[101]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_100_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[100]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_99_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[99]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_98_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[98]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_97_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[97]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_96_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[96]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_95_ ( .D(N231), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[95]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_94_ ( .D(N230), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[94]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_93_ ( .D(N229), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[93]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_92_ ( .D(N228), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[92]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_91_ ( .D(N227), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[91]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_90_ ( .D(N226), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[90]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_89_ ( .D(N225), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[89]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_88_ ( .D(N224), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[88]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_87_ ( .D(N223), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[87]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_86_ ( .D(N222), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[86]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_85_ ( .D(N221), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[85]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_84_ ( .D(N220), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[84]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_83_ ( .D(N219), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[83]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_82_ ( .D(N218), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[82]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_81_ ( .D(N217), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[81]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_80_ ( .D(N216), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[80]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_79_ ( .D(N215), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[79]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_78_ ( .D(N214), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[78]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_77_ ( .D(N213), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[77]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_76_ ( .D(N212), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[76]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_75_ ( .D(N211), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[75]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_74_ ( .D(N210), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[74]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_73_ ( .D(N209), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[73]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_72_ ( .D(N208), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[72]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_71_ ( .D(N207), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[71]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_70_ ( .D(N206), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[70]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_69_ ( .D(N205), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[69]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_68_ ( .D(N204), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[68]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_67_ ( .D(N203), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[67]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_66_ ( .D(N202), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[66]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_65_ ( .D(N201), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[65]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_data_latch_reg_64_ ( .D(N200), .CP(
        CLK), .Q(wire_tree_level_2__i_data_latch[64]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_3_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[3]) );
  DFQD1BWP30P140LVT wire_tree_level_2__i_valid_latch_reg_2_ ( .D(N233), .CP(
        CLK), .Q(wire_tree_level_2__i_valid_latch[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N297), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N296), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N295), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N294), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N293), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N292), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N291), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N290), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N289), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N288), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N287), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N286), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N285), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N284), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N283), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N282), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N281), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N280), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N279), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N278), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N277), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N276), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N275), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N274), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N273), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N272), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N271), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N270), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N269), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N268), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N267), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N266), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_1_ ( .D(N299), .CP(CLK), .Q(o_valid[1]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N299), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N363), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N362), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N361), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N360), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N359), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N358), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N357), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N356), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N355), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N354), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N353), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N352), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N351), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N350), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N349), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N348), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N347), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N346), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N345), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_3_ ( .D(N365), .CP(CLK), .Q(o_valid[3]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_2_ ( .D(N365), .CP(CLK), .Q(o_valid[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(N429), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(N428), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(N427), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(N426), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(N425), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(N424), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(N423), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(N422), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(N421), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(N420), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N419), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N418), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N417), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N416), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N415), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N414), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N413), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N412), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N411), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N410), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N409), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N408), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N407), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N406), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N405), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N404), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N403), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N402), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N401), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_5_ ( .D(N431), .CP(CLK), .Q(o_valid[5]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_4_ ( .D(N431), .CP(CLK), .Q(o_valid[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N495), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N494), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N493), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N492), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N491), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N490), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N489), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N488), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N487), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N486), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N485), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N484), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N483), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N482), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N481), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N480), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N479), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N478), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N477), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N476), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N475), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N474), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N473), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N472), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N471), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N470), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N469), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N468), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N467), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N466), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N465), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N464), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_7_ ( .D(N497), .CP(CLK), .Q(o_valid[7]) );
  DFQD1BWP30P140LVT o_valid_reg_reg_6_ ( .D(N497), .CP(CLK), .Q(o_valid[6]) );
  CKAN2D1BWP30P140LVT U3 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[96]), 
        .Z(N464) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[6]), 
        .Z(N272) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[3]), 
        .Z(N497) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[97]), 
        .Z(N465) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[98]), 
        .Z(N466) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[99]), 
        .Z(N467) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[100]), .Z(N468) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[101]), .Z(N469) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[102]), .Z(N470) );
  CKAN2D1BWP30P140LVT U12 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[103]), .Z(N471) );
  CKAN2D1BWP30P140LVT U13 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[104]), .Z(N472) );
  CKAN2D1BWP30P140LVT U14 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[105]), .Z(N473) );
  CKAN2D1BWP30P140LVT U15 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[106]), .Z(N474) );
  CKAN2D1BWP30P140LVT U16 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[107]), .Z(N475) );
  CKAN2D1BWP30P140LVT U17 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[108]), .Z(N476) );
  CKAN2D1BWP30P140LVT U18 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[109]), .Z(N477) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[110]), .Z(N478) );
  CKAN2D1BWP30P140LVT U20 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[111]), .Z(N479) );
  CKAN2D1BWP30P140LVT U21 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[112]), .Z(N480) );
  CKAN2D1BWP30P140LVT U22 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[113]), .Z(N481) );
  CKAN2D1BWP30P140LVT U23 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[114]), .Z(N482) );
  CKAN2D1BWP30P140LVT U24 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[115]), .Z(N483) );
  CKAN2D1BWP30P140LVT U25 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[116]), .Z(N484) );
  CKAN2D1BWP30P140LVT U26 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[117]), .Z(N485) );
  CKAN2D1BWP30P140LVT U27 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[118]), .Z(N486) );
  CKAN2D1BWP30P140LVT U28 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[82]), .Z(N416) );
  CKAN2D1BWP30P140LVT U29 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[86]), .Z(N420) );
  CKAN2D1BWP30P140LVT U30 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[61]), .Z(N361) );
  CKAN2D1BWP30P140LVT U31 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[63]), .Z(N363) );
  CKAN2D1BWP30P140LVT U32 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[2]), 
        .Z(N268) );
  CKAN2D1BWP30P140LVT U33 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[44]), 
        .Z(N212) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[47]), 
        .Z(N215) );
  CKAN2D1BWP30P140LVT U35 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[51]), 
        .Z(N219) );
  CKAN2D1BWP30P140LVT U36 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[58]), 
        .Z(N226) );
  CKAN2D1BWP30P140LVT U37 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[62]), 
        .Z(N230) );
  CKAN2D1BWP30P140LVT U38 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[1]), 
        .Z(N135) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[2]), 
        .Z(N136) );
  CKAN2D1BWP30P140LVT U40 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[3]), 
        .Z(N137) );
  CKAN2D1BWP30P140LVT U41 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[4]), 
        .Z(N138) );
  CKAN2D1BWP30P140LVT U42 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[5]), 
        .Z(N139) );
  CKAN2D1BWP30P140LVT U43 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[6]), 
        .Z(N140) );
  CKAN2D1BWP30P140LVT U44 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[7]), 
        .Z(N141) );
  CKAN2D1BWP30P140LVT U45 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[8]), 
        .Z(N142) );
  CKAN2D1BWP30P140LVT U46 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[9]), 
        .Z(N143) );
  CKAN2D1BWP30P140LVT U47 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[10]), 
        .Z(N144) );
  CKAN2D1BWP30P140LVT U48 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[11]), 
        .Z(N145) );
  CKAN2D1BWP30P140LVT U49 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[12]), 
        .Z(N146) );
  CKAN2D1BWP30P140LVT U50 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[13]), 
        .Z(N147) );
  CKAN2D1BWP30P140LVT U51 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[14]), 
        .Z(N148) );
  CKAN2D1BWP30P140LVT U52 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[15]), 
        .Z(N149) );
  CKAN2D1BWP30P140LVT U53 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[16]), 
        .Z(N150) );
  CKAN2D1BWP30P140LVT U54 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[17]), 
        .Z(N151) );
  CKAN2D1BWP30P140LVT U55 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[18]), 
        .Z(N152) );
  CKAN2D1BWP30P140LVT U56 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[19]), 
        .Z(N153) );
  CKAN2D1BWP30P140LVT U57 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[20]), 
        .Z(N154) );
  CKAN2D1BWP30P140LVT U58 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[21]), 
        .Z(N155) );
  CKAN2D1BWP30P140LVT U59 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[22]), 
        .Z(N156) );
  CKAN2D1BWP30P140LVT U60 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[23]), 
        .Z(N157) );
  CKAN2D1BWP30P140LVT U61 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[24]), 
        .Z(N158) );
  CKAN2D1BWP30P140LVT U62 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[25]), 
        .Z(N159) );
  CKAN2D1BWP30P140LVT U63 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[26]), 
        .Z(N160) );
  CKAN2D1BWP30P140LVT U64 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[27]), 
        .Z(N161) );
  CKAN2D1BWP30P140LVT U65 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[28]), 
        .Z(N162) );
  CKAN2D1BWP30P140LVT U66 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[29]), 
        .Z(N163) );
  CKAN2D1BWP30P140LVT U67 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[30]), 
        .Z(N164) );
  CKAN2D1BWP30P140LVT U68 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[31]), 
        .Z(N165) );
  CKAN2D1BWP30P140LVT U69 ( .A1(n1), .A2(wire_tree_level_0__i_valid_latch_0_), 
        .Z(N101) );
  CKAN2D1BWP30P140LVT U70 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[0]), 
        .Z(N68) );
  CKAN2D1BWP30P140LVT U71 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[1]), 
        .Z(N69) );
  CKAN2D1BWP30P140LVT U72 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[2]), 
        .Z(N70) );
  CKAN2D1BWP30P140LVT U73 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[3]), 
        .Z(N71) );
  CKAN2D1BWP30P140LVT U74 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[4]), 
        .Z(N72) );
  CKAN2D1BWP30P140LVT U75 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[5]), 
        .Z(N73) );
  CKAN2D1BWP30P140LVT U76 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[6]), 
        .Z(N74) );
  CKAN2D1BWP30P140LVT U77 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[7]), 
        .Z(N75) );
  CKAN2D1BWP30P140LVT U78 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[8]), 
        .Z(N76) );
  CKAN2D1BWP30P140LVT U79 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[9]), 
        .Z(N77) );
  CKAN2D1BWP30P140LVT U80 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[10]), 
        .Z(N78) );
  CKAN2D1BWP30P140LVT U81 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[11]), 
        .Z(N79) );
  CKAN2D1BWP30P140LVT U82 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[12]), 
        .Z(N80) );
  CKAN2D1BWP30P140LVT U83 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[13]), 
        .Z(N81) );
  CKAN2D1BWP30P140LVT U84 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[14]), 
        .Z(N82) );
  CKAN2D1BWP30P140LVT U85 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[15]), 
        .Z(N83) );
  CKAN2D1BWP30P140LVT U86 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[16]), 
        .Z(N84) );
  CKAN2D1BWP30P140LVT U87 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[17]), 
        .Z(N85) );
  CKAN2D1BWP30P140LVT U88 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[18]), 
        .Z(N86) );
  CKAN2D1BWP30P140LVT U89 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[19]), 
        .Z(N87) );
  CKAN2D1BWP30P140LVT U90 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[20]), 
        .Z(N88) );
  CKAN2D1BWP30P140LVT U91 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[21]), 
        .Z(N89) );
  CKAN2D1BWP30P140LVT U92 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[22]), 
        .Z(N90) );
  CKAN2D1BWP30P140LVT U93 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[23]), 
        .Z(N91) );
  CKAN2D1BWP30P140LVT U94 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[24]), 
        .Z(N92) );
  CKAN2D1BWP30P140LVT U95 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[25]), 
        .Z(N93) );
  CKAN2D1BWP30P140LVT U96 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[26]), 
        .Z(N94) );
  CKAN2D1BWP30P140LVT U97 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[27]), 
        .Z(N95) );
  CKAN2D1BWP30P140LVT U98 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[28]), 
        .Z(N96) );
  CKAN2D1BWP30P140LVT U99 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[29]), 
        .Z(N97) );
  CKAN2D1BWP30P140LVT U100 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[30]), 
        .Z(N98) );
  CKAN2D1BWP30P140LVT U101 ( .A1(n1), .A2(wire_tree_level_0__i_data_latch[31]), 
        .Z(N99) );
  CKAN2D1BWP30P140LVT U102 ( .A1(n1), .A2(i_data_bus[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U103 ( .A1(n1), .A2(i_data_bus[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U104 ( .A1(n1), .A2(i_data_bus[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U105 ( .A1(n1), .A2(i_data_bus[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U106 ( .A1(n1), .A2(i_data_bus[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U107 ( .A1(n1), .A2(i_data_bus[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U108 ( .A1(n1), .A2(i_data_bus[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U109 ( .A1(n1), .A2(i_data_bus[7]), .Z(N10) );
  CKAN2D1BWP30P140LVT U110 ( .A1(n1), .A2(i_data_bus[8]), .Z(N11) );
  CKAN2D1BWP30P140LVT U111 ( .A1(n1), .A2(i_data_bus[9]), .Z(N12) );
  CKAN2D1BWP30P140LVT U112 ( .A1(n1), .A2(i_data_bus[10]), .Z(N13) );
  CKAN2D1BWP30P140LVT U113 ( .A1(n1), .A2(i_data_bus[11]), .Z(N14) );
  CKAN2D1BWP30P140LVT U114 ( .A1(n1), .A2(i_data_bus[12]), .Z(N15) );
  CKAN2D1BWP30P140LVT U115 ( .A1(n1), .A2(i_data_bus[13]), .Z(N16) );
  CKAN2D1BWP30P140LVT U116 ( .A1(n1), .A2(i_data_bus[14]), .Z(N17) );
  CKAN2D1BWP30P140LVT U117 ( .A1(n1), .A2(i_data_bus[15]), .Z(N18) );
  CKAN2D1BWP30P140LVT U118 ( .A1(n1), .A2(i_data_bus[16]), .Z(N19) );
  CKAN2D1BWP30P140LVT U119 ( .A1(n1), .A2(i_data_bus[17]), .Z(N20) );
  CKAN2D1BWP30P140LVT U120 ( .A1(n1), .A2(i_data_bus[18]), .Z(N21) );
  CKAN2D1BWP30P140LVT U121 ( .A1(n1), .A2(i_data_bus[19]), .Z(N22) );
  CKAN2D1BWP30P140LVT U122 ( .A1(n1), .A2(i_data_bus[20]), .Z(N23) );
  CKAN2D1BWP30P140LVT U123 ( .A1(n1), .A2(i_data_bus[21]), .Z(N24) );
  CKAN2D1BWP30P140LVT U124 ( .A1(n1), .A2(i_data_bus[22]), .Z(N25) );
  CKAN2D1BWP30P140LVT U125 ( .A1(n1), .A2(i_data_bus[23]), .Z(N26) );
  CKAN2D1BWP30P140LVT U126 ( .A1(n1), .A2(i_data_bus[24]), .Z(N27) );
  CKAN2D1BWP30P140LVT U127 ( .A1(n1), .A2(i_data_bus[25]), .Z(N28) );
  CKAN2D1BWP30P140LVT U128 ( .A1(n1), .A2(i_data_bus[26]), .Z(N29) );
  CKAN2D1BWP30P140LVT U129 ( .A1(n1), .A2(i_data_bus[27]), .Z(N30) );
  CKAN2D1BWP30P140LVT U130 ( .A1(n1), .A2(i_data_bus[28]), .Z(N31) );
  CKAN2D1BWP30P140LVT U131 ( .A1(n1), .A2(i_data_bus[29]), .Z(N32) );
  CKAN2D1BWP30P140LVT U132 ( .A1(n1), .A2(i_data_bus[30]), .Z(N33) );
  CKAN2D1BWP30P140LVT U133 ( .A1(n1), .A2(i_data_bus[31]), .Z(N34) );
  CKAN2D1BWP30P140LVT U134 ( .A1(n1), .A2(i_valid[0]), .Z(N35) );
  INR2D2BWP30P140LVT U135 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U136 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[0]), 
        .Z(N134) );
  CKAN2D1BWP30P140LVT U137 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[0]), 
        .Z(N167) );
  CKAN2D1BWP30P140LVT U138 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[63]), 
        .Z(N231) );
  CKAN2D1BWP30P140LVT U139 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[61]), 
        .Z(N229) );
  CKAN2D1BWP30P140LVT U140 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[60]), 
        .Z(N228) );
  CKAN2D1BWP30P140LVT U141 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[59]), 
        .Z(N227) );
  CKAN2D1BWP30P140LVT U142 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[57]), 
        .Z(N225) );
  CKAN2D1BWP30P140LVT U143 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[56]), 
        .Z(N224) );
  CKAN2D1BWP30P140LVT U144 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[55]), 
        .Z(N223) );
  CKAN2D1BWP30P140LVT U145 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[54]), 
        .Z(N222) );
  CKAN2D1BWP30P140LVT U146 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[53]), 
        .Z(N221) );
  CKAN2D1BWP30P140LVT U147 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[52]), 
        .Z(N220) );
  CKAN2D1BWP30P140LVT U148 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[50]), 
        .Z(N218) );
  CKAN2D1BWP30P140LVT U149 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[49]), 
        .Z(N217) );
  CKAN2D1BWP30P140LVT U150 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[48]), 
        .Z(N216) );
  CKAN2D1BWP30P140LVT U151 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[46]), 
        .Z(N214) );
  CKAN2D1BWP30P140LVT U152 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[45]), 
        .Z(N213) );
  CKAN2D1BWP30P140LVT U153 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[43]), 
        .Z(N211) );
  CKAN2D1BWP30P140LVT U154 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[42]), 
        .Z(N210) );
  CKAN2D1BWP30P140LVT U155 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[41]), 
        .Z(N209) );
  CKAN2D1BWP30P140LVT U156 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[40]), 
        .Z(N208) );
  CKAN2D1BWP30P140LVT U157 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[39]), 
        .Z(N207) );
  CKAN2D1BWP30P140LVT U158 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[38]), 
        .Z(N206) );
  CKAN2D1BWP30P140LVT U159 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[37]), 
        .Z(N205) );
  CKAN2D1BWP30P140LVT U160 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[36]), 
        .Z(N204) );
  CKAN2D1BWP30P140LVT U161 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[35]), 
        .Z(N203) );
  CKAN2D1BWP30P140LVT U162 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[34]), 
        .Z(N202) );
  CKAN2D1BWP30P140LVT U163 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[33]), 
        .Z(N201) );
  CKAN2D1BWP30P140LVT U164 ( .A1(n1), .A2(wire_tree_level_1__i_data_latch[32]), 
        .Z(N200) );
  CKAN2D1BWP30P140LVT U165 ( .A1(n1), .A2(wire_tree_level_1__i_valid_latch[1]), 
        .Z(N233) );
  CKAN2D1BWP30P140LVT U166 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[0]), 
        .Z(N299) );
  CKAN2D1BWP30P140LVT U167 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[2]), 
        .Z(N431) );
  CKAN2D1BWP30P140LVT U168 ( .A1(n1), .A2(wire_tree_level_2__i_valid_latch[1]), 
        .Z(N365) );
  CKAN2D1BWP30P140LVT U169 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[31]), .Z(N297) );
  CKAN2D1BWP30P140LVT U170 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[29]), .Z(N295) );
  CKAN2D1BWP30P140LVT U171 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[28]), .Z(N294) );
  CKAN2D1BWP30P140LVT U172 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[27]), .Z(N293) );
  CKAN2D1BWP30P140LVT U173 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[26]), .Z(N292) );
  CKAN2D1BWP30P140LVT U174 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[25]), .Z(N291) );
  CKAN2D1BWP30P140LVT U175 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[24]), .Z(N290) );
  CKAN2D1BWP30P140LVT U176 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[23]), .Z(N289) );
  CKAN2D1BWP30P140LVT U177 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[22]), .Z(N288) );
  CKAN2D1BWP30P140LVT U178 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[21]), .Z(N287) );
  CKAN2D1BWP30P140LVT U179 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[20]), .Z(N286) );
  CKAN2D1BWP30P140LVT U180 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[30]), .Z(N296) );
  CKAN2D1BWP30P140LVT U181 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[17]), .Z(N283) );
  CKAN2D1BWP30P140LVT U182 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[16]), .Z(N282) );
  CKAN2D1BWP30P140LVT U183 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[15]), .Z(N281) );
  CKAN2D1BWP30P140LVT U184 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[14]), .Z(N280) );
  CKAN2D1BWP30P140LVT U185 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[13]), .Z(N279) );
  CKAN2D1BWP30P140LVT U186 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[12]), .Z(N278) );
  CKAN2D1BWP30P140LVT U187 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[11]), .Z(N277) );
  CKAN2D1BWP30P140LVT U188 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[10]), .Z(N276) );
  CKAN2D1BWP30P140LVT U189 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[9]), .Z(N275) );
  CKAN2D1BWP30P140LVT U190 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[8]), .Z(N274) );
  CKAN2D1BWP30P140LVT U191 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[7]), .Z(N273) );
  CKAN2D1BWP30P140LVT U192 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[4]), .Z(N270) );
  CKAN2D1BWP30P140LVT U193 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[3]), .Z(N269) );
  CKAN2D1BWP30P140LVT U194 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[1]), .Z(N267) );
  CKAN2D1BWP30P140LVT U195 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[0]), .Z(N266) );
  CKAN2D1BWP30P140LVT U196 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[18]), .Z(N284) );
  CKAN2D1BWP30P140LVT U197 ( .A1(n1), .A2(buf_in_last_level_3__i_data_o_buf[5]), .Z(N271) );
  CKAN2D1BWP30P140LVT U198 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[19]), .Z(N285) );
  CKAN2D1BWP30P140LVT U199 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[62]), .Z(N362) );
  CKAN2D1BWP30P140LVT U200 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[60]), .Z(N360) );
  CKAN2D1BWP30P140LVT U201 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[59]), .Z(N359) );
  CKAN2D1BWP30P140LVT U202 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[58]), .Z(N358) );
  CKAN2D1BWP30P140LVT U203 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[57]), .Z(N357) );
  CKAN2D1BWP30P140LVT U204 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[56]), .Z(N356) );
  CKAN2D1BWP30P140LVT U205 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[55]), .Z(N355) );
  CKAN2D1BWP30P140LVT U206 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[54]), .Z(N354) );
  CKAN2D1BWP30P140LVT U207 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[53]), .Z(N353) );
  CKAN2D1BWP30P140LVT U208 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[52]), .Z(N352) );
  CKAN2D1BWP30P140LVT U209 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[51]), .Z(N351) );
  CKAN2D1BWP30P140LVT U210 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[50]), .Z(N350) );
  CKAN2D1BWP30P140LVT U211 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[49]), .Z(N349) );
  CKAN2D1BWP30P140LVT U212 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[48]), .Z(N348) );
  CKAN2D1BWP30P140LVT U213 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[47]), .Z(N347) );
  CKAN2D1BWP30P140LVT U214 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[46]), .Z(N346) );
  CKAN2D1BWP30P140LVT U215 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[45]), .Z(N345) );
  CKAN2D1BWP30P140LVT U216 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[44]), .Z(N344) );
  CKAN2D1BWP30P140LVT U217 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[43]), .Z(N343) );
  CKAN2D1BWP30P140LVT U218 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[42]), .Z(N342) );
  CKAN2D1BWP30P140LVT U219 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[41]), .Z(N341) );
  CKAN2D1BWP30P140LVT U220 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[40]), .Z(N340) );
  CKAN2D1BWP30P140LVT U221 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[39]), .Z(N339) );
  CKAN2D1BWP30P140LVT U222 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[38]), .Z(N338) );
  CKAN2D1BWP30P140LVT U223 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[37]), .Z(N337) );
  CKAN2D1BWP30P140LVT U224 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[124]), .Z(N492) );
  CKAN2D1BWP30P140LVT U225 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[125]), .Z(N493) );
  CKAN2D1BWP30P140LVT U226 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[126]), .Z(N494) );
  CKAN2D1BWP30P140LVT U227 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[127]), .Z(N495) );
  CKAN2D1BWP30P140LVT U228 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[119]), .Z(N487) );
  CKAN2D1BWP30P140LVT U229 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[120]), .Z(N488) );
  CKAN2D1BWP30P140LVT U230 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[121]), .Z(N489) );
  CKAN2D1BWP30P140LVT U231 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[122]), .Z(N490) );
  CKAN2D1BWP30P140LVT U232 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[123]), .Z(N491) );
  CKAN2D1BWP30P140LVT U233 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[32]), .Z(N332) );
  CKAN2D1BWP30P140LVT U234 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[33]), .Z(N333) );
  CKAN2D1BWP30P140LVT U235 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[34]), .Z(N334) );
  CKAN2D1BWP30P140LVT U236 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[35]), .Z(N335) );
  CKAN2D1BWP30P140LVT U237 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[36]), .Z(N336) );
  CKAN2D1BWP30P140LVT U238 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[64]), .Z(N398) );
  CKAN2D1BWP30P140LVT U239 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[65]), .Z(N399) );
  CKAN2D1BWP30P140LVT U240 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[66]), .Z(N400) );
  CKAN2D1BWP30P140LVT U241 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[67]), .Z(N401) );
  CKAN2D1BWP30P140LVT U242 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[68]), .Z(N402) );
  CKAN2D1BWP30P140LVT U243 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[69]), .Z(N403) );
  CKAN2D1BWP30P140LVT U244 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[70]), .Z(N404) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[72]), .Z(N406) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[73]), .Z(N407) );
  CKAN2D1BWP30P140LVT U247 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[74]), .Z(N408) );
  CKAN2D1BWP30P140LVT U248 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[75]), .Z(N409) );
  CKAN2D1BWP30P140LVT U249 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[76]), .Z(N410) );
  CKAN2D1BWP30P140LVT U250 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[77]), .Z(N411) );
  CKAN2D1BWP30P140LVT U251 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[78]), .Z(N412) );
  CKAN2D1BWP30P140LVT U252 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[79]), .Z(N413) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[80]), .Z(N414) );
  CKAN2D1BWP30P140LVT U254 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[81]), .Z(N415) );
  CKAN2D1BWP30P140LVT U255 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[83]), .Z(N417) );
  CKAN2D1BWP30P140LVT U256 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[84]), .Z(N418) );
  CKAN2D1BWP30P140LVT U257 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[85]), .Z(N419) );
  CKAN2D1BWP30P140LVT U258 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[87]), .Z(N421) );
  CKAN2D1BWP30P140LVT U259 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[88]), .Z(N422) );
  CKAN2D1BWP30P140LVT U260 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[89]), .Z(N423) );
  CKAN2D1BWP30P140LVT U261 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[90]), .Z(N424) );
  CKAN2D1BWP30P140LVT U262 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[91]), .Z(N425) );
  CKAN2D1BWP30P140LVT U263 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[92]), .Z(N426) );
  CKAN2D1BWP30P140LVT U264 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[93]), .Z(N427) );
  CKAN2D1BWP30P140LVT U265 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[95]), .Z(N429) );
  CKAN2D1BWP30P140LVT U266 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[94]), .Z(N428) );
  CKAN2D1BWP30P140LVT U267 ( .A1(n1), .A2(
        buf_in_last_level_3__i_data_o_buf[71]), .Z(N405) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule


module crossbar_one_hot_seq ( CLK, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [63:0] i_cmd;
  input CLK, rst, i_en;
  wire   n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528;
  wire   [63:0] o_inner_cmd_wire;
  wire   [255:0] bottom_half_0__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_0__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_1__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_1__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_2__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_2__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_3__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_3__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_4__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_4__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_5__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_5__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_6__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_6__inner_valid_i_mux_tree_wire;
  wire   [255:0] bottom_half_7__inner_data_i_mux_tree_wire;
  wire   [7:0] bottom_half_7__inner_valid_i_mux_tree_wire;

  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 top_half_0__wire_pipeline ( 
        .CLK(CLK), .rst(rst), .i_valid(i_valid[0]), .i_data_bus(
        i_data_bus[31:0]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[0], 
        bottom_half_6__inner_valid_i_mux_tree_wire[0], 
        bottom_half_5__inner_valid_i_mux_tree_wire[0], 
        bottom_half_4__inner_valid_i_mux_tree_wire[0], 
        bottom_half_3__inner_valid_i_mux_tree_wire[0], 
        bottom_half_2__inner_valid_i_mux_tree_wire[0], 
        bottom_half_1__inner_valid_i_mux_tree_wire[0], 
        bottom_half_0__inner_valid_i_mux_tree_wire[0]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_6__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_5__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_4__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_3__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_2__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_1__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_0__inner_data_i_mux_tree_wire[31:0]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 top_half_1__wire_pipeline ( 
        .CLK(CLK), .rst(rst), .i_valid(i_valid[1]), .i_data_bus(
        i_data_bus[63:32]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[1], 
        bottom_half_6__inner_valid_i_mux_tree_wire[1], 
        bottom_half_5__inner_valid_i_mux_tree_wire[1], 
        bottom_half_4__inner_valid_i_mux_tree_wire[1], 
        bottom_half_3__inner_valid_i_mux_tree_wire[1], 
        bottom_half_2__inner_valid_i_mux_tree_wire[1], 
        bottom_half_1__inner_valid_i_mux_tree_wire[1], 
        bottom_half_0__inner_valid_i_mux_tree_wire[1]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_6__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_5__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_4__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_3__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_2__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_1__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_0__inner_data_i_mux_tree_wire[63:32]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 top_half_2__wire_pipeline ( 
        .CLK(CLK), .rst(rst), .i_valid(i_valid[2]), .i_data_bus(
        i_data_bus[95:64]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[2], 
        bottom_half_6__inner_valid_i_mux_tree_wire[2], 
        bottom_half_5__inner_valid_i_mux_tree_wire[2], 
        bottom_half_4__inner_valid_i_mux_tree_wire[2], 
        bottom_half_3__inner_valid_i_mux_tree_wire[2], 
        bottom_half_2__inner_valid_i_mux_tree_wire[2], 
        bottom_half_1__inner_valid_i_mux_tree_wire[2], 
        bottom_half_0__inner_valid_i_mux_tree_wire[2]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_6__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_5__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_4__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_3__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_2__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_1__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_0__inner_data_i_mux_tree_wire[95:64]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 top_half_3__wire_pipeline ( 
        .CLK(CLK), .rst(rst), .i_valid(i_valid[3]), .i_data_bus(
        i_data_bus[127:96]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[3], 
        bottom_half_6__inner_valid_i_mux_tree_wire[3], 
        bottom_half_5__inner_valid_i_mux_tree_wire[3], 
        bottom_half_4__inner_valid_i_mux_tree_wire[3], 
        bottom_half_3__inner_valid_i_mux_tree_wire[3], 
        bottom_half_2__inner_valid_i_mux_tree_wire[3], 
        bottom_half_1__inner_valid_i_mux_tree_wire[3], 
        bottom_half_0__inner_valid_i_mux_tree_wire[3]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_6__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_5__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_4__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_3__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_2__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_1__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_0__inner_data_i_mux_tree_wire[127:96]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 top_half_4__wire_pipeline ( 
        .CLK(CLK), .rst(rst), .i_valid(i_valid[4]), .i_data_bus(
        i_data_bus[159:128]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[4], 
        bottom_half_6__inner_valid_i_mux_tree_wire[4], 
        bottom_half_5__inner_valid_i_mux_tree_wire[4], 
        bottom_half_4__inner_valid_i_mux_tree_wire[4], 
        bottom_half_3__inner_valid_i_mux_tree_wire[4], 
        bottom_half_2__inner_valid_i_mux_tree_wire[4], 
        bottom_half_1__inner_valid_i_mux_tree_wire[4], 
        bottom_half_0__inner_valid_i_mux_tree_wire[4]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_6__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_5__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_4__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_3__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_2__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_1__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_0__inner_data_i_mux_tree_wire[159:128]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 top_half_5__wire_pipeline ( 
        .CLK(CLK), .rst(rst), .i_valid(i_valid[5]), .i_data_bus(
        i_data_bus[191:160]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[5], 
        bottom_half_6__inner_valid_i_mux_tree_wire[5], 
        bottom_half_5__inner_valid_i_mux_tree_wire[5], 
        bottom_half_4__inner_valid_i_mux_tree_wire[5], 
        bottom_half_3__inner_valid_i_mux_tree_wire[5], 
        bottom_half_2__inner_valid_i_mux_tree_wire[5], 
        bottom_half_1__inner_valid_i_mux_tree_wire[5], 
        bottom_half_0__inner_valid_i_mux_tree_wire[5]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_6__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_5__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_4__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_3__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_2__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_1__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_0__inner_data_i_mux_tree_wire[191:160]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 top_half_6__wire_pipeline ( 
        .CLK(CLK), .rst(rst), .i_valid(i_valid[6]), .i_data_bus(
        i_data_bus[223:192]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[6], 
        bottom_half_6__inner_valid_i_mux_tree_wire[6], 
        bottom_half_5__inner_valid_i_mux_tree_wire[6], 
        bottom_half_4__inner_valid_i_mux_tree_wire[6], 
        bottom_half_3__inner_valid_i_mux_tree_wire[6], 
        bottom_half_2__inner_valid_i_mux_tree_wire[6], 
        bottom_half_1__inner_valid_i_mux_tree_wire[6], 
        bottom_half_0__inner_valid_i_mux_tree_wire[6]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_6__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_5__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_4__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_3__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_2__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_1__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_0__inner_data_i_mux_tree_wire[223:192]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 top_half_7__wire_pipeline ( 
        .CLK(CLK), .rst(rst), .i_valid(i_valid[7]), .i_data_bus(
        i_data_bus[255:224]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[7], 
        bottom_half_6__inner_valid_i_mux_tree_wire[7], 
        bottom_half_5__inner_valid_i_mux_tree_wire[7], 
        bottom_half_4__inner_valid_i_mux_tree_wire[7], 
        bottom_half_3__inner_valid_i_mux_tree_wire[7], 
        bottom_half_2__inner_valid_i_mux_tree_wire[7], 
        bottom_half_1__inner_valid_i_mux_tree_wire[7], 
        bottom_half_0__inner_valid_i_mux_tree_wire[7]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_6__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_5__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_4__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_3__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_2__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_1__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_0__inner_data_i_mux_tree_wire[255:224]}), .i_en(i_en) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 i_cmd_id_0__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[0]), .o_cmd_1(
        o_inner_cmd_wire[8]), .o_cmd_2(o_inner_cmd_wire[16]), .o_cmd_3(
        o_inner_cmd_wire[24]), .o_cmd_4(o_inner_cmd_wire[32]), .o_cmd_5(
        o_inner_cmd_wire[40]), .o_cmd_6(o_inner_cmd_wire[48]), .o_cmd_7(
        o_inner_cmd_wire[56]), .i_en(i_en), .i_cmd(i_cmd[7:0]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 i_cmd_id_1__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[1]), .o_cmd_1(
        o_inner_cmd_wire[9]), .o_cmd_2(o_inner_cmd_wire[17]), .o_cmd_3(
        o_inner_cmd_wire[25]), .o_cmd_4(o_inner_cmd_wire[33]), .o_cmd_5(
        o_inner_cmd_wire[41]), .o_cmd_6(o_inner_cmd_wire[49]), .o_cmd_7(
        o_inner_cmd_wire[57]), .i_en(i_en), .i_cmd(i_cmd[15:8]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 i_cmd_id_2__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[2]), .o_cmd_1(
        o_inner_cmd_wire[10]), .o_cmd_2(o_inner_cmd_wire[18]), .o_cmd_3(
        o_inner_cmd_wire[26]), .o_cmd_4(o_inner_cmd_wire[34]), .o_cmd_5(
        o_inner_cmd_wire[42]), .o_cmd_6(o_inner_cmd_wire[50]), .o_cmd_7(
        o_inner_cmd_wire[58]), .i_en(i_en), .i_cmd(i_cmd[23:16]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 i_cmd_id_3__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[3]), .o_cmd_1(
        o_inner_cmd_wire[11]), .o_cmd_2(o_inner_cmd_wire[19]), .o_cmd_3(
        o_inner_cmd_wire[27]), .o_cmd_4(o_inner_cmd_wire[35]), .o_cmd_5(
        o_inner_cmd_wire[43]), .o_cmd_6(o_inner_cmd_wire[51]), .o_cmd_7(
        o_inner_cmd_wire[59]), .i_en(i_en), .i_cmd(i_cmd[31:24]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 i_cmd_id_4__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[4]), .o_cmd_1(
        o_inner_cmd_wire[12]), .o_cmd_2(o_inner_cmd_wire[20]), .o_cmd_3(
        o_inner_cmd_wire[28]), .o_cmd_4(o_inner_cmd_wire[36]), .o_cmd_5(
        o_inner_cmd_wire[44]), .o_cmd_6(o_inner_cmd_wire[52]), .o_cmd_7(
        o_inner_cmd_wire[60]), .i_en(i_en), .i_cmd(i_cmd[39:32]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 i_cmd_id_5__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[5]), .o_cmd_1(
        o_inner_cmd_wire[13]), .o_cmd_2(o_inner_cmd_wire[21]), .o_cmd_3(
        o_inner_cmd_wire[29]), .o_cmd_4(o_inner_cmd_wire[37]), .o_cmd_5(
        o_inner_cmd_wire[45]), .o_cmd_6(o_inner_cmd_wire[53]), .o_cmd_7(
        o_inner_cmd_wire[61]), .i_en(i_en), .i_cmd(i_cmd[47:40]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 i_cmd_id_6__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[6]), .o_cmd_1(
        o_inner_cmd_wire[14]), .o_cmd_2(o_inner_cmd_wire[22]), .o_cmd_3(
        o_inner_cmd_wire[30]), .o_cmd_4(o_inner_cmd_wire[38]), .o_cmd_5(
        o_inner_cmd_wire[46]), .o_cmd_6(o_inner_cmd_wire[54]), .o_cmd_7(
        o_inner_cmd_wire[62]), .i_en(i_en), .i_cmd(i_cmd[55:48]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 i_cmd_id_7__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[7]), .o_cmd_1(
        o_inner_cmd_wire[15]), .o_cmd_2(o_inner_cmd_wire[23]), .o_cmd_3(
        o_inner_cmd_wire[31]), .o_cmd_4(o_inner_cmd_wire[39]), .o_cmd_5(
        o_inner_cmd_wire[47]), .o_cmd_6(o_inner_cmd_wire[55]), .o_cmd_7(
        o_inner_cmd_wire[63]), .i_en(i_en), .i_cmd(i_cmd[63:56]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_0 bottom_half_0__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_0__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_0__inner_data_i_mux_tree_wire), .o_valid(n272), 
        .o_data_bus({n497, n498, n499, n500, n501, n502, n503, n504, n505, 
        n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
        n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[7:0]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_7 bottom_half_1__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_1__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_1__inner_data_i_mux_tree_wire), .o_valid(n271), 
        .o_data_bus({n465, n466, n467, n468, n469, n470, n471, n472, n473, 
        n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, 
        n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[15:8]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_6 bottom_half_2__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_2__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_2__inner_data_i_mux_tree_wire), .o_valid(n270), 
        .o_data_bus({n433, n434, n435, n436, n437, n438, n439, n440, n441, 
        n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
        n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[23:16]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_5 bottom_half_3__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_3__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_3__inner_data_i_mux_tree_wire), .o_valid(n269), 
        .o_data_bus({n401, n402, n403, n404, n405, n406, n407, n408, n409, 
        n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
        n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[31:24]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_4 bottom_half_4__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_4__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_4__inner_data_i_mux_tree_wire), .o_valid(n268), 
        .o_data_bus({n369, n370, n371, n372, n373, n374, n375, n376, n377, 
        n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
        n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[39:32]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_3 bottom_half_5__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_5__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_5__inner_data_i_mux_tree_wire), .o_valid(n267), 
        .o_data_bus({n337, n338, n339, n340, n341, n342, n343, n344, n345, 
        n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
        n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[47:40]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_2 bottom_half_6__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_6__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_6__inner_data_i_mux_tree_wire), .o_valid(n266), 
        .o_data_bus({n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[55:48]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_1 bottom_half_7__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_7__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_7__inner_data_i_mux_tree_wire), .o_valid(n265), 
        .o_data_bus({n273, n274, n275, n276, n277, n278, n279, n280, n281, 
        n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
        n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[63:56]) );
  BUFFD6BWP30P140LVT U1 ( .I(n528), .Z(o_data_bus[0]) );
  BUFFD6BWP30P140LVT U2 ( .I(n527), .Z(o_data_bus[1]) );
  BUFFD6BWP30P140LVT U3 ( .I(n526), .Z(o_data_bus[2]) );
  BUFFD6BWP30P140LVT U4 ( .I(n525), .Z(o_data_bus[3]) );
  BUFFD6BWP30P140LVT U5 ( .I(n524), .Z(o_data_bus[4]) );
  BUFFD6BWP30P140LVT U6 ( .I(n523), .Z(o_data_bus[5]) );
  BUFFD6BWP30P140LVT U7 ( .I(n522), .Z(o_data_bus[6]) );
  BUFFD6BWP30P140LVT U8 ( .I(n521), .Z(o_data_bus[7]) );
  BUFFD6BWP30P140LVT U9 ( .I(n520), .Z(o_data_bus[8]) );
  BUFFD6BWP30P140LVT U10 ( .I(n519), .Z(o_data_bus[9]) );
  BUFFD6BWP30P140LVT U11 ( .I(n518), .Z(o_data_bus[10]) );
  BUFFD6BWP30P140LVT U12 ( .I(n517), .Z(o_data_bus[11]) );
  BUFFD6BWP30P140LVT U13 ( .I(n516), .Z(o_data_bus[12]) );
  BUFFD6BWP30P140LVT U14 ( .I(n515), .Z(o_data_bus[13]) );
  BUFFD6BWP30P140LVT U15 ( .I(n514), .Z(o_data_bus[14]) );
  BUFFD6BWP30P140LVT U16 ( .I(n513), .Z(o_data_bus[15]) );
  BUFFD6BWP30P140LVT U17 ( .I(n512), .Z(o_data_bus[16]) );
  BUFFD6BWP30P140LVT U18 ( .I(n511), .Z(o_data_bus[17]) );
  BUFFD6BWP30P140LVT U19 ( .I(n510), .Z(o_data_bus[18]) );
  BUFFD6BWP30P140LVT U20 ( .I(n509), .Z(o_data_bus[19]) );
  BUFFD6BWP30P140LVT U21 ( .I(n508), .Z(o_data_bus[20]) );
  BUFFD6BWP30P140LVT U22 ( .I(n507), .Z(o_data_bus[21]) );
  BUFFD6BWP30P140LVT U23 ( .I(n506), .Z(o_data_bus[22]) );
  BUFFD6BWP30P140LVT U24 ( .I(n505), .Z(o_data_bus[23]) );
  BUFFD6BWP30P140LVT U25 ( .I(n504), .Z(o_data_bus[24]) );
  BUFFD6BWP30P140LVT U26 ( .I(n503), .Z(o_data_bus[25]) );
  BUFFD6BWP30P140LVT U27 ( .I(n502), .Z(o_data_bus[26]) );
  BUFFD6BWP30P140LVT U28 ( .I(n501), .Z(o_data_bus[27]) );
  BUFFD6BWP30P140LVT U29 ( .I(n500), .Z(o_data_bus[28]) );
  BUFFD6BWP30P140LVT U30 ( .I(n499), .Z(o_data_bus[29]) );
  BUFFD6BWP30P140LVT U31 ( .I(n498), .Z(o_data_bus[30]) );
  BUFFD6BWP30P140LVT U32 ( .I(n497), .Z(o_data_bus[31]) );
  BUFFD6BWP30P140LVT U33 ( .I(n496), .Z(o_data_bus[32]) );
  BUFFD6BWP30P140LVT U34 ( .I(n495), .Z(o_data_bus[33]) );
  BUFFD6BWP30P140LVT U35 ( .I(n494), .Z(o_data_bus[34]) );
  BUFFD6BWP30P140LVT U36 ( .I(n493), .Z(o_data_bus[35]) );
  BUFFD6BWP30P140LVT U37 ( .I(n492), .Z(o_data_bus[36]) );
  BUFFD6BWP30P140LVT U38 ( .I(n491), .Z(o_data_bus[37]) );
  BUFFD6BWP30P140LVT U39 ( .I(n490), .Z(o_data_bus[38]) );
  BUFFD6BWP30P140LVT U40 ( .I(n489), .Z(o_data_bus[39]) );
  BUFFD6BWP30P140LVT U41 ( .I(n488), .Z(o_data_bus[40]) );
  BUFFD6BWP30P140LVT U42 ( .I(n487), .Z(o_data_bus[41]) );
  BUFFD6BWP30P140LVT U43 ( .I(n486), .Z(o_data_bus[42]) );
  BUFFD6BWP30P140LVT U44 ( .I(n485), .Z(o_data_bus[43]) );
  BUFFD6BWP30P140LVT U45 ( .I(n484), .Z(o_data_bus[44]) );
  BUFFD6BWP30P140LVT U46 ( .I(n483), .Z(o_data_bus[45]) );
  BUFFD6BWP30P140LVT U47 ( .I(n482), .Z(o_data_bus[46]) );
  BUFFD6BWP30P140LVT U48 ( .I(n481), .Z(o_data_bus[47]) );
  BUFFD6BWP30P140LVT U49 ( .I(n480), .Z(o_data_bus[48]) );
  BUFFD6BWP30P140LVT U50 ( .I(n479), .Z(o_data_bus[49]) );
  BUFFD6BWP30P140LVT U51 ( .I(n478), .Z(o_data_bus[50]) );
  BUFFD6BWP30P140LVT U52 ( .I(n477), .Z(o_data_bus[51]) );
  BUFFD6BWP30P140LVT U53 ( .I(n476), .Z(o_data_bus[52]) );
  BUFFD6BWP30P140LVT U54 ( .I(n475), .Z(o_data_bus[53]) );
  BUFFD6BWP30P140LVT U55 ( .I(n474), .Z(o_data_bus[54]) );
  BUFFD6BWP30P140LVT U56 ( .I(n473), .Z(o_data_bus[55]) );
  BUFFD6BWP30P140LVT U57 ( .I(n472), .Z(o_data_bus[56]) );
  BUFFD6BWP30P140LVT U58 ( .I(n471), .Z(o_data_bus[57]) );
  BUFFD6BWP30P140LVT U59 ( .I(n470), .Z(o_data_bus[58]) );
  BUFFD6BWP30P140LVT U60 ( .I(n469), .Z(o_data_bus[59]) );
  BUFFD6BWP30P140LVT U61 ( .I(n468), .Z(o_data_bus[60]) );
  BUFFD6BWP30P140LVT U62 ( .I(n467), .Z(o_data_bus[61]) );
  BUFFD6BWP30P140LVT U63 ( .I(n466), .Z(o_data_bus[62]) );
  BUFFD6BWP30P140LVT U64 ( .I(n465), .Z(o_data_bus[63]) );
  BUFFD6BWP30P140LVT U65 ( .I(n464), .Z(o_data_bus[64]) );
  BUFFD6BWP30P140LVT U66 ( .I(n463), .Z(o_data_bus[65]) );
  BUFFD6BWP30P140LVT U67 ( .I(n462), .Z(o_data_bus[66]) );
  BUFFD6BWP30P140LVT U68 ( .I(n461), .Z(o_data_bus[67]) );
  BUFFD6BWP30P140LVT U69 ( .I(n460), .Z(o_data_bus[68]) );
  BUFFD6BWP30P140LVT U70 ( .I(n459), .Z(o_data_bus[69]) );
  BUFFD6BWP30P140LVT U71 ( .I(n458), .Z(o_data_bus[70]) );
  BUFFD6BWP30P140LVT U72 ( .I(n457), .Z(o_data_bus[71]) );
  BUFFD6BWP30P140LVT U73 ( .I(n456), .Z(o_data_bus[72]) );
  BUFFD6BWP30P140LVT U74 ( .I(n455), .Z(o_data_bus[73]) );
  BUFFD6BWP30P140LVT U75 ( .I(n454), .Z(o_data_bus[74]) );
  BUFFD6BWP30P140LVT U76 ( .I(n453), .Z(o_data_bus[75]) );
  BUFFD6BWP30P140LVT U77 ( .I(n452), .Z(o_data_bus[76]) );
  BUFFD6BWP30P140LVT U78 ( .I(n451), .Z(o_data_bus[77]) );
  BUFFD6BWP30P140LVT U79 ( .I(n450), .Z(o_data_bus[78]) );
  BUFFD6BWP30P140LVT U80 ( .I(n449), .Z(o_data_bus[79]) );
  BUFFD6BWP30P140LVT U81 ( .I(n448), .Z(o_data_bus[80]) );
  BUFFD6BWP30P140LVT U82 ( .I(n447), .Z(o_data_bus[81]) );
  BUFFD6BWP30P140LVT U83 ( .I(n446), .Z(o_data_bus[82]) );
  BUFFD6BWP30P140LVT U84 ( .I(n445), .Z(o_data_bus[83]) );
  BUFFD6BWP30P140LVT U85 ( .I(n444), .Z(o_data_bus[84]) );
  BUFFD6BWP30P140LVT U86 ( .I(n443), .Z(o_data_bus[85]) );
  BUFFD6BWP30P140LVT U87 ( .I(n442), .Z(o_data_bus[86]) );
  BUFFD6BWP30P140LVT U88 ( .I(n441), .Z(o_data_bus[87]) );
  BUFFD6BWP30P140LVT U89 ( .I(n440), .Z(o_data_bus[88]) );
  BUFFD6BWP30P140LVT U90 ( .I(n439), .Z(o_data_bus[89]) );
  BUFFD6BWP30P140LVT U91 ( .I(n438), .Z(o_data_bus[90]) );
  BUFFD6BWP30P140LVT U92 ( .I(n437), .Z(o_data_bus[91]) );
  BUFFD6BWP30P140LVT U93 ( .I(n436), .Z(o_data_bus[92]) );
  BUFFD6BWP30P140LVT U94 ( .I(n435), .Z(o_data_bus[93]) );
  BUFFD6BWP30P140LVT U95 ( .I(n434), .Z(o_data_bus[94]) );
  BUFFD6BWP30P140LVT U96 ( .I(n433), .Z(o_data_bus[95]) );
  BUFFD6BWP30P140LVT U97 ( .I(n432), .Z(o_data_bus[96]) );
  BUFFD6BWP30P140LVT U98 ( .I(n431), .Z(o_data_bus[97]) );
  BUFFD6BWP30P140LVT U99 ( .I(n430), .Z(o_data_bus[98]) );
  BUFFD6BWP30P140LVT U100 ( .I(n429), .Z(o_data_bus[99]) );
  BUFFD6BWP30P140LVT U101 ( .I(n428), .Z(o_data_bus[100]) );
  BUFFD6BWP30P140LVT U102 ( .I(n427), .Z(o_data_bus[101]) );
  BUFFD6BWP30P140LVT U103 ( .I(n426), .Z(o_data_bus[102]) );
  BUFFD6BWP30P140LVT U104 ( .I(n425), .Z(o_data_bus[103]) );
  BUFFD6BWP30P140LVT U105 ( .I(n424), .Z(o_data_bus[104]) );
  BUFFD6BWP30P140LVT U106 ( .I(n423), .Z(o_data_bus[105]) );
  BUFFD6BWP30P140LVT U107 ( .I(n422), .Z(o_data_bus[106]) );
  BUFFD6BWP30P140LVT U108 ( .I(n421), .Z(o_data_bus[107]) );
  BUFFD6BWP30P140LVT U109 ( .I(n420), .Z(o_data_bus[108]) );
  BUFFD6BWP30P140LVT U110 ( .I(n419), .Z(o_data_bus[109]) );
  BUFFD6BWP30P140LVT U111 ( .I(n418), .Z(o_data_bus[110]) );
  BUFFD6BWP30P140LVT U112 ( .I(n417), .Z(o_data_bus[111]) );
  BUFFD6BWP30P140LVT U113 ( .I(n416), .Z(o_data_bus[112]) );
  BUFFD6BWP30P140LVT U114 ( .I(n415), .Z(o_data_bus[113]) );
  BUFFD6BWP30P140LVT U115 ( .I(n414), .Z(o_data_bus[114]) );
  BUFFD6BWP30P140LVT U116 ( .I(n413), .Z(o_data_bus[115]) );
  BUFFD6BWP30P140LVT U117 ( .I(n412), .Z(o_data_bus[116]) );
  BUFFD6BWP30P140LVT U118 ( .I(n411), .Z(o_data_bus[117]) );
  BUFFD6BWP30P140LVT U119 ( .I(n410), .Z(o_data_bus[118]) );
  BUFFD6BWP30P140LVT U120 ( .I(n409), .Z(o_data_bus[119]) );
  BUFFD6BWP30P140LVT U121 ( .I(n408), .Z(o_data_bus[120]) );
  BUFFD6BWP30P140LVT U122 ( .I(n407), .Z(o_data_bus[121]) );
  BUFFD6BWP30P140LVT U123 ( .I(n406), .Z(o_data_bus[122]) );
  BUFFD6BWP30P140LVT U124 ( .I(n405), .Z(o_data_bus[123]) );
  BUFFD6BWP30P140LVT U125 ( .I(n404), .Z(o_data_bus[124]) );
  BUFFD6BWP30P140LVT U126 ( .I(n403), .Z(o_data_bus[125]) );
  BUFFD6BWP30P140LVT U127 ( .I(n402), .Z(o_data_bus[126]) );
  BUFFD6BWP30P140LVT U128 ( .I(n401), .Z(o_data_bus[127]) );
  BUFFD6BWP30P140LVT U129 ( .I(n400), .Z(o_data_bus[128]) );
  BUFFD6BWP30P140LVT U130 ( .I(n399), .Z(o_data_bus[129]) );
  BUFFD6BWP30P140LVT U131 ( .I(n398), .Z(o_data_bus[130]) );
  BUFFD6BWP30P140LVT U132 ( .I(n397), .Z(o_data_bus[131]) );
  BUFFD6BWP30P140LVT U133 ( .I(n396), .Z(o_data_bus[132]) );
  BUFFD6BWP30P140LVT U134 ( .I(n395), .Z(o_data_bus[133]) );
  BUFFD6BWP30P140LVT U135 ( .I(n394), .Z(o_data_bus[134]) );
  BUFFD6BWP30P140LVT U136 ( .I(n393), .Z(o_data_bus[135]) );
  BUFFD6BWP30P140LVT U137 ( .I(n392), .Z(o_data_bus[136]) );
  BUFFD6BWP30P140LVT U138 ( .I(n391), .Z(o_data_bus[137]) );
  BUFFD6BWP30P140LVT U139 ( .I(n390), .Z(o_data_bus[138]) );
  BUFFD6BWP30P140LVT U140 ( .I(n389), .Z(o_data_bus[139]) );
  BUFFD6BWP30P140LVT U141 ( .I(n388), .Z(o_data_bus[140]) );
  BUFFD6BWP30P140LVT U142 ( .I(n387), .Z(o_data_bus[141]) );
  BUFFD6BWP30P140LVT U143 ( .I(n386), .Z(o_data_bus[142]) );
  BUFFD6BWP30P140LVT U144 ( .I(n385), .Z(o_data_bus[143]) );
  BUFFD6BWP30P140LVT U145 ( .I(n384), .Z(o_data_bus[144]) );
  BUFFD6BWP30P140LVT U146 ( .I(n383), .Z(o_data_bus[145]) );
  BUFFD6BWP30P140LVT U147 ( .I(n382), .Z(o_data_bus[146]) );
  BUFFD6BWP30P140LVT U148 ( .I(n381), .Z(o_data_bus[147]) );
  BUFFD6BWP30P140LVT U149 ( .I(n380), .Z(o_data_bus[148]) );
  BUFFD6BWP30P140LVT U150 ( .I(n379), .Z(o_data_bus[149]) );
  BUFFD6BWP30P140LVT U151 ( .I(n378), .Z(o_data_bus[150]) );
  BUFFD6BWP30P140LVT U152 ( .I(n377), .Z(o_data_bus[151]) );
  BUFFD6BWP30P140LVT U153 ( .I(n376), .Z(o_data_bus[152]) );
  BUFFD6BWP30P140LVT U154 ( .I(n375), .Z(o_data_bus[153]) );
  BUFFD6BWP30P140LVT U155 ( .I(n374), .Z(o_data_bus[154]) );
  BUFFD6BWP30P140LVT U156 ( .I(n373), .Z(o_data_bus[155]) );
  BUFFD6BWP30P140LVT U157 ( .I(n372), .Z(o_data_bus[156]) );
  BUFFD6BWP30P140LVT U158 ( .I(n371), .Z(o_data_bus[157]) );
  BUFFD6BWP30P140LVT U159 ( .I(n370), .Z(o_data_bus[158]) );
  BUFFD6BWP30P140LVT U160 ( .I(n369), .Z(o_data_bus[159]) );
  BUFFD6BWP30P140LVT U161 ( .I(n368), .Z(o_data_bus[160]) );
  BUFFD6BWP30P140LVT U162 ( .I(n367), .Z(o_data_bus[161]) );
  BUFFD6BWP30P140LVT U163 ( .I(n366), .Z(o_data_bus[162]) );
  BUFFD6BWP30P140LVT U164 ( .I(n365), .Z(o_data_bus[163]) );
  BUFFD6BWP30P140LVT U165 ( .I(n364), .Z(o_data_bus[164]) );
  BUFFD6BWP30P140LVT U166 ( .I(n363), .Z(o_data_bus[165]) );
  BUFFD6BWP30P140LVT U167 ( .I(n362), .Z(o_data_bus[166]) );
  BUFFD6BWP30P140LVT U168 ( .I(n361), .Z(o_data_bus[167]) );
  BUFFD6BWP30P140LVT U169 ( .I(n360), .Z(o_data_bus[168]) );
  BUFFD6BWP30P140LVT U170 ( .I(n359), .Z(o_data_bus[169]) );
  BUFFD6BWP30P140LVT U171 ( .I(n358), .Z(o_data_bus[170]) );
  BUFFD6BWP30P140LVT U172 ( .I(n357), .Z(o_data_bus[171]) );
  BUFFD6BWP30P140LVT U173 ( .I(n356), .Z(o_data_bus[172]) );
  BUFFD6BWP30P140LVT U174 ( .I(n355), .Z(o_data_bus[173]) );
  BUFFD6BWP30P140LVT U175 ( .I(n354), .Z(o_data_bus[174]) );
  BUFFD6BWP30P140LVT U176 ( .I(n353), .Z(o_data_bus[175]) );
  BUFFD6BWP30P140LVT U177 ( .I(n352), .Z(o_data_bus[176]) );
  BUFFD6BWP30P140LVT U178 ( .I(n351), .Z(o_data_bus[177]) );
  BUFFD6BWP30P140LVT U179 ( .I(n350), .Z(o_data_bus[178]) );
  BUFFD6BWP30P140LVT U180 ( .I(n349), .Z(o_data_bus[179]) );
  BUFFD6BWP30P140LVT U181 ( .I(n348), .Z(o_data_bus[180]) );
  BUFFD6BWP30P140LVT U182 ( .I(n347), .Z(o_data_bus[181]) );
  BUFFD6BWP30P140LVT U183 ( .I(n346), .Z(o_data_bus[182]) );
  BUFFD6BWP30P140LVT U184 ( .I(n345), .Z(o_data_bus[183]) );
  BUFFD6BWP30P140LVT U185 ( .I(n344), .Z(o_data_bus[184]) );
  BUFFD6BWP30P140LVT U186 ( .I(n343), .Z(o_data_bus[185]) );
  BUFFD6BWP30P140LVT U187 ( .I(n342), .Z(o_data_bus[186]) );
  BUFFD6BWP30P140LVT U188 ( .I(n341), .Z(o_data_bus[187]) );
  BUFFD6BWP30P140LVT U189 ( .I(n340), .Z(o_data_bus[188]) );
  BUFFD6BWP30P140LVT U190 ( .I(n339), .Z(o_data_bus[189]) );
  BUFFD6BWP30P140LVT U191 ( .I(n338), .Z(o_data_bus[190]) );
  BUFFD6BWP30P140LVT U192 ( .I(n337), .Z(o_data_bus[191]) );
  BUFFD6BWP30P140LVT U193 ( .I(n336), .Z(o_data_bus[192]) );
  BUFFD6BWP30P140LVT U194 ( .I(n335), .Z(o_data_bus[193]) );
  BUFFD6BWP30P140LVT U195 ( .I(n334), .Z(o_data_bus[194]) );
  BUFFD6BWP30P140LVT U196 ( .I(n333), .Z(o_data_bus[195]) );
  BUFFD6BWP30P140LVT U197 ( .I(n332), .Z(o_data_bus[196]) );
  BUFFD6BWP30P140LVT U198 ( .I(n331), .Z(o_data_bus[197]) );
  BUFFD6BWP30P140LVT U199 ( .I(n330), .Z(o_data_bus[198]) );
  BUFFD6BWP30P140LVT U200 ( .I(n329), .Z(o_data_bus[199]) );
  BUFFD6BWP30P140LVT U201 ( .I(n328), .Z(o_data_bus[200]) );
  BUFFD6BWP30P140LVT U202 ( .I(n327), .Z(o_data_bus[201]) );
  BUFFD6BWP30P140LVT U203 ( .I(n326), .Z(o_data_bus[202]) );
  BUFFD6BWP30P140LVT U204 ( .I(n325), .Z(o_data_bus[203]) );
  BUFFD6BWP30P140LVT U205 ( .I(n324), .Z(o_data_bus[204]) );
  BUFFD6BWP30P140LVT U206 ( .I(n323), .Z(o_data_bus[205]) );
  BUFFD6BWP30P140LVT U207 ( .I(n322), .Z(o_data_bus[206]) );
  BUFFD6BWP30P140LVT U208 ( .I(n321), .Z(o_data_bus[207]) );
  BUFFD6BWP30P140LVT U209 ( .I(n320), .Z(o_data_bus[208]) );
  BUFFD6BWP30P140LVT U210 ( .I(n319), .Z(o_data_bus[209]) );
  BUFFD6BWP30P140LVT U211 ( .I(n318), .Z(o_data_bus[210]) );
  BUFFD6BWP30P140LVT U212 ( .I(n317), .Z(o_data_bus[211]) );
  BUFFD6BWP30P140LVT U213 ( .I(n316), .Z(o_data_bus[212]) );
  BUFFD6BWP30P140LVT U214 ( .I(n315), .Z(o_data_bus[213]) );
  BUFFD6BWP30P140LVT U215 ( .I(n314), .Z(o_data_bus[214]) );
  BUFFD6BWP30P140LVT U216 ( .I(n313), .Z(o_data_bus[215]) );
  BUFFD6BWP30P140LVT U217 ( .I(n312), .Z(o_data_bus[216]) );
  BUFFD6BWP30P140LVT U218 ( .I(n311), .Z(o_data_bus[217]) );
  BUFFD6BWP30P140LVT U219 ( .I(n310), .Z(o_data_bus[218]) );
  BUFFD6BWP30P140LVT U220 ( .I(n309), .Z(o_data_bus[219]) );
  BUFFD6BWP30P140LVT U221 ( .I(n308), .Z(o_data_bus[220]) );
  BUFFD6BWP30P140LVT U222 ( .I(n307), .Z(o_data_bus[221]) );
  BUFFD6BWP30P140LVT U223 ( .I(n306), .Z(o_data_bus[222]) );
  BUFFD6BWP30P140LVT U224 ( .I(n305), .Z(o_data_bus[223]) );
  BUFFD6BWP30P140LVT U225 ( .I(n304), .Z(o_data_bus[224]) );
  BUFFD6BWP30P140LVT U226 ( .I(n303), .Z(o_data_bus[225]) );
  BUFFD6BWP30P140LVT U227 ( .I(n302), .Z(o_data_bus[226]) );
  BUFFD6BWP30P140LVT U228 ( .I(n301), .Z(o_data_bus[227]) );
  BUFFD6BWP30P140LVT U229 ( .I(n300), .Z(o_data_bus[228]) );
  BUFFD6BWP30P140LVT U230 ( .I(n299), .Z(o_data_bus[229]) );
  BUFFD6BWP30P140LVT U231 ( .I(n298), .Z(o_data_bus[230]) );
  BUFFD6BWP30P140LVT U232 ( .I(n297), .Z(o_data_bus[231]) );
  BUFFD6BWP30P140LVT U233 ( .I(n296), .Z(o_data_bus[232]) );
  BUFFD6BWP30P140LVT U234 ( .I(n295), .Z(o_data_bus[233]) );
  BUFFD6BWP30P140LVT U235 ( .I(n294), .Z(o_data_bus[234]) );
  BUFFD6BWP30P140LVT U236 ( .I(n293), .Z(o_data_bus[235]) );
  BUFFD6BWP30P140LVT U237 ( .I(n292), .Z(o_data_bus[236]) );
  BUFFD6BWP30P140LVT U238 ( .I(n291), .Z(o_data_bus[237]) );
  BUFFD6BWP30P140LVT U239 ( .I(n290), .Z(o_data_bus[238]) );
  BUFFD6BWP30P140LVT U240 ( .I(n289), .Z(o_data_bus[239]) );
  BUFFD6BWP30P140LVT U241 ( .I(n288), .Z(o_data_bus[240]) );
  BUFFD6BWP30P140LVT U242 ( .I(n287), .Z(o_data_bus[241]) );
  BUFFD6BWP30P140LVT U243 ( .I(n286), .Z(o_data_bus[242]) );
  BUFFD6BWP30P140LVT U244 ( .I(n285), .Z(o_data_bus[243]) );
  BUFFD6BWP30P140LVT U245 ( .I(n284), .Z(o_data_bus[244]) );
  BUFFD6BWP30P140LVT U246 ( .I(n283), .Z(o_data_bus[245]) );
  BUFFD6BWP30P140LVT U247 ( .I(n282), .Z(o_data_bus[246]) );
  BUFFD6BWP30P140LVT U248 ( .I(n281), .Z(o_data_bus[247]) );
  BUFFD6BWP30P140LVT U249 ( .I(n280), .Z(o_data_bus[248]) );
  BUFFD6BWP30P140LVT U250 ( .I(n279), .Z(o_data_bus[249]) );
  BUFFD6BWP30P140LVT U251 ( .I(n278), .Z(o_data_bus[250]) );
  BUFFD6BWP30P140LVT U252 ( .I(n277), .Z(o_data_bus[251]) );
  BUFFD6BWP30P140LVT U253 ( .I(n276), .Z(o_data_bus[252]) );
  BUFFD6BWP30P140LVT U254 ( .I(n275), .Z(o_data_bus[253]) );
  BUFFD6BWP30P140LVT U255 ( .I(n274), .Z(o_data_bus[254]) );
  BUFFD6BWP30P140LVT U256 ( .I(n273), .Z(o_data_bus[255]) );
  BUFFD6BWP30P140LVT U257 ( .I(n272), .Z(o_valid[0]) );
  BUFFD6BWP30P140LVT U258 ( .I(n271), .Z(o_valid[1]) );
  BUFFD6BWP30P140LVT U259 ( .I(n270), .Z(o_valid[2]) );
  BUFFD6BWP30P140LVT U260 ( .I(n269), .Z(o_valid[3]) );
  BUFFD6BWP30P140LVT U261 ( .I(n268), .Z(o_valid[4]) );
  BUFFD6BWP30P140LVT U262 ( .I(n267), .Z(o_valid[5]) );
  BUFFD6BWP30P140LVT U263 ( .I(n266), .Z(o_valid[6]) );
  BUFFD6BWP30P140LVT U264 ( .I(n265), .Z(o_valid[7]) );
endmodule

