`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

//module glob_pe_controller(CLK, reset, boot_up, boot_up_local, boot_up_table_update, start, init_sram, table_parse, input_valid, glob_scen_noc_input_valid, delay_matrix_element, obj_id_element,from_glob_prefetch_start,  from_glob_prefetch_dest,  scenario_update, local_controller_id, from_glob_prefetch_stop, hardware_latency1, hardware_latency2, scenario_len, data_in, noc_out_0, noc_out_1, noc_out_2, noc_out_3, noc_out_4, noc_out_5, noc_out_6, noc_out_7, noc_out_8, noc_out_9, noc_out_10, noc_out_11, noc_out_12, noc_out_13, noc_out_14, noc_out_15, final_out_0, final_out_1, final_out_2, final_out_3, valid_bit, h_tree_input_data, htree_connected_addr, from_noc_output_valid_0, from_noc_output_valid_1, scenario_update_to_loc, prefetch_enable, direct_tap, ready);
//module glob_pe_controller(CLK, reset, boot_up, boot_up_local, boot_up_table_update, start, init_sram, table_parse, input_valid, glob_scen_noc_input_valid, delay_matrix_element, obj_id_element,from_glob_prefetch_start,  from_glob_prefetch_dest, local_controller_id, from_glob_prefetch_stop, hardware_latency1, hardware_latency2, scenario_len, data_in, noc_out_0, noc_out_1, noc_out_2, noc_out_3, noc_out_4, noc_out_5, noc_out_6, noc_out_7, noc_out_8, noc_out_9, noc_out_10, noc_out_11, noc_out_12, noc_out_13, noc_out_14, noc_out_15, final_out_0, final_out_1, final_out_2, valid_bit, h_tree_input_data, htree_connected_addr, from_noc_output_valid_0, from_noc_output_valid_1, scenario_update_to_loc, prefetch_enable, direct_tap, ready,scenario_update_global, input_block_scen_pipeline, load_same_scenario,  input_block_latency);
module glob_pe_controller(CLK, reset, boot_up_ext, boot_up_local_ext, boot_up_table_update_ext, start_ext, init_sram_ext, table_parse_ext, dft_clk_out, delay_matrix_element, obj_id_element,from_glob_prefetch_start,  from_glob_prefetch_dest, local_controller_id, from_glob_prefetch_stop, hardware_latency1, hardware_latency2, scenario_len, data_in, noc_out_0, noc_out_1, noc_out_2, noc_out_3, noc_out_4, noc_out_5, noc_out_6, noc_out_7, noc_out_8, noc_out_9, noc_out_10, noc_out_11, noc_out_12, noc_out_13, noc_out_14, noc_out_15, final_out_0, final_out_1, final_out_2, valid_bit, h_tree_input_data, htree_connected_addr, from_noc_output_valid_0, from_noc_output_valid_1, scenario_update_to_loc, prefetch_enable, direct_tap, ready,scenario_update_global, input_block_scen_pipeline, load_same_scenario,  input_block_latency, pe_controller_latency, interp_time_block_latency, doppler_time_block_latency, scenario_update_interp, scenario_update_doppler, scenario_update_rx, input_latency, loc_controller_latency, ddnoc_latency, scenario_update_doppler_real,pre_cycle_doppler,scenario_global_latency2, scenario_update_global2, scenario_interp_latency2, scenario_update_interp2, boot_up, boot_up_local, boot_up_table_update, start, init_sram, table_parse, dft_program_delay, scen_del_pe_config, scenario_del_global_internal_config);

    // parameter
    	parameter N_sample = 1024;
	parameter datawidth = 16;
	parameter address_vector_width = 4; //4; //can be 200 or 8: 8 for small tapeout
	parameter full_address_vector_width = 8; //4; //can be 200 or 8: 8 for small tapeout
	parameter N_obj = 4; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 4; // 16 local controllers in subscaled system
	parameter sample_address_width = 10; /// assuming 256 words: needs to change if arrangement is different
	parameter pe_sample_address_width = 8; /// assuming 256 words: needs to change if arrangement is different
	parameter packet_width = 2+2*datawidth + full_address_vector_width;
	parameter delay_length = 14; // log(id_width*N_sample)
	parameter obj_id_width = 2; // log(N_obj)
	parameter tapping_loc_packet_width = sample_address_width + obj_id_width; // log(N_obj)
	parameter scen_len_width = 14;   //needs to be revised
	parameter noc_output_half = 8;   //needs to be revised
	parameter num_loc_controller = 16;	
	parameter num_prefetch_config_width = 25;
	parameter scen_del_width = 3;   ///increase if pipelining increases
	parameter latency_width = 7;

//=== IO Ports ===//

     // Normal Mode Input
    	input CLK; // system clock, generated by VCO
	input reset;
	input start_ext;
	input init_sram_ext;
	input boot_up_ext;
	input boot_up_local_ext;
	input boot_up_table_update_ext;
	input table_parse_ext;
	//input input_valid;
	//input glob_scen_noc_input_valid;
	input [delay_length - 1:0] delay_matrix_element;
	input [obj_id_width - 1:0] obj_id_element;
	input [delay_length - 1:0] hardware_latency1;   ///keep as config to be input through spi?
	input [delay_length - 1:0] hardware_latency2;   /// keep as config to be input through spi?
	input [scen_len_width - 1:0] scenario_len;   /// keep as config to be input through spi?
	input [2*datawidth - 1:0] data_in;   /// keep as config to be input through spi?
        input [2*datawidth-1:0] noc_out_0;   
        input [2*datawidth-1:0] noc_out_1;   
        input [2*datawidth-1:0] noc_out_2;   
        input [2*datawidth-1:0] noc_out_3;   
        input [2*datawidth-1:0] noc_out_4;   
        input [2*datawidth-1:0] noc_out_5;   
        input [2*datawidth-1:0] noc_out_6;   
        input [2*datawidth-1:0] noc_out_7;    
        input [2*datawidth-1:0] noc_out_8;   
        input [2*datawidth-1:0] noc_out_9;   
        input [2*datawidth-1:0] noc_out_10;   
        input [2*datawidth-1:0] noc_out_11;   
        input [2*datawidth-1:0] noc_out_12;   
        input [2*datawidth-1:0] noc_out_13;   
        input [2*datawidth-1:0] noc_out_14;   
        input [2*datawidth-1:0] noc_out_15;   
	input [noc_output_half - 1:0] from_noc_output_valid_0;
	input [noc_output_half - 1:0] from_noc_output_valid_1;
	input direct_tap;
	input [delay_length - 1:0] input_block_latency;
	input [delay_length - 1:0] input_block_scen_pipeline;
	input load_same_scenario;
	input [latency_width - 1:0] scenario_global_latency2;
	input [latency_width - 1:0] scenario_interp_latency2;
	input [latency_width - 1:0] input_latency;
	input [latency_width - 1:0] loc_controller_latency;
	input [latency_width - 1:0] ddnoc_latency;
	input [latency_width - 1:0] pe_controller_latency;
	input [latency_width - 1:0] interp_time_block_latency;
	input [latency_width - 1:0] doppler_time_block_latency;
	input [8:0] pre_cycle_doppler;
	input dft_clk_out;
	input [5:0] dft_program_delay;
	input [latency_width - 1:0] scen_del_pe_config;
	input [latency_width - 1:0] scenario_del_global_internal_config;

    // output
	output [address_vector_width - 1:0] from_glob_prefetch_dest;
	output [sample_address_width - 1:0] from_glob_prefetch_start;
	output [sample_address_width - 1:0] from_glob_prefetch_stop;
	output prefetch_enable;
	output [id_width - 1:0] local_controller_id;
	output valid_bit;


	output reg [2*datawidth-1:0] final_out_0;
	output reg [2*datawidth-1:0] final_out_1;
	output reg [2*datawidth-1:0] final_out_2;
	//output reg [2*datawidth-1:0] final_out_3;

	output [11:0] htree_connected_addr;  //no of bits needs to be fixed once Htree is fixed
	output [2*datawidth - 1:0] h_tree_input_data;
	output scenario_update_to_loc;
	output scenario_update_global;
	output scenario_update_global2;

 	output ready;
	output scenario_update_interp;
	output scenario_update_interp2;
	output scenario_update_doppler;
	output scenario_update_rx;
	output scenario_update_doppler_real;
	output reg start;
	output reg init_sram;
	output reg boot_up;
	output reg boot_up_local;
	output reg boot_up_table_update;
	output reg table_parse;

endmodule    

