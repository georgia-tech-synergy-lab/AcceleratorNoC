
module crossbar_one_hot_comb ( i_valid, i_data_bus, o_valid, o_data_bus, i_en, 
        i_cmd );
  input [31:0] i_valid;
  input [1023:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [255:0] i_cmd;
  input i_en;
  wire   n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528;

  NR3D0P7BWP30P140LVT U6684 ( .A1(i_cmd[87]), .A2(i_cmd[95]), .A3(i_cmd[79]), 
        .ZN(n6418) );
  INVD1BWP30P140LVT U6685 ( .I(n6418), .ZN(n6420) );
  MAOI222D1BWP30P140LVT U6686 ( .A(i_cmd[87]), .B(i_cmd[95]), .C(i_cmd[79]), 
        .ZN(n6419) );
  ND2D1BWP30P140LVT U6687 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  MUX2D0BWP30P140LVT U6688 ( .I0(n6421), .I1(n6420), .S(i_cmd[71]), .Z(n6447)
         );
  NR3D0P7BWP30P140LVT U6689 ( .A1(i_cmd[127]), .A2(i_cmd[111]), .A3(i_cmd[119]), .ZN(n6422) );
  INVD1BWP30P140LVT U6690 ( .I(n6422), .ZN(n6424) );
  MAOI222D1BWP30P140LVT U6691 ( .A(i_cmd[127]), .B(i_cmd[111]), .C(i_cmd[119]), 
        .ZN(n6423) );
  ND2D1BWP30P140LVT U6692 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  MUX2NUD1BWP30P140LVT U6693 ( .I0(n6425), .I1(n6424), .S(i_cmd[103]), .ZN(
        n6465) );
  ND2D1BWP30P140LVT U6694 ( .A1(i_en), .A2(n6465), .ZN(n6462) );
  NR3D0P7BWP30P140LVT U6695 ( .A1(i_cmd[63]), .A2(i_cmd[55]), .A3(i_cmd[47]), 
        .ZN(n6426) );
  INVD1BWP30P140LVT U6696 ( .I(n6426), .ZN(n7662) );
  MAOI222D1BWP30P140LVT U6697 ( .A(i_cmd[63]), .B(i_cmd[55]), .C(i_cmd[47]), 
        .ZN(n6427) );
  ND2D1BWP30P140LVT U6698 ( .A1(n7662), .A2(n6427), .ZN(n6428) );
  MUX2NUD1BWP30P140LVT U6699 ( .I0(n6428), .I1(n7662), .S(i_cmd[39]), .ZN(
        n6461) );
  ND2D1BWP30P140LVT U6700 ( .A1(i_en), .A2(n6461), .ZN(n6464) );
  ND2D1BWP30P140LVT U6701 ( .A1(n6462), .A2(n6464), .ZN(n6452) );
  INVD1BWP30P140LVT U6702 ( .I(i_en), .ZN(n6832) );
  NR3D0P7BWP30P140LVT U6703 ( .A1(i_cmd[191]), .A2(i_cmd[183]), .A3(i_cmd[175]), .ZN(n6429) );
  INVD1BWP30P140LVT U6704 ( .I(n6429), .ZN(n6431) );
  MAOI222D1BWP30P140LVT U6705 ( .A(i_cmd[191]), .B(i_cmd[183]), .C(i_cmd[175]), 
        .ZN(n6430) );
  ND2D1BWP30P140LVT U6706 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  MUX2D0BWP30P140LVT U6707 ( .I0(n6432), .I1(n6431), .S(i_cmd[167]), .Z(n6456)
         );
  NR2D1BWP30P140LVT U6708 ( .A1(n6832), .A2(n6456), .ZN(n6469) );
  NR3D0P7BWP30P140LVT U6709 ( .A1(i_cmd[223]), .A2(i_cmd[215]), .A3(i_cmd[207]), .ZN(n6433) );
  INVD1BWP30P140LVT U6710 ( .I(n6433), .ZN(n7649) );
  MAOI222D1BWP30P140LVT U6711 ( .A(i_cmd[223]), .B(i_cmd[215]), .C(i_cmd[207]), 
        .ZN(n6434) );
  ND2D1BWP30P140LVT U6712 ( .A1(n7649), .A2(n6434), .ZN(n6435) );
  MUX2D0BWP30P140LVT U6713 ( .I0(n6435), .I1(n7649), .S(i_cmd[199]), .Z(n6468)
         );
  NR2D1BWP30P140LVT U6714 ( .A1(n6832), .A2(n6468), .ZN(n6455) );
  NR2D1BWP30P140LVT U6715 ( .A1(n6469), .A2(n6455), .ZN(n6473) );
  NR3D0P7BWP30P140LVT U6716 ( .A1(i_cmd[151]), .A2(i_cmd[143]), .A3(i_cmd[159]), .ZN(n6436) );
  INVD1BWP30P140LVT U6717 ( .I(n6436), .ZN(n6439) );
  MAOI222D1BWP30P140LVT U6718 ( .A(i_cmd[151]), .B(i_cmd[143]), .C(i_cmd[159]), 
        .ZN(n6437) );
  AOI21D1BWP30P140LVT U6719 ( .A1(n6437), .A2(n6439), .B(i_cmd[135]), .ZN(
        n6438) );
  AOI211D1BWP30P140LVT U6720 ( .A1(i_cmd[135]), .A2(n6439), .B(n6832), .C(
        n6438), .ZN(n6472) );
  INR2D1BWP30P140LVT U6721 ( .A1(n6473), .B1(n6472), .ZN(n6457) );
  INVD1BWP30P140LVT U6722 ( .I(i_cmd[7]), .ZN(n7652) );
  NR2D1BWP30P140LVT U6723 ( .A1(i_cmd[31]), .A2(n7652), .ZN(n6443) );
  INVD1BWP30P140LVT U6724 ( .I(i_cmd[31]), .ZN(n7647) );
  NR2D1BWP30P140LVT U6725 ( .A1(i_cmd[7]), .A2(n7647), .ZN(n6442) );
  INVD1BWP30P140LVT U6726 ( .I(i_cmd[15]), .ZN(n7646) );
  INVD1BWP30P140LVT U6727 ( .I(i_cmd[23]), .ZN(n7653) );
  AOI22D1BWP30P140LVT U6728 ( .A1(i_cmd[23]), .A2(i_cmd[15]), .B1(n7646), .B2(
        n7653), .ZN(n6441) );
  OAI22D1BWP30P140LVT U6729 ( .A1(i_cmd[23]), .A2(i_cmd[15]), .B1(i_cmd[31]), 
        .B2(i_cmd[7]), .ZN(n6440) );
  OAI31D1BWP30P140LVT U6730 ( .A1(n6443), .A2(n6442), .A3(n6441), .B(n6440), 
        .ZN(n6470) );
  INVD1BWP30P140LVT U6731 ( .I(n6470), .ZN(n6454) );
  ND2D1BWP30P140LVT U6732 ( .A1(i_en), .A2(n6454), .ZN(n6458) );
  ND2D1BWP30P140LVT U6733 ( .A1(n6457), .A2(n6458), .ZN(n6460) );
  NR2D1BWP30P140LVT U6734 ( .A1(n6452), .A2(n6460), .ZN(n6448) );
  NR3D0P7BWP30P140LVT U6735 ( .A1(i_cmd[247]), .A2(i_cmd[239]), .A3(i_cmd[255]), .ZN(n6444) );
  INVD1BWP30P140LVT U6736 ( .I(n6444), .ZN(n7661) );
  MAOI222D1BWP30P140LVT U6737 ( .A(i_cmd[247]), .B(i_cmd[239]), .C(i_cmd[255]), 
        .ZN(n6445) );
  ND2D1BWP30P140LVT U6738 ( .A1(n7661), .A2(n6445), .ZN(n6446) );
  MUX2D0BWP30P140LVT U6739 ( .I0(n6446), .I1(n7661), .S(i_cmd[231]), .Z(n6449)
         );
  NR2D1BWP30P140LVT U6740 ( .A1(n6832), .A2(n6449), .ZN(n6450) );
  ND3D1BWP30P140LVT U6741 ( .A1(n6447), .A2(n6448), .A3(n6450), .ZN(n7673) );
  NR2D1BWP30P140LVT U6742 ( .A1(n6832), .A2(n6447), .ZN(n6451) );
  ND3D1BWP30P140LVT U6743 ( .A1(n6451), .A2(n6449), .A3(n6448), .ZN(n7670) );
  INVD1BWP30P140LVT U6744 ( .I(n7670), .ZN(n7669) );
  NR2D1BWP30P140LVT U6745 ( .A1(n6451), .A2(n6450), .ZN(n6459) );
  INR2D1BWP30P140LVT U6746 ( .A1(n6459), .B1(n6452), .ZN(n6471) );
  IND2D1BWP30P140LVT U6747 ( .A1(n6472), .B1(n6471), .ZN(n6453) );
  NR2D1BWP30P140LVT U6748 ( .A1(n6454), .A2(n6453), .ZN(n6467) );
  ND3D1BWP30P140LVT U6749 ( .A1(n6456), .A2(n6455), .A3(n6467), .ZN(n7650) );
  IND3D1BWP30P140LVT U6750 ( .A1(n6458), .B1(n6457), .B2(n6471), .ZN(n7654) );
  IND2D1BWP30P140LVT U6751 ( .A1(n6460), .B1(n6459), .ZN(n6463) );
  NR3D0P7BWP30P140LVT U6752 ( .A1(n6462), .A2(n6461), .A3(n6463), .ZN(n7672)
         );
  INVD1BWP30P140LVT U6753 ( .I(n7672), .ZN(n7659) );
  OR3D1BWP30P140LVT U6754 ( .A1(n6465), .A2(n6464), .A3(n6463), .Z(n7674) );
  ND4D1BWP30P140LVT U6755 ( .A1(n7650), .A2(n7654), .A3(n7659), .A4(n7674), 
        .ZN(n6466) );
  INR3D0BWP30P140LVT U6756 ( .A1(n7673), .B1(n7669), .B2(n6466), .ZN(n6474) );
  ND3D1BWP30P140LVT U6757 ( .A1(n6469), .A2(n6468), .A3(n6467), .ZN(n7651) );
  ND4D1BWP30P140LVT U6758 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), 
        .ZN(n7664) );
  ND3D3BWP30P140LVT U6759 ( .A1(n6474), .A2(n7651), .A3(n7664), .ZN(o_valid[7]) );
  NR3D0P7BWP30P140LVT U6760 ( .A1(i_cmd[181]), .A2(i_cmd[189]), .A3(i_cmd[173]), .ZN(n6475) );
  INVD1BWP30P140LVT U6761 ( .I(n6475), .ZN(n6477) );
  MAOI222D1BWP30P140LVT U6762 ( .A(i_cmd[181]), .B(i_cmd[189]), .C(i_cmd[173]), 
        .ZN(n6476) );
  ND2D1BWP30P140LVT U6763 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  MUX2D0BWP30P140LVT U6764 ( .I0(n6478), .I1(n6477), .S(i_cmd[165]), .Z(n6521)
         );
  NR2D1BWP30P140LVT U6765 ( .A1(n6832), .A2(n6521), .ZN(n6525) );
  NR3D0P7BWP30P140LVT U6766 ( .A1(i_cmd[213]), .A2(i_cmd[205]), .A3(i_cmd[221]), .ZN(n6479) );
  INVD1BWP30P140LVT U6767 ( .I(n6479), .ZN(n6481) );
  MAOI222D1BWP30P140LVT U6768 ( .A(i_cmd[213]), .B(i_cmd[205]), .C(i_cmd[221]), 
        .ZN(n6480) );
  ND2D1BWP30P140LVT U6769 ( .A1(n6481), .A2(n6480), .ZN(n6482) );
  MUX2D0BWP30P140LVT U6770 ( .I0(n6482), .I1(n6481), .S(i_cmd[197]), .Z(n6524)
         );
  NR2D1BWP30P140LVT U6771 ( .A1(n6832), .A2(n6524), .ZN(n6520) );
  NR2D1BWP30P140LVT U6772 ( .A1(n6525), .A2(n6520), .ZN(n6511) );
  INVD1BWP30P140LVT U6773 ( .I(i_cmd[253]), .ZN(n6483) );
  INVD1BWP30P140LVT U6774 ( .I(i_cmd[237]), .ZN(n6485) );
  INVD1BWP30P140LVT U6775 ( .I(i_cmd[229]), .ZN(n6484) );
  ND4D1BWP30P140LVT U6776 ( .A1(n6483), .A2(n6485), .A3(n6484), .A4(i_cmd[245]), .ZN(n7549) );
  OR4D1BWP30P140LVT U6777 ( .A1(i_cmd[245]), .A2(i_cmd[229]), .A3(i_cmd[237]), 
        .A4(n6483), .Z(n7545) );
  OR4D1BWP30P140LVT U6778 ( .A1(i_cmd[245]), .A2(i_cmd[253]), .A3(i_cmd[237]), 
        .A4(n6484), .Z(n7556) );
  OR4D1BWP30P140LVT U6779 ( .A1(i_cmd[245]), .A2(i_cmd[253]), .A3(i_cmd[229]), 
        .A4(n6485), .Z(n7546) );
  ND4D1BWP30P140LVT U6780 ( .A1(n7549), .A2(n7545), .A3(n7556), .A4(n7546), 
        .ZN(n6518) );
  CKAN2D1BWP30P140LVT U6781 ( .A1(n6518), .A2(i_en), .Z(n6512) );
  INR2D1BWP30P140LVT U6782 ( .A1(n6511), .B1(n6512), .ZN(n6530) );
  NR3D0P7BWP30P140LVT U6783 ( .A1(i_cmd[29]), .A2(i_cmd[13]), .A3(i_cmd[21]), 
        .ZN(n6486) );
  INVD1BWP30P140LVT U6784 ( .I(n6486), .ZN(n6489) );
  MAOI222D1BWP30P140LVT U6785 ( .A(i_cmd[29]), .B(i_cmd[13]), .C(i_cmd[21]), 
        .ZN(n6487) );
  AOI21D1BWP30P140LVT U6786 ( .A1(n6489), .A2(n6487), .B(i_cmd[5]), .ZN(n6488)
         );
  AOI21D1BWP30P140LVT U6787 ( .A1(i_cmd[5]), .A2(n6489), .B(n6488), .ZN(n6528)
         );
  CKAN2D1BWP30P140LVT U6788 ( .A1(n6528), .A2(i_en), .Z(n6510) );
  INR2D1BWP30P140LVT U6789 ( .A1(n6530), .B1(n6510), .ZN(n6515) );
  NR3D0P7BWP30P140LVT U6790 ( .A1(i_cmd[141]), .A2(i_cmd[157]), .A3(i_cmd[149]), .ZN(n6493) );
  INVD1BWP30P140LVT U6791 ( .I(i_cmd[133]), .ZN(n6492) );
  MAOI222D1BWP30P140LVT U6792 ( .A(i_cmd[141]), .B(i_cmd[157]), .C(i_cmd[149]), 
        .ZN(n6490) );
  AOI21D1BWP30P140LVT U6793 ( .A1(n6490), .A2(n6492), .B(n6493), .ZN(n6491) );
  AOI211D1BWP30P140LVT U6794 ( .A1(n6493), .A2(n6492), .B(n6491), .C(n6832), 
        .ZN(n6531) );
  INR2D1BWP30P140LVT U6795 ( .A1(n6515), .B1(n6531), .ZN(n6506) );
  NR3D0P7BWP30P140LVT U6796 ( .A1(i_cmd[53]), .A2(i_cmd[61]), .A3(i_cmd[45]), 
        .ZN(n6494) );
  INVD1BWP30P140LVT U6797 ( .I(n6494), .ZN(n6496) );
  MAOI222D1BWP30P140LVT U6798 ( .A(i_cmd[53]), .B(i_cmd[61]), .C(i_cmd[45]), 
        .ZN(n6495) );
  ND2D1BWP30P140LVT U6799 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  MUX2NUD1BWP30P140LVT U6800 ( .I0(n6497), .I1(n6496), .S(i_cmd[37]), .ZN(
        n6527) );
  INR2D1BWP30P140LVT U6801 ( .A1(n6527), .B1(n6832), .ZN(n6507) );
  NR3D0P7BWP30P140LVT U6802 ( .A1(i_cmd[117]), .A2(i_cmd[125]), .A3(i_cmd[109]), .ZN(n6498) );
  INVD1BWP30P140LVT U6803 ( .I(n6498), .ZN(n7566) );
  MAOI222D1BWP30P140LVT U6804 ( .A(i_cmd[117]), .B(i_cmd[125]), .C(i_cmd[109]), 
        .ZN(n6499) );
  ND2D1BWP30P140LVT U6805 ( .A1(n7566), .A2(n6499), .ZN(n6500) );
  MUX2NUD1BWP30P140LVT U6806 ( .I0(n6500), .I1(n7566), .S(i_cmd[101]), .ZN(
        n6517) );
  ND2D1BWP30P140LVT U6807 ( .A1(i_en), .A2(n6517), .ZN(n6505) );
  NR3D0P7BWP30P140LVT U6808 ( .A1(i_cmd[85]), .A2(i_cmd[93]), .A3(i_cmd[77]), 
        .ZN(n6501) );
  INVD1BWP30P140LVT U6809 ( .I(n6501), .ZN(n7561) );
  MAOI222D1BWP30P140LVT U6810 ( .A(i_cmd[85]), .B(i_cmd[93]), .C(i_cmd[77]), 
        .ZN(n6502) );
  ND2D1BWP30P140LVT U6811 ( .A1(n7561), .A2(n6502), .ZN(n6503) );
  MUX2NUD1BWP30P140LVT U6812 ( .I0(n6503), .I1(n7561), .S(i_cmd[69]), .ZN(
        n6504) );
  ND2D1BWP30P140LVT U6813 ( .A1(i_en), .A2(n6504), .ZN(n6513) );
  ND2D1BWP30P140LVT U6814 ( .A1(n6505), .A2(n6513), .ZN(n6526) );
  INVD1BWP30P140LVT U6815 ( .I(n6526), .ZN(n6508) );
  ND3D1BWP30P140LVT U6816 ( .A1(n6506), .A2(n6507), .A3(n6508), .ZN(n7569) );
  INVD1BWP30P140LVT U6817 ( .I(n7569), .ZN(n7571) );
  INR4D0BWP30P140LVT U6818 ( .A1(n6506), .B1(n6527), .B2(n6505), .B3(n6504), 
        .ZN(n7568) );
  NR2D1BWP30P140LVT U6819 ( .A1(n6531), .A2(n6507), .ZN(n6514) );
  ND2D1BWP30P140LVT U6820 ( .A1(n6508), .A2(n6514), .ZN(n6509) );
  IND3D1BWP30P140LVT U6821 ( .A1(n6509), .B1(n6510), .B2(n6530), .ZN(n7557) );
  NR2D1BWP30P140LVT U6822 ( .A1(n6510), .A2(n6509), .ZN(n6519) );
  ND3D1BWP30P140LVT U6823 ( .A1(n6512), .A2(n6511), .A3(n6519), .ZN(n7555) );
  INVD1BWP30P140LVT U6824 ( .I(n6513), .ZN(n6516) );
  IND4D1BWP30P140LVT U6825 ( .A1(n6517), .B1(n6516), .B2(n6515), .B3(n6514), 
        .ZN(n7560) );
  INR2D1BWP30P140LVT U6826 ( .A1(n6519), .B1(n6518), .ZN(n6523) );
  ND3D1BWP30P140LVT U6827 ( .A1(n6521), .A2(n6520), .A3(n6523), .ZN(n7558) );
  ND4D1BWP30P140LVT U6828 ( .A1(n7557), .A2(n7555), .A3(n7560), .A4(n7558), 
        .ZN(n6522) );
  NR3D0P7BWP30P140LVT U6829 ( .A1(n7571), .A2(n7568), .A3(n6522), .ZN(n6532)
         );
  ND3D1BWP30P140LVT U6830 ( .A1(n6525), .A2(n6524), .A3(n6523), .ZN(n7559) );
  NR3D0P7BWP30P140LVT U6831 ( .A1(n6528), .A2(n6527), .A3(n6526), .ZN(n6529)
         );
  ND3D1BWP30P140LVT U6832 ( .A1(n6531), .A2(n6530), .A3(n6529), .ZN(n7572) );
  ND3D3BWP30P140LVT U6833 ( .A1(n6532), .A2(n7559), .A3(n7572), .ZN(o_valid[5]) );
  NR3D0P7BWP30P140LVT U6834 ( .A1(i_cmd[140]), .A2(i_cmd[156]), .A3(i_cmd[148]), .ZN(n6533) );
  INVD1BWP30P140LVT U6835 ( .I(n6533), .ZN(n9736) );
  MAOI222D1BWP30P140LVT U6836 ( .A(i_cmd[140]), .B(i_cmd[156]), .C(i_cmd[148]), 
        .ZN(n6534) );
  ND2D1BWP30P140LVT U6837 ( .A1(n9736), .A2(n6534), .ZN(n6535) );
  MUX2NUD1BWP30P140LVT U6838 ( .I0(n6535), .I1(n9736), .S(i_cmd[132]), .ZN(
        n6568) );
  ND2D1BWP30P140LVT U6839 ( .A1(i_en), .A2(n6568), .ZN(n6559) );
  NR3D0P7BWP30P140LVT U6840 ( .A1(i_cmd[116]), .A2(i_cmd[124]), .A3(i_cmd[108]), .ZN(n6536) );
  INVD1BWP30P140LVT U6841 ( .I(n6536), .ZN(n6539) );
  MAOI222D1BWP30P140LVT U6842 ( .A(i_cmd[116]), .B(i_cmd[124]), .C(i_cmd[108]), 
        .ZN(n6537) );
  AOI21D1BWP30P140LVT U6843 ( .A1(n6539), .A2(n6537), .B(i_cmd[100]), .ZN(
        n6538) );
  AO21D1BWP30P140LVT U6844 ( .A1(i_cmd[100]), .A2(n6539), .B(n6538), .Z(n6571)
         );
  NR2D1BWP30P140LVT U6845 ( .A1(n6571), .A2(n6832), .ZN(n6585) );
  NR3D0P7BWP30P140LVT U6846 ( .A1(i_cmd[84]), .A2(i_cmd[92]), .A3(i_cmd[76]), 
        .ZN(n6540) );
  INVD1BWP30P140LVT U6847 ( .I(n6540), .ZN(n9751) );
  MAOI222D1BWP30P140LVT U6848 ( .A(i_cmd[84]), .B(i_cmd[92]), .C(i_cmd[76]), 
        .ZN(n6541) );
  AOI21D1BWP30P140LVT U6849 ( .A1(n9751), .A2(n6541), .B(i_cmd[68]), .ZN(n6542) );
  AO21D1BWP30P140LVT U6850 ( .A1(i_cmd[68]), .A2(n9751), .B(n6542), .Z(n6584)
         );
  NR2D1BWP30P140LVT U6851 ( .A1(n6584), .A2(n6832), .ZN(n6570) );
  NR2D1BWP30P140LVT U6852 ( .A1(n6585), .A2(n6570), .ZN(n6560) );
  NR3D0P7BWP30P140LVT U6853 ( .A1(i_cmd[52]), .A2(i_cmd[60]), .A3(i_cmd[44]), 
        .ZN(n6543) );
  INVD1BWP30P140LVT U6854 ( .I(n6543), .ZN(n6545) );
  MAOI222D1BWP30P140LVT U6855 ( .A(i_cmd[52]), .B(i_cmd[60]), .C(i_cmd[44]), 
        .ZN(n6544) );
  ND2D1BWP30P140LVT U6856 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  MUX2NUD1BWP30P140LVT U6857 ( .I0(n6546), .I1(n6545), .S(i_cmd[36]), .ZN(
        n6563) );
  INR2D1BWP30P140LVT U6858 ( .A1(n6563), .B1(n6832), .ZN(n6581) );
  NR3D0P7BWP30P140LVT U6859 ( .A1(i_cmd[28]), .A2(i_cmd[12]), .A3(i_cmd[20]), 
        .ZN(n6547) );
  INVD1BWP30P140LVT U6860 ( .I(n6547), .ZN(n9734) );
  MAOI222D1BWP30P140LVT U6861 ( .A(i_cmd[28]), .B(i_cmd[12]), .C(i_cmd[20]), 
        .ZN(n6548) );
  ND2D1BWP30P140LVT U6862 ( .A1(n9734), .A2(n6548), .ZN(n6549) );
  MUX2NUD1BWP30P140LVT U6863 ( .I0(n6549), .I1(n9734), .S(i_cmd[4]), .ZN(n6582) );
  ND2D1BWP30P140LVT U6864 ( .A1(i_en), .A2(n6582), .ZN(n6562) );
  IND2D1BWP30P140LVT U6865 ( .A1(n6581), .B1(n6562), .ZN(n6565) );
  NR3D0P7BWP30P140LVT U6866 ( .A1(i_cmd[180]), .A2(i_cmd[188]), .A3(i_cmd[172]), .ZN(n6550) );
  INVD1BWP30P140LVT U6867 ( .I(n6550), .ZN(n9761) );
  MAOI222D1BWP30P140LVT U6868 ( .A(i_cmd[180]), .B(i_cmd[188]), .C(i_cmd[172]), 
        .ZN(n6551) );
  AOI21D1BWP30P140LVT U6869 ( .A1(n9761), .A2(n6551), .B(i_cmd[164]), .ZN(
        n6552) );
  AO21D1BWP30P140LVT U6870 ( .A1(i_cmd[164]), .A2(n9761), .B(n6552), .Z(n6578)
         );
  NR2D1BWP30P140LVT U6871 ( .A1(n6578), .A2(n6832), .ZN(n6575) );
  NR3D0P7BWP30P140LVT U6872 ( .A1(i_cmd[212]), .A2(i_cmd[204]), .A3(i_cmd[220]), .ZN(n6553) );
  INVD1BWP30P140LVT U6873 ( .I(n6553), .ZN(n9763) );
  MAOI222D1BWP30P140LVT U6874 ( .A(i_cmd[212]), .B(i_cmd[204]), .C(i_cmd[220]), 
        .ZN(n6554) );
  AOI21D1BWP30P140LVT U6875 ( .A1(n9763), .A2(n6554), .B(i_cmd[196]), .ZN(
        n6555) );
  AO21D1BWP30P140LVT U6876 ( .A1(i_cmd[196]), .A2(n9763), .B(n6555), .Z(n6574)
         );
  NR2D1BWP30P140LVT U6877 ( .A1(n6574), .A2(n6832), .ZN(n6577) );
  NR2D1BWP30P140LVT U6878 ( .A1(n6575), .A2(n6577), .ZN(n6566) );
  NR2D1BWP30P140LVT U6879 ( .A1(i_cmd[252]), .A2(i_cmd[236]), .ZN(n6556) );
  INVD1BWP30P140LVT U6880 ( .I(i_cmd[228]), .ZN(n6558) );
  ND3D1BWP30P140LVT U6881 ( .A1(n6556), .A2(i_cmd[244]), .A3(n6558), .ZN(n9743) );
  INVD1BWP30P140LVT U6882 ( .I(i_cmd[244]), .ZN(n6557) );
  IND4D1BWP30P140LVT U6883 ( .A1(i_cmd[252]), .B1(i_cmd[236]), .B2(n6558), 
        .B3(n6557), .ZN(n9756) );
  OR4D1BWP30P140LVT U6884 ( .A1(i_cmd[252]), .A2(i_cmd[236]), .A3(i_cmd[244]), 
        .A4(n6558), .Z(n9752) );
  IND4D1BWP30P140LVT U6885 ( .A1(i_cmd[236]), .B1(i_cmd[252]), .B2(n6558), 
        .B3(n6557), .ZN(n9735) );
  ND4D1BWP30P140LVT U6886 ( .A1(n9743), .A2(n9756), .A3(n9752), .A4(n9735), 
        .ZN(n6572) );
  ND2D1BWP30P140LVT U6887 ( .A1(n6572), .A2(i_en), .ZN(n6567) );
  ND2D1BWP30P140LVT U6888 ( .A1(n6566), .A2(n6567), .ZN(n6561) );
  NR2D1BWP30P140LVT U6889 ( .A1(n6565), .A2(n6561), .ZN(n6569) );
  IND3D1BWP30P140LVT U6890 ( .A1(n6559), .B1(n6560), .B2(n6569), .ZN(n9754) );
  ND2D1BWP30P140LVT U6891 ( .A1(n6560), .A2(n6559), .ZN(n6564) );
  NR2D1BWP30P140LVT U6892 ( .A1(n6564), .A2(n6561), .ZN(n6580) );
  INR3D0BWP30P140LVT U6893 ( .A1(n6580), .B1(n6563), .B2(n6562), .ZN(n9753) );
  NR2D1BWP30P140LVT U6894 ( .A1(n6565), .A2(n6564), .ZN(n6573) );
  IND3D1BWP30P140LVT U6895 ( .A1(n6567), .B1(n6566), .B2(n6573), .ZN(n9755) );
  INR2D1BWP30P140LVT U6896 ( .A1(n6569), .B1(n6568), .ZN(n6583) );
  ND3D1BWP30P140LVT U6897 ( .A1(n6571), .A2(n6570), .A3(n6583), .ZN(n9750) );
  INR2D1BWP30P140LVT U6898 ( .A1(n6573), .B1(n6572), .ZN(n6576) );
  ND3D1BWP30P140LVT U6899 ( .A1(n6575), .A2(n6574), .A3(n6576), .ZN(n9764) );
  ND3D1BWP30P140LVT U6900 ( .A1(n6578), .A2(n6577), .A3(n6576), .ZN(n9762) );
  ND4D1BWP30P140LVT U6901 ( .A1(n9755), .A2(n9750), .A3(n9764), .A4(n9762), 
        .ZN(n6579) );
  INR3D0BWP30P140LVT U6902 ( .A1(n9754), .B1(n9753), .B2(n6579), .ZN(n6586) );
  IND3D1BWP30P140LVT U6903 ( .A1(n6582), .B1(n6581), .B2(n6580), .ZN(n9749) );
  ND3D1BWP30P140LVT U6904 ( .A1(n6585), .A2(n6584), .A3(n6583), .ZN(n9748) );
  ND3D3BWP30P140LVT U6905 ( .A1(n6586), .A2(n9749), .A3(n9748), .ZN(o_valid[4]) );
  NR3D0P7BWP30P140LVT U6906 ( .A1(i_cmd[107]), .A2(i_cmd[115]), .A3(i_cmd[123]), .ZN(n6587) );
  INVD1BWP30P140LVT U6907 ( .I(n6587), .ZN(n6590) );
  MAOI222D1BWP30P140LVT U6908 ( .A(i_cmd[107]), .B(i_cmd[115]), .C(i_cmd[123]), 
        .ZN(n6588) );
  AOI21D1BWP30P140LVT U6909 ( .A1(n6590), .A2(n6588), .B(i_cmd[99]), .ZN(n6589) );
  AO21D1BWP30P140LVT U6910 ( .A1(i_cmd[99]), .A2(n6590), .B(n6589), .Z(n6614)
         );
  NR3D0P7BWP30P140LVT U6911 ( .A1(i_cmd[139]), .A2(i_cmd[155]), .A3(i_cmd[147]), .ZN(n6591) );
  INVD1BWP30P140LVT U6912 ( .I(n6591), .ZN(n11712) );
  MAOI222D1BWP30P140LVT U6913 ( .A(i_cmd[139]), .B(i_cmd[155]), .C(i_cmd[147]), 
        .ZN(n6592) );
  AOI21D1BWP30P140LVT U6914 ( .A1(n11712), .A2(n6592), .B(i_cmd[131]), .ZN(
        n6593) );
  AO21D1BWP30P140LVT U6915 ( .A1(i_cmd[131]), .A2(n11712), .B(n6593), .Z(n6622) );
  NR2D1BWP30P140LVT U6916 ( .A1(n6622), .A2(n6832), .ZN(n6641) );
  NR3D0P7BWP30P140LVT U6917 ( .A1(i_cmd[27]), .A2(i_cmd[11]), .A3(i_cmd[19]), 
        .ZN(n6594) );
  INVD1BWP30P140LVT U6918 ( .I(n6594), .ZN(n11702) );
  MAOI222D1BWP30P140LVT U6919 ( .A(i_cmd[27]), .B(i_cmd[11]), .C(i_cmd[19]), 
        .ZN(n6595) );
  AOI21D1BWP30P140LVT U6920 ( .A1(n11702), .A2(n6595), .B(i_cmd[3]), .ZN(n6596) );
  AO21D1BWP30P140LVT U6921 ( .A1(i_cmd[3]), .A2(n11702), .B(n6596), .Z(n6640)
         );
  NR2D1BWP30P140LVT U6922 ( .A1(n6640), .A2(n6832), .ZN(n6621) );
  NR2D1BWP30P140LVT U6923 ( .A1(n6641), .A2(n6621), .ZN(n6625) );
  NR3D0P7BWP30P140LVT U6924 ( .A1(i_cmd[179]), .A2(i_cmd[187]), .A3(i_cmd[171]), .ZN(n6597) );
  INVD1BWP30P140LVT U6925 ( .I(n6597), .ZN(n11746) );
  MAOI222D1BWP30P140LVT U6926 ( .A(i_cmd[179]), .B(i_cmd[187]), .C(i_cmd[171]), 
        .ZN(n6598) );
  ND2D1BWP30P140LVT U6927 ( .A1(n11746), .A2(n6598), .ZN(n6599) );
  MUX2D0BWP30P140LVT U6928 ( .I0(n6599), .I1(n11746), .S(i_cmd[163]), .Z(n6634) );
  NR2D1BWP30P140LVT U6929 ( .A1(n6832), .A2(n6634), .ZN(n6631) );
  NR3D0P7BWP30P140LVT U6930 ( .A1(i_cmd[211]), .A2(i_cmd[203]), .A3(i_cmd[219]), .ZN(n6600) );
  INVD1BWP30P140LVT U6931 ( .I(n6600), .ZN(n6602) );
  MAOI222D1BWP30P140LVT U6932 ( .A(i_cmd[211]), .B(i_cmd[203]), .C(i_cmd[219]), 
        .ZN(n6601) );
  ND2D1BWP30P140LVT U6933 ( .A1(n6602), .A2(n6601), .ZN(n6603) );
  MUX2D0BWP30P140LVT U6934 ( .I0(n6603), .I1(n6602), .S(i_cmd[195]), .Z(n6630)
         );
  NR2D1BWP30P140LVT U6935 ( .A1(n6832), .A2(n6630), .ZN(n6633) );
  NR2D1BWP30P140LVT U6936 ( .A1(n6631), .A2(n6633), .ZN(n6626) );
  INVD1BWP30P140LVT U6937 ( .I(i_cmd[227]), .ZN(n6605) );
  INVD1BWP30P140LVT U6938 ( .I(i_cmd[243]), .ZN(n6606) );
  INVD1BWP30P140LVT U6939 ( .I(i_cmd[235]), .ZN(n6604) );
  ND4D1BWP30P140LVT U6940 ( .A1(n6605), .A2(n6606), .A3(n6604), .A4(i_cmd[251]), .ZN(n11716) );
  OR4D1BWP30P140LVT U6941 ( .A1(i_cmd[251]), .A2(i_cmd[227]), .A3(i_cmd[243]), 
        .A4(n6604), .Z(n11739) );
  OR4D1BWP30P140LVT U6942 ( .A1(i_cmd[251]), .A2(i_cmd[235]), .A3(i_cmd[243]), 
        .A4(n6605), .Z(n11734) );
  OR4D1BWP30P140LVT U6943 ( .A1(i_cmd[251]), .A2(i_cmd[227]), .A3(i_cmd[235]), 
        .A4(n6606), .Z(n11714) );
  ND4D1BWP30P140LVT U6944 ( .A1(n11716), .A2(n11739), .A3(n11734), .A4(n11714), 
        .ZN(n6628) );
  CKAN2D1BWP30P140LVT U6945 ( .A1(n6628), .A2(i_en), .Z(n6627) );
  INR2D1BWP30P140LVT U6946 ( .A1(n6626), .B1(n6627), .ZN(n6618) );
  ND2D1BWP30P140LVT U6947 ( .A1(n6625), .A2(n6618), .ZN(n6616) );
  NR3D0P7BWP30P140LVT U6948 ( .A1(i_cmd[51]), .A2(i_cmd[59]), .A3(i_cmd[43]), 
        .ZN(n6607) );
  INVD1BWP30P140LVT U6949 ( .I(n6607), .ZN(n11720) );
  MAOI222D1BWP30P140LVT U6950 ( .A(i_cmd[51]), .B(i_cmd[59]), .C(i_cmd[43]), 
        .ZN(n6608) );
  ND2D1BWP30P140LVT U6951 ( .A1(n11720), .A2(n6608), .ZN(n6609) );
  MUX2NUD1BWP30P140LVT U6952 ( .I0(n6609), .I1(n11720), .S(i_cmd[35]), .ZN(
        n6620) );
  NR2D1BWP30P140LVT U6953 ( .A1(n6616), .A2(n6620), .ZN(n6636) );
  NR3D0P7BWP30P140LVT U6954 ( .A1(i_cmd[83]), .A2(i_cmd[91]), .A3(i_cmd[75]), 
        .ZN(n6610) );
  INVD1BWP30P140LVT U6955 ( .I(n6610), .ZN(n6613) );
  MAOI222D1BWP30P140LVT U6956 ( .A(i_cmd[83]), .B(i_cmd[91]), .C(i_cmd[75]), 
        .ZN(n6611) );
  AOI21D1BWP30P140LVT U6957 ( .A1(n6613), .A2(n6611), .B(i_cmd[67]), .ZN(n6612) );
  AO21D1BWP30P140LVT U6958 ( .A1(i_cmd[67]), .A2(n6613), .B(n6612), .Z(n6637)
         );
  NR2D1BWP30P140LVT U6959 ( .A1(n6637), .A2(n6832), .ZN(n6615) );
  ND3D1BWP30P140LVT U6960 ( .A1(n6614), .A2(n6636), .A3(n6615), .ZN(n11730) );
  CKAN2D1BWP30P140LVT U6961 ( .A1(n6620), .A2(i_en), .Z(n6624) );
  NR2D1BWP30P140LVT U6962 ( .A1(n6614), .A2(n6832), .ZN(n6638) );
  NR2D1BWP30P140LVT U6963 ( .A1(n6638), .A2(n6615), .ZN(n6617) );
  INVD1BWP30P140LVT U6964 ( .I(n6617), .ZN(n6623) );
  INR3D0BWP30P140LVT U6965 ( .A1(n6624), .B1(n6616), .B2(n6623), .ZN(n11729)
         );
  ND2D1BWP30P140LVT U6966 ( .A1(n6618), .A2(n6617), .ZN(n6619) );
  NR2D1BWP30P140LVT U6967 ( .A1(n6620), .A2(n6619), .ZN(n6639) );
  ND3D1BWP30P140LVT U6968 ( .A1(n6622), .A2(n6621), .A3(n6639), .ZN(n11736) );
  INR3D0BWP30P140LVT U6969 ( .A1(n6625), .B1(n6624), .B2(n6623), .ZN(n6629) );
  ND3D1BWP30P140LVT U6970 ( .A1(n6627), .A2(n6626), .A3(n6629), .ZN(n11738) );
  INR2D1BWP30P140LVT U6971 ( .A1(n6629), .B1(n6628), .ZN(n6632) );
  ND3D1BWP30P140LVT U6972 ( .A1(n6631), .A2(n6630), .A3(n6632), .ZN(n11755) );
  ND3D1BWP30P140LVT U6973 ( .A1(n6634), .A2(n6633), .A3(n6632), .ZN(n11752) );
  ND4D1BWP30P140LVT U6974 ( .A1(n11736), .A2(n11738), .A3(n11755), .A4(n11752), 
        .ZN(n6635) );
  INR3D0BWP30P140LVT U6975 ( .A1(n11730), .B1(n11729), .B2(n6635), .ZN(n6642)
         );
  ND3D1BWP30P140LVT U6976 ( .A1(n6638), .A2(n6637), .A3(n6636), .ZN(n11718) );
  ND3D1BWP30P140LVT U6977 ( .A1(n6641), .A2(n6640), .A3(n6639), .ZN(n11732) );
  ND3D3BWP30P140LVT U6978 ( .A1(n6642), .A2(n11718), .A3(n11732), .ZN(
        o_valid[3]) );
  NR3D0P7BWP30P140LVT U6979 ( .A1(i_cmd[112]), .A2(i_cmd[120]), .A3(i_cmd[104]), .ZN(n6643) );
  INVD1BWP30P140LVT U6980 ( .I(n6643), .ZN(n7767) );
  MAOI222D1BWP30P140LVT U6981 ( .A(i_cmd[112]), .B(i_cmd[120]), .C(i_cmd[104]), 
        .ZN(n6644) );
  AOI21D1BWP30P140LVT U6982 ( .A1(n7767), .A2(n6644), .B(i_cmd[96]), .ZN(n6645) );
  AO21D1BWP30P140LVT U6983 ( .A1(i_cmd[96]), .A2(n7767), .B(n6645), .Z(n6667)
         );
  NR3D0P7BWP30P140LVT U6984 ( .A1(i_cmd[24]), .A2(i_cmd[8]), .A3(i_cmd[16]), 
        .ZN(n6646) );
  INVD1BWP30P140LVT U6985 ( .I(n6646), .ZN(n7755) );
  MAOI222D1BWP30P140LVT U6986 ( .A(i_cmd[24]), .B(i_cmd[8]), .C(i_cmd[16]), 
        .ZN(n6647) );
  ND2D1BWP30P140LVT U6987 ( .A1(n7755), .A2(n6647), .ZN(n6648) );
  MUX2NUD1BWP30P140LVT U6988 ( .I0(n6648), .I1(n7755), .S(i_cmd[0]), .ZN(n6689) );
  ND2D1BWP30P140LVT U6989 ( .A1(i_en), .A2(n6689), .ZN(n6687) );
  NR3D0P7BWP30P140LVT U6990 ( .A1(i_cmd[136]), .A2(i_cmd[152]), .A3(i_cmd[144]), .ZN(n6649) );
  INVD1BWP30P140LVT U6991 ( .I(n6649), .ZN(n6651) );
  MAOI222D1BWP30P140LVT U6992 ( .A(i_cmd[136]), .B(i_cmd[152]), .C(i_cmd[144]), 
        .ZN(n6650) );
  ND2D1BWP30P140LVT U6993 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  MUX2NUD1BWP30P140LVT U6994 ( .I0(n6652), .I1(n6651), .S(i_cmd[128]), .ZN(
        n6686) );
  ND2D1BWP30P140LVT U6995 ( .A1(i_en), .A2(n6686), .ZN(n6688) );
  ND2D1BWP30P140LVT U6996 ( .A1(n6687), .A2(n6688), .ZN(n6669) );
  INVD1BWP30P140LVT U6997 ( .I(i_cmd[232]), .ZN(n6654) );
  OR4D1BWP30P140LVT U6998 ( .A1(i_cmd[224]), .A2(i_cmd[240]), .A3(i_cmd[248]), 
        .A4(n6654), .Z(n7757) );
  INVD1BWP30P140LVT U6999 ( .I(i_cmd[248]), .ZN(n6653) );
  IND4D1BWP30P140LVT U7000 ( .A1(i_cmd[224]), .B1(i_cmd[240]), .B2(n6653), 
        .B3(n6654), .ZN(n7751) );
  IND4D1BWP30P140LVT U7001 ( .A1(i_cmd[240]), .B1(i_cmd[224]), .B2(n6653), 
        .B3(n6654), .ZN(n7750) );
  NR2D1BWP30P140LVT U7002 ( .A1(i_cmd[224]), .A2(i_cmd[240]), .ZN(n6655) );
  ND3D1BWP30P140LVT U7003 ( .A1(i_cmd[248]), .A2(n6655), .A3(n6654), .ZN(n7754) );
  AN4D0BWP30P140LVT U7004 ( .A1(n7757), .A2(n7751), .A3(n7750), .A4(n7754), 
        .Z(n6670) );
  NR2D1BWP30P140LVT U7005 ( .A1(n6670), .A2(n6832), .ZN(n6678) );
  NR3D0P7BWP30P140LVT U7006 ( .A1(i_cmd[208]), .A2(i_cmd[200]), .A3(i_cmd[216]), .ZN(n6656) );
  INVD1BWP30P140LVT U7007 ( .I(n6656), .ZN(n7765) );
  MAOI222D1BWP30P140LVT U7008 ( .A(i_cmd[208]), .B(i_cmd[200]), .C(i_cmd[216]), 
        .ZN(n6657) );
  AOI21D1BWP30P140LVT U7009 ( .A1(n7765), .A2(n6657), .B(i_cmd[192]), .ZN(
        n6658) );
  AOI21D1BWP30P140LVT U7010 ( .A1(i_cmd[192]), .A2(n7765), .B(n6658), .ZN(
        n6671) );
  CKAN2D1BWP30P140LVT U7011 ( .A1(n6671), .A2(i_en), .Z(n6682) );
  OR3D1BWP30P140LVT U7012 ( .A1(i_cmd[176]), .A2(i_cmd[184]), .A3(i_cmd[168]), 
        .Z(n7775) );
  MAOI222D1BWP30P140LVT U7013 ( .A(i_cmd[176]), .B(i_cmd[184]), .C(i_cmd[168]), 
        .ZN(n6659) );
  AOI21D1BWP30P140LVT U7014 ( .A1(n7775), .A2(n6659), .B(i_cmd[160]), .ZN(
        n6660) );
  AO21D1BWP30P140LVT U7015 ( .A1(i_cmd[160]), .A2(n7775), .B(n6660), .Z(n6681)
         );
  NR2D1BWP30P140LVT U7016 ( .A1(n6681), .A2(n6832), .ZN(n6672) );
  NR2D1BWP30P140LVT U7017 ( .A1(n6682), .A2(n6672), .ZN(n6677) );
  IND2D1BWP30P140LVT U7018 ( .A1(n6678), .B1(n6677), .ZN(n6693) );
  NR2D1BWP30P140LVT U7019 ( .A1(n6669), .A2(n6693), .ZN(n6680) );
  NR3D0P7BWP30P140LVT U7020 ( .A1(i_cmd[48]), .A2(i_cmd[56]), .A3(i_cmd[40]), 
        .ZN(n6661) );
  INVD1BWP30P140LVT U7021 ( .I(n6661), .ZN(n6663) );
  MAOI222D1BWP30P140LVT U7022 ( .A(i_cmd[48]), .B(i_cmd[56]), .C(i_cmd[40]), 
        .ZN(n6662) );
  ND2D1BWP30P140LVT U7023 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  MUX2NUD1BWP30P140LVT U7024 ( .I0(n6664), .I1(n6663), .S(i_cmd[32]), .ZN(
        n6690) );
  INR2D1BWP30P140LVT U7025 ( .A1(n6680), .B1(n6690), .ZN(n6673) );
  OR3D1BWP30P140LVT U7026 ( .A1(i_cmd[80]), .A2(i_cmd[88]), .A3(i_cmd[72]), 
        .Z(n7752) );
  MAOI222D1BWP30P140LVT U7027 ( .A(i_cmd[80]), .B(i_cmd[88]), .C(i_cmd[72]), 
        .ZN(n6665) );
  AOI21D1BWP30P140LVT U7028 ( .A1(n7752), .A2(n6665), .B(i_cmd[64]), .ZN(n6666) );
  AO21D1BWP30P140LVT U7029 ( .A1(i_cmd[64]), .A2(n7752), .B(n6666), .Z(n6675)
         );
  NR2D1BWP30P140LVT U7030 ( .A1(n6675), .A2(n6832), .ZN(n6668) );
  AN3D1BWP30P140LVT U7031 ( .A1(n6667), .A2(n6673), .A3(n6668), .Z(n7778) );
  INR2D1BWP30P140LVT U7032 ( .A1(n6690), .B1(n6832), .ZN(n6679) );
  NR2D1BWP30P140LVT U7033 ( .A1(n6667), .A2(n6832), .ZN(n6674) );
  NR2D1BWP30P140LVT U7034 ( .A1(n6674), .A2(n6668), .ZN(n6691) );
  IND2D1BWP30P140LVT U7035 ( .A1(n6679), .B1(n6691), .ZN(n6685) );
  NR2D1BWP30P140LVT U7036 ( .A1(n6669), .A2(n6685), .ZN(n6676) );
  ND2D1BWP30P140LVT U7037 ( .A1(n6670), .A2(n6676), .ZN(n6683) );
  INR3D0BWP30P140LVT U7038 ( .A1(n6672), .B1(n6671), .B2(n6683), .ZN(n7776) );
  ND3D1BWP30P140LVT U7039 ( .A1(n6675), .A2(n6674), .A3(n6673), .ZN(n7774) );
  ND3D1BWP30P140LVT U7040 ( .A1(n6678), .A2(n6677), .A3(n6676), .ZN(n7756) );
  ND3D1BWP30P140LVT U7041 ( .A1(n6680), .A2(n6679), .A3(n6691), .ZN(n7760) );
  IND3D1BWP30P140LVT U7042 ( .A1(n6683), .B1(n6682), .B2(n6681), .ZN(n7779) );
  ND4D1BWP30P140LVT U7043 ( .A1(n7774), .A2(n7756), .A3(n7760), .A4(n7779), 
        .ZN(n6684) );
  NR3D0P7BWP30P140LVT U7044 ( .A1(n7778), .A2(n7776), .A3(n6684), .ZN(n6694)
         );
  OR4D1BWP30P140LVT U7045 ( .A1(n6687), .A2(n6686), .A3(n6693), .A4(n6685), 
        .Z(n7759) );
  INR4D0BWP30P140LVT U7046 ( .A1(n6691), .B1(n6690), .B2(n6689), .B3(n6688), 
        .ZN(n6692) );
  IND2D1BWP30P140LVT U7047 ( .A1(n6693), .B1(n6692), .ZN(n7769) );
  ND3D3BWP30P140LVT U7048 ( .A1(n6694), .A2(n7759), .A3(n7769), .ZN(o_valid[0]) );
  NR3D0P7BWP30P140LVT U7049 ( .A1(i_cmd[81]), .A2(i_cmd[73]), .A3(i_cmd[89]), 
        .ZN(n6695) );
  INVD1BWP30P140LVT U7050 ( .I(n6695), .ZN(n6698) );
  MAOI222D1BWP30P140LVT U7051 ( .A(i_cmd[81]), .B(i_cmd[73]), .C(i_cmd[89]), 
        .ZN(n6696) );
  AOI21D1BWP30P140LVT U7052 ( .A1(n6698), .A2(n6696), .B(i_cmd[65]), .ZN(n6697) );
  AO21D1BWP30P140LVT U7053 ( .A1(i_cmd[65]), .A2(n6698), .B(n6697), .Z(n6723)
         );
  NR3D0P7BWP30P140LVT U7054 ( .A1(i_cmd[113]), .A2(i_cmd[121]), .A3(i_cmd[105]), .ZN(n6699) );
  INVD1BWP30P140LVT U7055 ( .I(n6699), .ZN(n11016) );
  MAOI222D1BWP30P140LVT U7056 ( .A(i_cmd[113]), .B(i_cmd[121]), .C(i_cmd[105]), 
        .ZN(n6700) );
  AOI21D1BWP30P140LVT U7057 ( .A1(n11016), .A2(n6700), .B(i_cmd[97]), .ZN(
        n6701) );
  AO21D1BWP30P140LVT U7058 ( .A1(i_cmd[97]), .A2(n11016), .B(n6701), .Z(n6738)
         );
  NR2D1BWP30P140LVT U7059 ( .A1(n6738), .A2(n6832), .ZN(n6724) );
  NR3D0P7BWP30P140LVT U7060 ( .A1(i_cmd[49]), .A2(i_cmd[57]), .A3(i_cmd[41]), 
        .ZN(n6702) );
  INVD1BWP30P140LVT U7061 ( .I(n6702), .ZN(n6704) );
  MAOI222D1BWP30P140LVT U7062 ( .A(i_cmd[49]), .B(i_cmd[57]), .C(i_cmd[41]), 
        .ZN(n6703) );
  ND2D1BWP30P140LVT U7063 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  MUX2D0BWP30P140LVT U7064 ( .I0(n6705), .I1(n6704), .S(i_cmd[33]), .Z(n6734)
         );
  NR3D0P7BWP30P140LVT U7065 ( .A1(i_cmd[177]), .A2(i_cmd[185]), .A3(i_cmd[169]), .ZN(n6706) );
  INVD1BWP30P140LVT U7066 ( .I(n6706), .ZN(n11021) );
  MAOI222D1BWP30P140LVT U7067 ( .A(i_cmd[177]), .B(i_cmd[185]), .C(i_cmd[169]), 
        .ZN(n6707) );
  AOI21D1BWP30P140LVT U7068 ( .A1(n11021), .A2(n6707), .B(i_cmd[161]), .ZN(
        n6708) );
  AO21D1BWP30P140LVT U7069 ( .A1(i_cmd[161]), .A2(n11021), .B(n6708), .Z(n6727) );
  NR2D1BWP30P140LVT U7070 ( .A1(n6727), .A2(n6832), .ZN(n6730) );
  NR3D0P7BWP30P140LVT U7071 ( .A1(i_cmd[209]), .A2(i_cmd[201]), .A3(i_cmd[217]), .ZN(n6709) );
  INVD1BWP30P140LVT U7072 ( .I(n6709), .ZN(n11022) );
  MAOI222D1BWP30P140LVT U7073 ( .A(i_cmd[209]), .B(i_cmd[201]), .C(i_cmd[217]), 
        .ZN(n6710) );
  AOI21D1BWP30P140LVT U7074 ( .A1(n11022), .A2(n6710), .B(i_cmd[193]), .ZN(
        n6711) );
  AO21D1BWP30P140LVT U7075 ( .A1(i_cmd[193]), .A2(n11022), .B(n6711), .Z(n6729) );
  NR2D1BWP30P140LVT U7076 ( .A1(n6729), .A2(n6832), .ZN(n6726) );
  NR2D1BWP30P140LVT U7077 ( .A1(n6730), .A2(n6726), .ZN(n6742) );
  NR2D1BWP30P140LVT U7078 ( .A1(i_cmd[225]), .A2(i_cmd[241]), .ZN(n6712) );
  INVD1BWP30P140LVT U7079 ( .I(i_cmd[233]), .ZN(n6714) );
  ND3D1BWP30P140LVT U7080 ( .A1(n6712), .A2(i_cmd[249]), .A3(n6714), .ZN(
        n11004) );
  OR4D1BWP30P140LVT U7081 ( .A1(i_cmd[225]), .A2(i_cmd[241]), .A3(i_cmd[249]), 
        .A4(n6714), .Z(n11005) );
  INVD1BWP30P140LVT U7082 ( .I(i_cmd[249]), .ZN(n6713) );
  IND4D1BWP30P140LVT U7083 ( .A1(i_cmd[241]), .B1(i_cmd[225]), .B2(n6714), 
        .B3(n6713), .ZN(n11014) );
  IND4D1BWP30P140LVT U7084 ( .A1(i_cmd[225]), .B1(i_cmd[241]), .B2(n6714), 
        .B3(n6713), .ZN(n11012) );
  ND4D1BWP30P140LVT U7085 ( .A1(n11004), .A2(n11005), .A3(n11014), .A4(n11012), 
        .ZN(n6725) );
  CKAN2D1BWP30P140LVT U7086 ( .A1(n6725), .A2(i_en), .Z(n6743) );
  INR2D1BWP30P140LVT U7087 ( .A1(n6742), .B1(n6743), .ZN(n6744) );
  NR3D0P7BWP30P140LVT U7088 ( .A1(i_cmd[25]), .A2(i_cmd[9]), .A3(i_cmd[17]), 
        .ZN(n6715) );
  INVD1BWP30P140LVT U7089 ( .I(n6715), .ZN(n6718) );
  MAOI222D1BWP30P140LVT U7090 ( .A(i_cmd[25]), .B(i_cmd[9]), .C(i_cmd[17]), 
        .ZN(n6716) );
  AOI21D1BWP30P140LVT U7091 ( .A1(n6716), .A2(n6718), .B(i_cmd[1]), .ZN(n6717)
         );
  AOI211D1BWP30P140LVT U7092 ( .A1(i_cmd[1]), .A2(n6718), .B(n6832), .C(n6717), 
        .ZN(n6746) );
  INR2D1BWP30P140LVT U7093 ( .A1(n6744), .B1(n6746), .ZN(n6733) );
  NR3D0P7BWP30P140LVT U7094 ( .A1(i_cmd[137]), .A2(i_cmd[153]), .A3(i_cmd[145]), .ZN(n6722) );
  INVD1BWP30P140LVT U7095 ( .I(i_cmd[129]), .ZN(n6721) );
  MAOI222D1BWP30P140LVT U7096 ( .A(i_cmd[137]), .B(i_cmd[153]), .C(i_cmd[145]), 
        .ZN(n6719) );
  AOI21D1BWP30P140LVT U7097 ( .A1(n6719), .A2(n6721), .B(n6722), .ZN(n6720) );
  AOI211D1BWP30P140LVT U7098 ( .A1(n6722), .A2(n6721), .B(n6720), .C(n6832), 
        .ZN(n6736) );
  INR2D1BWP30P140LVT U7099 ( .A1(n6733), .B1(n6736), .ZN(n6731) );
  CKAN2D1BWP30P140LVT U7100 ( .A1(n6734), .A2(n6731), .Z(n6737) );
  ND3D1BWP30P140LVT U7101 ( .A1(n6723), .A2(n6724), .A3(n6737), .ZN(n11024) );
  NR2D1BWP30P140LVT U7102 ( .A1(n6723), .A2(n6832), .ZN(n6739) );
  NR2D1BWP30P140LVT U7103 ( .A1(n6739), .A2(n6724), .ZN(n6735) );
  NR2D1BWP30P140LVT U7104 ( .A1(n6832), .A2(n6734), .ZN(n6732) );
  INR3D0BWP30P140LVT U7105 ( .A1(n6735), .B1(n6736), .B2(n6732), .ZN(n6745) );
  INR2D1BWP30P140LVT U7106 ( .A1(n6745), .B1(n6746), .ZN(n6741) );
  INR2D1BWP30P140LVT U7107 ( .A1(n6741), .B1(n6725), .ZN(n6728) );
  ND3D1BWP30P140LVT U7108 ( .A1(n6727), .A2(n6726), .A3(n6728), .ZN(n11034) );
  ND3D1BWP30P140LVT U7109 ( .A1(n6730), .A2(n6729), .A3(n6728), .ZN(n11031) );
  ND3D1BWP30P140LVT U7110 ( .A1(n6735), .A2(n6732), .A3(n6731), .ZN(n11033) );
  ND4D1BWP30P140LVT U7111 ( .A1(n11024), .A2(n11034), .A3(n11031), .A4(n11033), 
        .ZN(n6740) );
  ND4D1BWP30P140LVT U7112 ( .A1(n6736), .A2(n6735), .A3(n6734), .A4(n6733), 
        .ZN(n11015) );
  ND3D1BWP30P140LVT U7113 ( .A1(n6739), .A2(n6738), .A3(n6737), .ZN(n11035) );
  IND3D1BWP30P140LVT U7114 ( .A1(n6740), .B1(n11015), .B2(n11035), .ZN(n6747)
         );
  ND3D1BWP30P140LVT U7115 ( .A1(n6743), .A2(n6742), .A3(n6741), .ZN(n11013) );
  ND3D1BWP30P140LVT U7116 ( .A1(n6746), .A2(n6745), .A3(n6744), .ZN(n11011) );
  IND3D4BWP30P140LVT U7117 ( .A1(n6747), .B1(n11013), .B2(n11011), .ZN(
        o_valid[1]) );
  NR3D0P7BWP30P140LVT U7118 ( .A1(i_cmd[182]), .A2(i_cmd[190]), .A3(i_cmd[174]), .ZN(n6748) );
  INVD1BWP30P140LVT U7119 ( .I(n6748), .ZN(n6751) );
  MAOI222D1BWP30P140LVT U7120 ( .A(i_cmd[182]), .B(i_cmd[190]), .C(i_cmd[174]), 
        .ZN(n6749) );
  AOI21D1BWP30P140LVT U7121 ( .A1(n6751), .A2(n6749), .B(i_cmd[166]), .ZN(
        n6750) );
  AO21D1BWP30P140LVT U7122 ( .A1(i_cmd[166]), .A2(n6751), .B(n6750), .Z(n6791)
         );
  NR2D1BWP30P140LVT U7123 ( .A1(n6791), .A2(n6832), .ZN(n6777) );
  NR3D0P7BWP30P140LVT U7124 ( .A1(i_cmd[214]), .A2(i_cmd[206]), .A3(i_cmd[222]), .ZN(n6752) );
  INVD1BWP30P140LVT U7125 ( .I(n6752), .ZN(n6755) );
  MAOI222D1BWP30P140LVT U7126 ( .A(i_cmd[214]), .B(i_cmd[206]), .C(i_cmd[222]), 
        .ZN(n6753) );
  AOI21D1BWP30P140LVT U7127 ( .A1(n6755), .A2(n6753), .B(i_cmd[198]), .ZN(
        n6754) );
  AO21D1BWP30P140LVT U7128 ( .A1(i_cmd[198]), .A2(n6755), .B(n6754), .Z(n6776)
         );
  NR3D0P7BWP30P140LVT U7129 ( .A1(i_cmd[86]), .A2(i_cmd[94]), .A3(i_cmd[78]), 
        .ZN(n6756) );
  INVD1BWP30P140LVT U7130 ( .I(n6756), .ZN(n6758) );
  MAOI222D1BWP30P140LVT U7131 ( .A(i_cmd[86]), .B(i_cmd[94]), .C(i_cmd[78]), 
        .ZN(n6757) );
  ND2D1BWP30P140LVT U7132 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  MUX2D0BWP30P140LVT U7133 ( .I0(n6759), .I1(n6758), .S(i_cmd[70]), .Z(n6785)
         );
  NR2D1BWP30P140LVT U7134 ( .A1(n6832), .A2(n6785), .ZN(n6781) );
  NR3D0P7BWP30P140LVT U7135 ( .A1(i_cmd[118]), .A2(i_cmd[126]), .A3(i_cmd[110]), .ZN(n6760) );
  INVD1BWP30P140LVT U7136 ( .I(n6760), .ZN(n10310) );
  MAOI222D1BWP30P140LVT U7137 ( .A(i_cmd[118]), .B(i_cmd[126]), .C(i_cmd[110]), 
        .ZN(n6761) );
  ND2D1BWP30P140LVT U7138 ( .A1(n10310), .A2(n6761), .ZN(n6762) );
  MUX2D0BWP30P140LVT U7139 ( .I0(n6762), .I1(n10310), .S(i_cmd[102]), .Z(n6780) );
  NR2D1BWP30P140LVT U7140 ( .A1(n6832), .A2(n6780), .ZN(n6784) );
  NR2D1BWP30P140LVT U7141 ( .A1(n6781), .A2(n6784), .ZN(n6800) );
  NR3D0P7BWP30P140LVT U7142 ( .A1(i_cmd[54]), .A2(i_cmd[62]), .A3(i_cmd[46]), 
        .ZN(n6763) );
  INVD1BWP30P140LVT U7143 ( .I(n6763), .ZN(n10321) );
  MAOI222D1BWP30P140LVT U7144 ( .A(i_cmd[54]), .B(i_cmd[62]), .C(i_cmd[46]), 
        .ZN(n6764) );
  AOI21D1BWP30P140LVT U7145 ( .A1(n10321), .A2(n6764), .B(i_cmd[38]), .ZN(
        n6765) );
  AO21D1BWP30P140LVT U7146 ( .A1(i_cmd[38]), .A2(n10321), .B(n6765), .Z(n6786)
         );
  NR2D1BWP30P140LVT U7147 ( .A1(n6786), .A2(n6832), .ZN(n6788) );
  NR3D0P7BWP30P140LVT U7148 ( .A1(i_cmd[142]), .A2(i_cmd[158]), .A3(i_cmd[150]), .ZN(n6766) );
  INVD1BWP30P140LVT U7149 ( .I(n6766), .ZN(n10317) );
  MAOI222D1BWP30P140LVT U7150 ( .A(i_cmd[142]), .B(i_cmd[158]), .C(i_cmd[150]), 
        .ZN(n6767) );
  AOI21D1BWP30P140LVT U7151 ( .A1(n10317), .A2(n6767), .B(i_cmd[134]), .ZN(
        n6768) );
  AO21D1BWP30P140LVT U7152 ( .A1(i_cmd[134]), .A2(n10317), .B(n6768), .Z(n6782) );
  NR2D1BWP30P140LVT U7153 ( .A1(n6782), .A2(n6832), .ZN(n6801) );
  INR3D0BWP30P140LVT U7154 ( .A1(n6800), .B1(n6788), .B2(n6801), .ZN(n6795) );
  NR3D0P7BWP30P140LVT U7155 ( .A1(i_cmd[30]), .A2(i_cmd[14]), .A3(i_cmd[22]), 
        .ZN(n6769) );
  INVD1BWP30P140LVT U7156 ( .I(n6769), .ZN(n6772) );
  MAOI222D1BWP30P140LVT U7157 ( .A(i_cmd[30]), .B(i_cmd[14]), .C(i_cmd[22]), 
        .ZN(n6770) );
  AOI21D1BWP30P140LVT U7158 ( .A1(n6772), .A2(n6770), .B(i_cmd[6]), .ZN(n6771)
         );
  AOI21D1BWP30P140LVT U7159 ( .A1(i_cmd[6]), .A2(n6772), .B(n6771), .ZN(n6798)
         );
  ND2D1BWP30P140LVT U7160 ( .A1(i_en), .A2(n6798), .ZN(n6779) );
  INVD1BWP30P140LVT U7161 ( .I(n6779), .ZN(n6793) );
  INVD1BWP30P140LVT U7162 ( .I(i_cmd[238]), .ZN(n6775) );
  INVD1BWP30P140LVT U7163 ( .I(i_cmd[254]), .ZN(n6774) );
  IND4D1BWP30P140LVT U7164 ( .A1(i_cmd[230]), .B1(i_cmd[246]), .B2(n6775), 
        .B3(n6774), .ZN(n10294) );
  NR2D1BWP30P140LVT U7165 ( .A1(i_cmd[230]), .A2(i_cmd[246]), .ZN(n6773) );
  ND3D1BWP30P140LVT U7166 ( .A1(i_cmd[254]), .A2(n6773), .A3(n6775), .ZN(
        n10293) );
  OR4D1BWP30P140LVT U7167 ( .A1(i_cmd[230]), .A2(i_cmd[246]), .A3(i_cmd[254]), 
        .A4(n6775), .Z(n10295) );
  IND4D1BWP30P140LVT U7168 ( .A1(i_cmd[246]), .B1(i_cmd[230]), .B2(n6775), 
        .B3(n6774), .ZN(n10297) );
  ND4D1BWP30P140LVT U7169 ( .A1(n10294), .A2(n10293), .A3(n10295), .A4(n10297), 
        .ZN(n6778) );
  INR3D0BWP30P140LVT U7170 ( .A1(n6795), .B1(n6793), .B2(n6778), .ZN(n6789) );
  ND3D1BWP30P140LVT U7171 ( .A1(n6777), .A2(n6776), .A3(n6789), .ZN(n10308) );
  NR2D1BWP30P140LVT U7172 ( .A1(n6776), .A2(n6832), .ZN(n6790) );
  NR2D1BWP30P140LVT U7173 ( .A1(n6777), .A2(n6790), .ZN(n6796) );
  CKAN2D1BWP30P140LVT U7174 ( .A1(n6778), .A2(i_en), .Z(n6797) );
  INR2D1BWP30P140LVT U7175 ( .A1(n6796), .B1(n6797), .ZN(n6792) );
  ND2D1BWP30P140LVT U7176 ( .A1(n6792), .A2(n6779), .ZN(n6783) );
  NR2D1BWP30P140LVT U7177 ( .A1(n6788), .A2(n6783), .ZN(n6799) );
  ND4D1BWP30P140LVT U7178 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6799), 
        .ZN(n10309) );
  NR2D1BWP30P140LVT U7179 ( .A1(n6801), .A2(n6783), .ZN(n6787) );
  ND4D1BWP30P140LVT U7180 ( .A1(n6786), .A2(n6785), .A3(n6784), .A4(n6787), 
        .ZN(n10322) );
  ND3D1BWP30P140LVT U7181 ( .A1(n6788), .A2(n6800), .A3(n6787), .ZN(n10323) );
  ND4D1BWP30P140LVT U7182 ( .A1(n10308), .A2(n10309), .A3(n10322), .A4(n10323), 
        .ZN(n6794) );
  ND3D1BWP30P140LVT U7183 ( .A1(n6791), .A2(n6790), .A3(n6789), .ZN(n10319) );
  ND3D1BWP30P140LVT U7184 ( .A1(n6795), .A2(n6793), .A3(n6792), .ZN(n10320) );
  IND3D1BWP30P140LVT U7185 ( .A1(n6794), .B1(n10319), .B2(n10320), .ZN(n6802)
         );
  IND4D1BWP30P140LVT U7186 ( .A1(n6798), .B1(n6797), .B2(n6796), .B3(n6795), 
        .ZN(n10296) );
  ND3D1BWP30P140LVT U7187 ( .A1(n6801), .A2(n6800), .A3(n6799), .ZN(n10316) );
  IND3D4BWP30P140LVT U7188 ( .A1(n6802), .B1(n10296), .B2(n10316), .ZN(
        o_valid[6]) );
  OR3D1BWP30P140LVT U7189 ( .A1(i_cmd[82]), .A2(i_cmd[90]), .A3(i_cmd[74]), 
        .Z(n6805) );
  MAOI222D1BWP30P140LVT U7190 ( .A(i_cmd[82]), .B(i_cmd[90]), .C(i_cmd[74]), 
        .ZN(n6803) );
  AOI21D1BWP30P140LVT U7191 ( .A1(n6805), .A2(n6803), .B(i_cmd[66]), .ZN(n6804) );
  AO21D1BWP30P140LVT U7192 ( .A1(i_cmd[66]), .A2(n6805), .B(n6804), .Z(n6828)
         );
  NR3D0P7BWP30P140LVT U7193 ( .A1(i_cmd[114]), .A2(i_cmd[122]), .A3(i_cmd[106]), .ZN(n6806) );
  INVD1BWP30P140LVT U7194 ( .I(n6806), .ZN(n6831) );
  MAOI222D1BWP30P140LVT U7195 ( .A(i_cmd[114]), .B(i_cmd[122]), .C(i_cmd[106]), 
        .ZN(n6807) );
  AOI21D1BWP30P140LVT U7196 ( .A1(n6831), .A2(n6807), .B(i_cmd[98]), .ZN(n6808) );
  AO21D1BWP30P140LVT U7197 ( .A1(i_cmd[98]), .A2(n6831), .B(n6808), .Z(n6830)
         );
  NR2D1BWP30P140LVT U7198 ( .A1(n6830), .A2(n6832), .ZN(n6834) );
  NR3D0P7BWP30P140LVT U7199 ( .A1(i_cmd[210]), .A2(i_cmd[202]), .A3(i_cmd[218]), .ZN(n6809) );
  INVD1BWP30P140LVT U7200 ( .I(n6809), .ZN(n6846) );
  MAOI222D1BWP30P140LVT U7201 ( .A(i_cmd[210]), .B(i_cmd[202]), .C(i_cmd[218]), 
        .ZN(n6810) );
  ND2D1BWP30P140LVT U7202 ( .A1(n6846), .A2(n6810), .ZN(n6811) );
  MUX2D0BWP30P140LVT U7203 ( .I0(n6811), .I1(n6846), .S(i_cmd[194]), .Z(n6842)
         );
  NR2D1BWP30P140LVT U7204 ( .A1(n6832), .A2(n6842), .ZN(n6839) );
  NR3D0P7BWP30P140LVT U7205 ( .A1(i_cmd[178]), .A2(i_cmd[186]), .A3(i_cmd[170]), .ZN(n6812) );
  INVD1BWP30P140LVT U7206 ( .I(n6812), .ZN(n6853) );
  MAOI222D1BWP30P140LVT U7207 ( .A(i_cmd[178]), .B(i_cmd[186]), .C(i_cmd[170]), 
        .ZN(n6813) );
  ND2D1BWP30P140LVT U7208 ( .A1(n6853), .A2(n6813), .ZN(n6814) );
  MUX2D0BWP30P140LVT U7209 ( .I0(n6814), .I1(n6853), .S(i_cmd[162]), .Z(n6838)
         );
  NR2D1BWP30P140LVT U7210 ( .A1(n6832), .A2(n6838), .ZN(n6841) );
  NR2D1BWP30P140LVT U7211 ( .A1(n6839), .A2(n6841), .ZN(n6860) );
  INVD1BWP30P140LVT U7212 ( .I(i_cmd[250]), .ZN(n6817) );
  INVD1BWP30P140LVT U7213 ( .I(i_cmd[234]), .ZN(n6816) );
  INVD1BWP30P140LVT U7214 ( .I(i_cmd[242]), .ZN(n6815) );
  ND4D1BWP30P140LVT U7215 ( .A1(n6817), .A2(n6816), .A3(n6815), .A4(i_cmd[226]), .ZN(n6870) );
  OR4D1BWP30P140LVT U7216 ( .A1(i_cmd[226]), .A2(i_cmd[250]), .A3(i_cmd[234]), 
        .A4(n6815), .Z(n6863) );
  OR4D1BWP30P140LVT U7217 ( .A1(i_cmd[226]), .A2(i_cmd[250]), .A3(i_cmd[242]), 
        .A4(n6816), .Z(n6872) );
  OR4D1BWP30P140LVT U7218 ( .A1(i_cmd[226]), .A2(i_cmd[242]), .A3(i_cmd[234]), 
        .A4(n6817), .Z(n6871) );
  ND4D1BWP30P140LVT U7219 ( .A1(n6870), .A2(n6863), .A3(n6872), .A4(n6871), 
        .ZN(n6837) );
  CKAN2D1BWP30P140LVT U7220 ( .A1(n6837), .A2(i_en), .Z(n6861) );
  INR2D1BWP30P140LVT U7221 ( .A1(n6860), .B1(n6861), .ZN(n6868) );
  NR3D0P7BWP30P140LVT U7222 ( .A1(i_cmd[26]), .A2(i_cmd[10]), .A3(i_cmd[18]), 
        .ZN(n6818) );
  INVD1BWP30P140LVT U7223 ( .I(n6818), .ZN(n6852) );
  MAOI222D1BWP30P140LVT U7224 ( .A(i_cmd[26]), .B(i_cmd[10]), .C(i_cmd[18]), 
        .ZN(n6819) );
  ND2D1BWP30P140LVT U7225 ( .A1(n6852), .A2(n6819), .ZN(n6820) );
  MUX2NUD1BWP30P140LVT U7226 ( .I0(n6820), .I1(n6852), .S(i_cmd[2]), .ZN(n6865) );
  INVD1BWP30P140LVT U7227 ( .I(n6865), .ZN(n6862) );
  NR2D1BWP30P140LVT U7228 ( .A1(n6832), .A2(n6862), .ZN(n6835) );
  NR3D0P7BWP30P140LVT U7229 ( .A1(i_cmd[138]), .A2(i_cmd[154]), .A3(i_cmd[146]), .ZN(n6824) );
  INVD1BWP30P140LVT U7230 ( .I(i_cmd[130]), .ZN(n6823) );
  MAOI222D1BWP30P140LVT U7231 ( .A(i_cmd[138]), .B(i_cmd[154]), .C(i_cmd[146]), 
        .ZN(n6821) );
  AOI21D1BWP30P140LVT U7232 ( .A1(n6821), .A2(n6823), .B(n6824), .ZN(n6822) );
  AOI211D1BWP30P140LVT U7233 ( .A1(n6824), .A2(n6823), .B(n6822), .C(n6832), 
        .ZN(n6869) );
  INR3D0BWP30P140LVT U7234 ( .A1(n6868), .B1(n6835), .B2(n6869), .ZN(n6845) );
  NR3D0P7BWP30P140LVT U7235 ( .A1(i_cmd[50]), .A2(i_cmd[58]), .A3(i_cmd[42]), 
        .ZN(n6825) );
  INVD1BWP30P140LVT U7236 ( .I(n6825), .ZN(n6851) );
  MAOI222D1BWP30P140LVT U7237 ( .A(i_cmd[50]), .B(i_cmd[58]), .C(i_cmd[42]), 
        .ZN(n6826) );
  ND2D1BWP30P140LVT U7238 ( .A1(n6851), .A2(n6826), .ZN(n6827) );
  MUX2NUD1BWP30P140LVT U7239 ( .I0(n6827), .I1(n6851), .S(i_cmd[34]), .ZN(
        n6866) );
  INR2D1BWP30P140LVT U7240 ( .A1(n6845), .B1(n6866), .ZN(n6829) );
  ND3D1BWP30P140LVT U7241 ( .A1(n6828), .A2(n6834), .A3(n6829), .ZN(n9731) );
  INVD1BWP30P140LVT U7242 ( .I(n9731), .ZN(n6858) );
  ND3D1BWP30P140LVT U7243 ( .A1(i_valid[13]), .A2(i_cmd[106]), .A3(n6858), 
        .ZN(n7437) );
  INVD1BWP30P140LVT U7244 ( .I(n7437), .ZN(n7523) );
  ND3D1BWP30P140LVT U7245 ( .A1(i_valid[15]), .A2(i_cmd[122]), .A3(n6858), 
        .ZN(n7524) );
  INVD1BWP30P140LVT U7246 ( .I(n7524), .ZN(n7459) );
  AOI22D1BWP30P140LVT U7247 ( .A1(i_data_bus[447]), .A2(n7523), .B1(
        i_data_bus[511]), .B2(n7459), .ZN(n6884) );
  NR2D1BWP30P140LVT U7248 ( .A1(n6828), .A2(n6832), .ZN(n6833) );
  AN3D1BWP30P140LVT U7249 ( .A1(n6830), .A2(n6829), .A3(n6833), .Z(n9728) );
  ND3D1BWP30P140LVT U7250 ( .A1(i_valid[8]), .A2(i_cmd[66]), .A3(n9728), .ZN(
        n7521) );
  INVD1BWP30P140LVT U7251 ( .I(n7521), .ZN(n7436) );
  INVD1BWP30P140LVT U7252 ( .I(i_valid[12]), .ZN(n11705) );
  NR3D0P7BWP30P140LVT U7253 ( .A1(n11705), .A2(n6831), .A3(n9731), .ZN(n7496)
         );
  AOI22D1BWP30P140LVT U7254 ( .A1(i_data_bus[287]), .A2(n7436), .B1(
        i_data_bus[415]), .B2(n7496), .ZN(n6883) );
  INVD1BWP30P140LVT U7255 ( .I(i_valid[1]), .ZN(n11737) );
  INR2D1BWP30P140LVT U7256 ( .A1(n6866), .B1(n6832), .ZN(n6843) );
  NR2D1BWP30P140LVT U7257 ( .A1(n6834), .A2(n6833), .ZN(n6844) );
  INVD1BWP30P140LVT U7258 ( .I(n6844), .ZN(n6864) );
  NR3D0P7BWP30P140LVT U7259 ( .A1(n6869), .A2(n6843), .A3(n6864), .ZN(n6859)
         );
  ND3D1BWP30P140LVT U7260 ( .A1(n6835), .A2(n6868), .A3(n6859), .ZN(n9724) );
  INR3D0BWP30P140LVT U7261 ( .A1(i_cmd[10]), .B1(n11737), .B2(n9724), .ZN(
        n7514) );
  INVD1BWP30P140LVT U7262 ( .I(i_valid[25]), .ZN(n11751) );
  IND2D1BWP30P140LVT U7263 ( .A1(n6835), .B1(n6859), .ZN(n6836) );
  NR2D1BWP30P140LVT U7264 ( .A1(n6837), .A2(n6836), .ZN(n6840) );
  ND3D1BWP30P140LVT U7265 ( .A1(n6839), .A2(n6838), .A3(n6840), .ZN(n9726) );
  INR3D0BWP30P140LVT U7266 ( .A1(i_cmd[202]), .B1(n11751), .B2(n9726), .ZN(
        n7513) );
  AOI22D1BWP30P140LVT U7267 ( .A1(i_data_bus[63]), .A2(n7514), .B1(
        i_data_bus[831]), .B2(n7513), .ZN(n6850) );
  INVD1BWP30P140LVT U7268 ( .I(i_valid[22]), .ZN(n11748) );
  ND3D1BWP30P140LVT U7269 ( .A1(n6842), .A2(n6841), .A3(n6840), .ZN(n9725) );
  INR3D0BWP30P140LVT U7270 ( .A1(i_cmd[178]), .B1(n11748), .B2(n9725), .ZN(
        n7510) );
  INVD1BWP30P140LVT U7271 ( .I(i_valid[23]), .ZN(n11750) );
  INR3D0BWP30P140LVT U7272 ( .A1(i_cmd[186]), .B1(n11750), .B2(n9725), .ZN(
        n7504) );
  AOI22D1BWP30P140LVT U7273 ( .A1(i_data_bus[735]), .A2(n7510), .B1(
        i_data_bus[767]), .B2(n7504), .ZN(n6849) );
  INVD1BWP30P140LVT U7274 ( .I(i_valid[3]), .ZN(n11726) );
  INR3D0BWP30P140LVT U7275 ( .A1(i_cmd[26]), .B1(n11726), .B2(n9724), .ZN(
        n7512) );
  INVD1BWP30P140LVT U7276 ( .I(i_valid[6]), .ZN(n11030) );
  ND3D1BWP30P140LVT U7277 ( .A1(n6845), .A2(n6844), .A3(n6843), .ZN(n9723) );
  INR3D0BWP30P140LVT U7278 ( .A1(i_cmd[50]), .B1(n11030), .B2(n9723), .ZN(
        n7502) );
  AOI22D1BWP30P140LVT U7279 ( .A1(i_data_bus[127]), .A2(n7512), .B1(
        i_data_bus[223]), .B2(n7502), .ZN(n6848) );
  INVD1BWP30P140LVT U7280 ( .I(i_valid[2]), .ZN(n11699) );
  INR3D0BWP30P140LVT U7281 ( .A1(i_cmd[18]), .B1(n11699), .B2(n9724), .ZN(
        n7511) );
  INVD1BWP30P140LVT U7282 ( .I(i_valid[24]), .ZN(n11754) );
  NR3D0P7BWP30P140LVT U7283 ( .A1(n11754), .A2(n6846), .A3(n9726), .ZN(n7516)
         );
  AOI22D1BWP30P140LVT U7284 ( .A1(i_data_bus[95]), .A2(n7511), .B1(
        i_data_bus[799]), .B2(n7516), .ZN(n6847) );
  AN4D0BWP30P140LVT U7285 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), 
        .Z(n6882) );
  ND3D1BWP30P140LVT U7286 ( .A1(i_valid[9]), .A2(i_cmd[74]), .A3(n9728), .ZN(
        n7394) );
  INVD1BWP30P140LVT U7287 ( .I(n7394), .ZN(n7494) );
  ND3D1BWP30P140LVT U7288 ( .A1(i_valid[11]), .A2(i_cmd[90]), .A3(n9728), .ZN(
        n7369) );
  INVD1BWP30P140LVT U7289 ( .I(n7369), .ZN(n7495) );
  AOI22D1BWP30P140LVT U7290 ( .A1(i_data_bus[319]), .A2(n7494), .B1(
        i_data_bus[383]), .B2(n7495), .ZN(n6880) );
  INVD1BWP30P140LVT U7291 ( .I(i_valid[26]), .ZN(n11745) );
  INR3D0BWP30P140LVT U7292 ( .A1(i_cmd[210]), .B1(n11745), .B2(n9726), .ZN(
        n7498) );
  INVD1BWP30P140LVT U7293 ( .I(i_valid[21]), .ZN(n11756) );
  INR3D0BWP30P140LVT U7294 ( .A1(i_cmd[170]), .B1(n11756), .B2(n9725), .ZN(
        n7509) );
  AOI22D1BWP30P140LVT U7295 ( .A1(i_data_bus[863]), .A2(n7498), .B1(
        i_data_bus[703]), .B2(n7509), .ZN(n6857) );
  INVD1BWP30P140LVT U7296 ( .I(i_valid[4]), .ZN(n11721) );
  NR3D0P7BWP30P140LVT U7297 ( .A1(n11721), .A2(n6851), .A3(n9723), .ZN(n7503)
         );
  INVD1BWP30P140LVT U7298 ( .I(i_valid[7]), .ZN(n11032) );
  INR3D0BWP30P140LVT U7299 ( .A1(i_cmd[58]), .B1(n11032), .B2(n9723), .ZN(
        n7501) );
  AOI22D1BWP30P140LVT U7300 ( .A1(i_data_bus[159]), .A2(n7503), .B1(
        i_data_bus[255]), .B2(n7501), .ZN(n6856) );
  INVD1BWP30P140LVT U7301 ( .I(i_valid[0]), .ZN(n11703) );
  NR3D0P7BWP30P140LVT U7302 ( .A1(n11703), .A2(n6852), .A3(n9724), .ZN(n7500)
         );
  INVD1BWP30P140LVT U7303 ( .I(i_valid[5]), .ZN(n11023) );
  INR3D0BWP30P140LVT U7304 ( .A1(i_cmd[42]), .B1(n11023), .B2(n9723), .ZN(
        n7515) );
  AOI22D1BWP30P140LVT U7305 ( .A1(i_data_bus[31]), .A2(n7500), .B1(
        i_data_bus[191]), .B2(n7515), .ZN(n6855) );
  INVD1BWP30P140LVT U7306 ( .I(i_valid[20]), .ZN(n11747) );
  NR3D0P7BWP30P140LVT U7307 ( .A1(n11747), .A2(n6853), .A3(n9725), .ZN(n7499)
         );
  INVD1BWP30P140LVT U7308 ( .I(i_valid[27]), .ZN(n11749) );
  INR3D0BWP30P140LVT U7309 ( .A1(i_cmd[218]), .B1(n11749), .B2(n9726), .ZN(
        n7497) );
  AOI22D1BWP30P140LVT U7310 ( .A1(i_data_bus[671]), .A2(n7499), .B1(
        i_data_bus[895]), .B2(n7497), .ZN(n6854) );
  ND4D1BWP30P140LVT U7311 ( .A1(n6857), .A2(n6856), .A3(n6855), .A4(n6854), 
        .ZN(n6879) );
  INVD1BWP30P140LVT U7312 ( .I(i_data_bus[479]), .ZN(n7766) );
  ND3D1BWP30P140LVT U7313 ( .A1(i_valid[14]), .A2(i_cmd[114]), .A3(n6858), 
        .ZN(n7522) );
  ND3D1BWP30P140LVT U7314 ( .A1(i_valid[10]), .A2(i_cmd[82]), .A3(n9728), .ZN(
        n7458) );
  INVD1BWP30P140LVT U7315 ( .I(n7458), .ZN(n7493) );
  MOAI22D1BWP30P140LVT U7316 ( .A1(n7766), .A2(n7522), .B1(i_data_bus[351]), 
        .B2(n7493), .ZN(n6878) );
  INVD1BWP30P140LVT U7317 ( .I(i_valid[30]), .ZN(n11715) );
  ND4D1BWP30P140LVT U7318 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), 
        .ZN(n9730) );
  NR3D0P7BWP30P140LVT U7319 ( .A1(n11715), .A2(n6863), .A3(n9730), .ZN(n7525)
         );
  INVD1BWP30P140LVT U7320 ( .I(i_valid[17]), .ZN(n11701) );
  NR3D0P7BWP30P140LVT U7321 ( .A1(n6866), .A2(n6865), .A3(n6864), .ZN(n6867)
         );
  ND3D1BWP30P140LVT U7322 ( .A1(n6869), .A2(n6868), .A3(n6867), .ZN(n9729) );
  INR3D0BWP30P140LVT U7323 ( .A1(i_cmd[138]), .B1(n11701), .B2(n9729), .ZN(
        n7526) );
  AOI22D1BWP30P140LVT U7324 ( .A1(i_data_bus[991]), .A2(n7525), .B1(
        i_data_bus[575]), .B2(n7526), .ZN(n6876) );
  INVD1BWP30P140LVT U7325 ( .I(i_valid[28]), .ZN(n11735) );
  NR3D0P7BWP30P140LVT U7326 ( .A1(n11735), .A2(n6870), .A3(n9730), .ZN(n7527)
         );
  INVD1BWP30P140LVT U7327 ( .I(i_valid[19]), .ZN(n11697) );
  INR3D0BWP30P140LVT U7328 ( .A1(i_cmd[154]), .B1(n11697), .B2(n9729), .ZN(
        n7529) );
  AOI22D1BWP30P140LVT U7329 ( .A1(i_data_bus[927]), .A2(n7527), .B1(
        i_data_bus[639]), .B2(n7529), .ZN(n6875) );
  INVD1BWP30P140LVT U7330 ( .I(i_valid[31]), .ZN(n11717) );
  NR3D0P7BWP30P140LVT U7331 ( .A1(n11717), .A2(n6871), .A3(n9730), .ZN(n7532)
         );
  INVD1BWP30P140LVT U7332 ( .I(i_valid[18]), .ZN(n11733) );
  INR3D0BWP30P140LVT U7333 ( .A1(i_cmd[146]), .B1(n11733), .B2(n9729), .ZN(
        n7531) );
  AOI22D1BWP30P140LVT U7334 ( .A1(i_data_bus[1023]), .A2(n7532), .B1(
        i_data_bus[607]), .B2(n7531), .ZN(n6874) );
  INVD1BWP30P140LVT U7335 ( .I(i_valid[16]), .ZN(n11713) );
  NR3D0P7BWP30P140LVT U7336 ( .A1(n11713), .A2(n6823), .A3(n9729), .ZN(n7530)
         );
  INVD1BWP30P140LVT U7337 ( .I(i_valid[29]), .ZN(n11740) );
  NR3D0P7BWP30P140LVT U7338 ( .A1(n11740), .A2(n6872), .A3(n9730), .ZN(n7528)
         );
  AOI22D1BWP30P140LVT U7339 ( .A1(i_data_bus[543]), .A2(n7530), .B1(
        i_data_bus[959]), .B2(n7528), .ZN(n6873) );
  ND4D1BWP30P140LVT U7340 ( .A1(n6876), .A2(n6875), .A3(n6874), .A4(n6873), 
        .ZN(n6877) );
  INR4D0BWP30P140LVT U7341 ( .A1(n6880), .B1(n6879), .B2(n6878), .B3(n6877), 
        .ZN(n6881) );
  ND4D4BWP30P140LVT U7342 ( .A1(n6884), .A2(n6883), .A3(n6882), .A4(n6881), 
        .ZN(o_data_bus[95]) );
  AOI22D1BWP30P140LVT U7343 ( .A1(i_data_bus[446]), .A2(n7523), .B1(
        i_data_bus[510]), .B2(n7459), .ZN(n6904) );
  AOI22D1BWP30P140LVT U7344 ( .A1(i_data_bus[350]), .A2(n7493), .B1(
        i_data_bus[318]), .B2(n7494), .ZN(n6903) );
  AOI22D1BWP30P140LVT U7345 ( .A1(i_data_bus[766]), .A2(n7504), .B1(
        i_data_bus[830]), .B2(n7513), .ZN(n6888) );
  AOI22D1BWP30P140LVT U7346 ( .A1(i_data_bus[670]), .A2(n7499), .B1(
        i_data_bus[190]), .B2(n7515), .ZN(n6887) );
  AOI22D1BWP30P140LVT U7347 ( .A1(i_data_bus[862]), .A2(n7498), .B1(
        i_data_bus[798]), .B2(n7516), .ZN(n6886) );
  AOI22D1BWP30P140LVT U7348 ( .A1(i_data_bus[62]), .A2(n7514), .B1(
        i_data_bus[894]), .B2(n7497), .ZN(n6885) );
  AN4D0BWP30P140LVT U7349 ( .A1(n6888), .A2(n6887), .A3(n6886), .A4(n6885), 
        .Z(n6902) );
  AOI22D1BWP30P140LVT U7350 ( .A1(i_data_bus[286]), .A2(n7436), .B1(
        i_data_bus[382]), .B2(n7495), .ZN(n6900) );
  AOI22D1BWP30P140LVT U7351 ( .A1(i_data_bus[734]), .A2(n7510), .B1(
        i_data_bus[158]), .B2(n7503), .ZN(n6892) );
  AOI22D1BWP30P140LVT U7352 ( .A1(i_data_bus[126]), .A2(n7512), .B1(
        i_data_bus[254]), .B2(n7501), .ZN(n6891) );
  AOI22D1BWP30P140LVT U7353 ( .A1(i_data_bus[94]), .A2(n7511), .B1(
        i_data_bus[222]), .B2(n7502), .ZN(n6890) );
  AOI22D1BWP30P140LVT U7354 ( .A1(i_data_bus[30]), .A2(n7500), .B1(
        i_data_bus[702]), .B2(n7509), .ZN(n6889) );
  ND4D1BWP30P140LVT U7355 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), 
        .ZN(n6899) );
  INVD1BWP30P140LVT U7356 ( .I(i_data_bus[414]), .ZN(n9224) );
  INVD1BWP30P140LVT U7357 ( .I(n7496), .ZN(n7411) );
  INVD1BWP30P140LVT U7358 ( .I(n7522), .ZN(n7472) );
  MOAI22D1BWP30P140LVT U7359 ( .A1(n9224), .A2(n7411), .B1(i_data_bus[478]), 
        .B2(n7472), .ZN(n6898) );
  AOI22D1BWP30P140LVT U7360 ( .A1(i_data_bus[958]), .A2(n7528), .B1(
        i_data_bus[1022]), .B2(n7532), .ZN(n6896) );
  AOI22D1BWP30P140LVT U7361 ( .A1(i_data_bus[926]), .A2(n7527), .B1(
        i_data_bus[990]), .B2(n7525), .ZN(n6895) );
  AOI22D1BWP30P140LVT U7362 ( .A1(i_data_bus[606]), .A2(n7531), .B1(
        i_data_bus[638]), .B2(n7529), .ZN(n6894) );
  AOI22D1BWP30P140LVT U7363 ( .A1(i_data_bus[542]), .A2(n7530), .B1(
        i_data_bus[574]), .B2(n7526), .ZN(n6893) );
  ND4D1BWP30P140LVT U7364 ( .A1(n6896), .A2(n6895), .A3(n6894), .A4(n6893), 
        .ZN(n6897) );
  INR4D0BWP30P140LVT U7365 ( .A1(n6900), .B1(n6899), .B2(n6898), .B3(n6897), 
        .ZN(n6901) );
  ND4D4BWP30P140LVT U7366 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), 
        .ZN(o_data_bus[94]) );
  AOI22D1BWP30P140LVT U7367 ( .A1(i_data_bus[365]), .A2(n7495), .B1(
        i_data_bus[461]), .B2(n7472), .ZN(n6924) );
  AOI22D1BWP30P140LVT U7368 ( .A1(i_data_bus[429]), .A2(n7523), .B1(
        i_data_bus[333]), .B2(n7493), .ZN(n6923) );
  AOI22D1BWP30P140LVT U7369 ( .A1(i_data_bus[525]), .A2(n7530), .B1(
        i_data_bus[621]), .B2(n7529), .ZN(n6908) );
  AOI22D1BWP30P140LVT U7370 ( .A1(i_data_bus[973]), .A2(n7525), .B1(
        i_data_bus[941]), .B2(n7528), .ZN(n6907) );
  AOI22D1BWP30P140LVT U7371 ( .A1(i_data_bus[557]), .A2(n7526), .B1(
        i_data_bus[1005]), .B2(n7532), .ZN(n6906) );
  AOI22D1BWP30P140LVT U7372 ( .A1(i_data_bus[909]), .A2(n7527), .B1(
        i_data_bus[589]), .B2(n7531), .ZN(n6905) );
  AN4D0BWP30P140LVT U7373 ( .A1(n6908), .A2(n6907), .A3(n6906), .A4(n6905), 
        .Z(n6922) );
  AOI22D1BWP30P140LVT U7374 ( .A1(i_data_bus[397]), .A2(n7496), .B1(
        i_data_bus[269]), .B2(n7436), .ZN(n6920) );
  INVD1BWP30P140LVT U7375 ( .I(i_data_bus[493]), .ZN(n8866) );
  MOAI22D1BWP30P140LVT U7376 ( .A1(n8866), .A2(n7524), .B1(i_data_bus[301]), 
        .B2(n7494), .ZN(n6919) );
  AOI22D1BWP30P140LVT U7377 ( .A1(i_data_bus[749]), .A2(n7504), .B1(
        i_data_bus[173]), .B2(n7515), .ZN(n6912) );
  AOI22D1BWP30P140LVT U7378 ( .A1(i_data_bus[77]), .A2(n7511), .B1(
        i_data_bus[141]), .B2(n7503), .ZN(n6911) );
  AOI22D1BWP30P140LVT U7379 ( .A1(i_data_bus[45]), .A2(n7514), .B1(
        i_data_bus[813]), .B2(n7513), .ZN(n6910) );
  AOI22D1BWP30P140LVT U7380 ( .A1(i_data_bus[781]), .A2(n7516), .B1(
        i_data_bus[205]), .B2(n7502), .ZN(n6909) );
  ND4D1BWP30P140LVT U7381 ( .A1(n6912), .A2(n6911), .A3(n6910), .A4(n6909), 
        .ZN(n6918) );
  AOI22D1BWP30P140LVT U7382 ( .A1(i_data_bus[685]), .A2(n7509), .B1(
        i_data_bus[717]), .B2(n7510), .ZN(n6916) );
  AOI22D1BWP30P140LVT U7383 ( .A1(i_data_bus[109]), .A2(n7512), .B1(
        i_data_bus[653]), .B2(n7499), .ZN(n6915) );
  AOI22D1BWP30P140LVT U7384 ( .A1(i_data_bus[13]), .A2(n7500), .B1(
        i_data_bus[877]), .B2(n7497), .ZN(n6914) );
  AOI22D1BWP30P140LVT U7385 ( .A1(i_data_bus[237]), .A2(n7501), .B1(
        i_data_bus[845]), .B2(n7498), .ZN(n6913) );
  ND4D1BWP30P140LVT U7386 ( .A1(n6916), .A2(n6915), .A3(n6914), .A4(n6913), 
        .ZN(n6917) );
  INR4D0BWP30P140LVT U7387 ( .A1(n6920), .B1(n6919), .B2(n6918), .B3(n6917), 
        .ZN(n6921) );
  ND4D4BWP30P140LVT U7388 ( .A1(n6924), .A2(n6923), .A3(n6922), .A4(n6921), 
        .ZN(o_data_bus[77]) );
  AOI22D1BWP30P140LVT U7389 ( .A1(i_data_bus[445]), .A2(n7523), .B1(
        i_data_bus[413]), .B2(n7496), .ZN(n6944) );
  AOI22D1BWP30P140LVT U7390 ( .A1(i_data_bus[349]), .A2(n7493), .B1(
        i_data_bus[477]), .B2(n7472), .ZN(n6943) );
  AOI22D1BWP30P140LVT U7391 ( .A1(i_data_bus[765]), .A2(n7504), .B1(
        i_data_bus[733]), .B2(n7510), .ZN(n6928) );
  AOI22D1BWP30P140LVT U7392 ( .A1(i_data_bus[29]), .A2(n7500), .B1(
        i_data_bus[61]), .B2(n7514), .ZN(n6927) );
  AOI22D1BWP30P140LVT U7393 ( .A1(i_data_bus[701]), .A2(n7509), .B1(
        i_data_bus[669]), .B2(n7499), .ZN(n6926) );
  AOI22D1BWP30P140LVT U7394 ( .A1(i_data_bus[861]), .A2(n7498), .B1(
        i_data_bus[221]), .B2(n7502), .ZN(n6925) );
  AN4D0BWP30P140LVT U7395 ( .A1(n6928), .A2(n6927), .A3(n6926), .A4(n6925), 
        .Z(n6942) );
  AOI22D1BWP30P140LVT U7396 ( .A1(i_data_bus[125]), .A2(n7512), .B1(
        i_data_bus[893]), .B2(n7497), .ZN(n6932) );
  AOI22D1BWP30P140LVT U7397 ( .A1(i_data_bus[93]), .A2(n7511), .B1(
        i_data_bus[797]), .B2(n7516), .ZN(n6931) );
  AOI22D1BWP30P140LVT U7398 ( .A1(i_data_bus[189]), .A2(n7515), .B1(
        i_data_bus[253]), .B2(n7501), .ZN(n6930) );
  AOI22D1BWP30P140LVT U7399 ( .A1(i_data_bus[157]), .A2(n7503), .B1(
        i_data_bus[829]), .B2(n7513), .ZN(n6929) );
  ND4D1BWP30P140LVT U7400 ( .A1(n6932), .A2(n6931), .A3(n6930), .A4(n6929), 
        .ZN(n6940) );
  INVD1BWP30P140LVT U7401 ( .I(i_data_bus[381]), .ZN(n7836) );
  INVD1BWP30P140LVT U7402 ( .I(i_data_bus[285]), .ZN(n8740) );
  OAI22D1BWP30P140LVT U7403 ( .A1(n7836), .A2(n7369), .B1(n8740), .B2(n7521), 
        .ZN(n6939) );
  INVD1BWP30P140LVT U7404 ( .I(i_data_bus[509]), .ZN(n7567) );
  MOAI22D1BWP30P140LVT U7405 ( .A1(n7567), .A2(n7524), .B1(i_data_bus[317]), 
        .B2(n7494), .ZN(n6938) );
  AOI22D1BWP30P140LVT U7406 ( .A1(i_data_bus[1021]), .A2(n7532), .B1(
        i_data_bus[541]), .B2(n7530), .ZN(n6936) );
  AOI22D1BWP30P140LVT U7407 ( .A1(i_data_bus[637]), .A2(n7529), .B1(
        i_data_bus[989]), .B2(n7525), .ZN(n6935) );
  AOI22D1BWP30P140LVT U7408 ( .A1(i_data_bus[925]), .A2(n7527), .B1(
        i_data_bus[605]), .B2(n7531), .ZN(n6934) );
  AOI22D1BWP30P140LVT U7409 ( .A1(i_data_bus[957]), .A2(n7528), .B1(
        i_data_bus[573]), .B2(n7526), .ZN(n6933) );
  ND4D1BWP30P140LVT U7410 ( .A1(n6936), .A2(n6935), .A3(n6934), .A4(n6933), 
        .ZN(n6937) );
  NR4D0BWP30P140LVT U7411 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), 
        .ZN(n6941) );
  ND4D4BWP30P140LVT U7412 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6941), 
        .ZN(o_data_bus[93]) );
  AOI22D1BWP30P140LVT U7413 ( .A1(i_data_bus[380]), .A2(n7495), .B1(
        i_data_bus[444]), .B2(n7523), .ZN(n6964) );
  AOI22D1BWP30P140LVT U7414 ( .A1(i_data_bus[508]), .A2(n7459), .B1(
        i_data_bus[316]), .B2(n7494), .ZN(n6963) );
  AOI22D1BWP30P140LVT U7415 ( .A1(i_data_bus[92]), .A2(n7511), .B1(
        i_data_bus[892]), .B2(n7497), .ZN(n6948) );
  AOI22D1BWP30P140LVT U7416 ( .A1(i_data_bus[764]), .A2(n7504), .B1(
        i_data_bus[860]), .B2(n7498), .ZN(n6947) );
  AOI22D1BWP30P140LVT U7417 ( .A1(i_data_bus[124]), .A2(n7512), .B1(
        i_data_bus[700]), .B2(n7509), .ZN(n6946) );
  AOI22D1BWP30P140LVT U7418 ( .A1(i_data_bus[796]), .A2(n7516), .B1(
        i_data_bus[156]), .B2(n7503), .ZN(n6945) );
  AN4D0BWP30P140LVT U7419 ( .A1(n6948), .A2(n6947), .A3(n6946), .A4(n6945), 
        .Z(n6962) );
  AOI22D1BWP30P140LVT U7420 ( .A1(i_data_bus[60]), .A2(n7514), .B1(
        i_data_bus[252]), .B2(n7501), .ZN(n6952) );
  AOI22D1BWP30P140LVT U7421 ( .A1(i_data_bus[28]), .A2(n7500), .B1(
        i_data_bus[668]), .B2(n7499), .ZN(n6951) );
  AOI22D1BWP30P140LVT U7422 ( .A1(i_data_bus[828]), .A2(n7513), .B1(
        i_data_bus[220]), .B2(n7502), .ZN(n6950) );
  AOI22D1BWP30P140LVT U7423 ( .A1(i_data_bus[732]), .A2(n7510), .B1(
        i_data_bus[188]), .B2(n7515), .ZN(n6949) );
  ND4D1BWP30P140LVT U7424 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(n6949), 
        .ZN(n6960) );
  INVD1BWP30P140LVT U7425 ( .I(i_data_bus[476]), .ZN(n8005) );
  INVD1BWP30P140LVT U7426 ( .I(i_data_bus[284]), .ZN(n8929) );
  OAI22D1BWP30P140LVT U7427 ( .A1(n8005), .A2(n7522), .B1(n8929), .B2(n7521), 
        .ZN(n6959) );
  INVD1BWP30P140LVT U7428 ( .I(i_data_bus[348]), .ZN(n9248) );
  INVD1BWP30P140LVT U7429 ( .I(i_data_bus[412]), .ZN(n9246) );
  OAI22D1BWP30P140LVT U7430 ( .A1(n9248), .A2(n7458), .B1(n9246), .B2(n7411), 
        .ZN(n6958) );
  AOI22D1BWP30P140LVT U7431 ( .A1(i_data_bus[988]), .A2(n7525), .B1(
        i_data_bus[956]), .B2(n7528), .ZN(n6956) );
  AOI22D1BWP30P140LVT U7432 ( .A1(i_data_bus[540]), .A2(n7530), .B1(
        i_data_bus[604]), .B2(n7531), .ZN(n6955) );
  AOI22D1BWP30P140LVT U7433 ( .A1(i_data_bus[924]), .A2(n7527), .B1(
        i_data_bus[1020]), .B2(n7532), .ZN(n6954) );
  AOI22D1BWP30P140LVT U7434 ( .A1(i_data_bus[636]), .A2(n7529), .B1(
        i_data_bus[572]), .B2(n7526), .ZN(n6953) );
  ND4D1BWP30P140LVT U7435 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), 
        .ZN(n6957) );
  NR4D0BWP30P140LVT U7436 ( .A1(n6960), .A2(n6959), .A3(n6958), .A4(n6957), 
        .ZN(n6961) );
  ND4D4BWP30P140LVT U7437 ( .A1(n6964), .A2(n6963), .A3(n6962), .A4(n6961), 
        .ZN(o_data_bus[92]) );
  AOI22D1BWP30P140LVT U7438 ( .A1(i_data_bus[315]), .A2(n7494), .B1(
        i_data_bus[475]), .B2(n7472), .ZN(n6984) );
  AOI22D1BWP30P140LVT U7439 ( .A1(i_data_bus[443]), .A2(n7523), .B1(
        i_data_bus[283]), .B2(n7436), .ZN(n6983) );
  AOI22D1BWP30P140LVT U7440 ( .A1(i_data_bus[891]), .A2(n7497), .B1(
        i_data_bus[859]), .B2(n7498), .ZN(n6968) );
  AOI22D1BWP30P140LVT U7441 ( .A1(i_data_bus[59]), .A2(n7514), .B1(
        i_data_bus[763]), .B2(n7504), .ZN(n6967) );
  AOI22D1BWP30P140LVT U7442 ( .A1(i_data_bus[219]), .A2(n7502), .B1(
        i_data_bus[187]), .B2(n7515), .ZN(n6966) );
  AOI22D1BWP30P140LVT U7443 ( .A1(i_data_bus[667]), .A2(n7499), .B1(
        i_data_bus[699]), .B2(n7509), .ZN(n6965) );
  AN4D0BWP30P140LVT U7444 ( .A1(n6968), .A2(n6967), .A3(n6966), .A4(n6965), 
        .Z(n6982) );
  AOI22D1BWP30P140LVT U7445 ( .A1(i_data_bus[123]), .A2(n7512), .B1(
        i_data_bus[795]), .B2(n7516), .ZN(n6972) );
  AOI22D1BWP30P140LVT U7446 ( .A1(i_data_bus[27]), .A2(n7500), .B1(
        i_data_bus[731]), .B2(n7510), .ZN(n6971) );
  AOI22D1BWP30P140LVT U7447 ( .A1(i_data_bus[91]), .A2(n7511), .B1(
        i_data_bus[251]), .B2(n7501), .ZN(n6970) );
  AOI22D1BWP30P140LVT U7448 ( .A1(i_data_bus[827]), .A2(n7513), .B1(
        i_data_bus[155]), .B2(n7503), .ZN(n6969) );
  ND4D1BWP30P140LVT U7449 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), 
        .ZN(n6980) );
  INVD1BWP30P140LVT U7450 ( .I(i_data_bus[379]), .ZN(n9605) );
  MOAI22D1BWP30P140LVT U7451 ( .A1(n9605), .A2(n7369), .B1(i_data_bus[507]), 
        .B2(n7459), .ZN(n6979) );
  INVD1BWP30P140LVT U7452 ( .I(i_data_bus[347]), .ZN(n7713) );
  MOAI22D1BWP30P140LVT U7453 ( .A1(n7713), .A2(n7458), .B1(i_data_bus[411]), 
        .B2(n7496), .ZN(n6978) );
  AOI22D1BWP30P140LVT U7454 ( .A1(i_data_bus[571]), .A2(n7526), .B1(
        i_data_bus[539]), .B2(n7530), .ZN(n6976) );
  AOI22D1BWP30P140LVT U7455 ( .A1(i_data_bus[987]), .A2(n7525), .B1(
        i_data_bus[603]), .B2(n7531), .ZN(n6975) );
  AOI22D1BWP30P140LVT U7456 ( .A1(i_data_bus[635]), .A2(n7529), .B1(
        i_data_bus[923]), .B2(n7527), .ZN(n6974) );
  AOI22D1BWP30P140LVT U7457 ( .A1(i_data_bus[1019]), .A2(n7532), .B1(
        i_data_bus[955]), .B2(n7528), .ZN(n6973) );
  ND4D1BWP30P140LVT U7458 ( .A1(n6976), .A2(n6975), .A3(n6974), .A4(n6973), 
        .ZN(n6977) );
  NR4D0BWP30P140LVT U7459 ( .A1(n6980), .A2(n6979), .A3(n6978), .A4(n6977), 
        .ZN(n6981) );
  ND4D4BWP30P140LVT U7460 ( .A1(n6984), .A2(n6983), .A3(n6982), .A4(n6981), 
        .ZN(o_data_bus[91]) );
  AOI22D1BWP30P140LVT U7461 ( .A1(i_data_bus[442]), .A2(n7523), .B1(
        i_data_bus[282]), .B2(n7436), .ZN(n7004) );
  AOI22D1BWP30P140LVT U7462 ( .A1(i_data_bus[314]), .A2(n7494), .B1(
        i_data_bus[346]), .B2(n7493), .ZN(n7003) );
  AOI22D1BWP30P140LVT U7463 ( .A1(i_data_bus[250]), .A2(n7501), .B1(
        i_data_bus[666]), .B2(n7499), .ZN(n6988) );
  AOI22D1BWP30P140LVT U7464 ( .A1(i_data_bus[826]), .A2(n7513), .B1(
        i_data_bus[186]), .B2(n7515), .ZN(n6987) );
  AOI22D1BWP30P140LVT U7465 ( .A1(i_data_bus[218]), .A2(n7502), .B1(
        i_data_bus[858]), .B2(n7498), .ZN(n6986) );
  AOI22D1BWP30P140LVT U7466 ( .A1(i_data_bus[698]), .A2(n7509), .B1(
        i_data_bus[762]), .B2(n7504), .ZN(n6985) );
  AN4D0BWP30P140LVT U7467 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), 
        .Z(n7002) );
  AOI22D1BWP30P140LVT U7468 ( .A1(i_data_bus[58]), .A2(n7514), .B1(
        i_data_bus[794]), .B2(n7516), .ZN(n6992) );
  AOI22D1BWP30P140LVT U7469 ( .A1(i_data_bus[26]), .A2(n7500), .B1(
        i_data_bus[154]), .B2(n7503), .ZN(n6991) );
  AOI22D1BWP30P140LVT U7470 ( .A1(i_data_bus[122]), .A2(n7512), .B1(
        i_data_bus[90]), .B2(n7511), .ZN(n6990) );
  AOI22D1BWP30P140LVT U7471 ( .A1(i_data_bus[890]), .A2(n7497), .B1(
        i_data_bus[730]), .B2(n7510), .ZN(n6989) );
  ND4D1BWP30P140LVT U7472 ( .A1(n6992), .A2(n6991), .A3(n6990), .A4(n6989), 
        .ZN(n7000) );
  INVD1BWP30P140LVT U7473 ( .I(i_data_bus[378]), .ZN(n9269) );
  MOAI22D1BWP30P140LVT U7474 ( .A1(n9269), .A2(n7369), .B1(i_data_bus[474]), 
        .B2(n7472), .ZN(n6999) );
  INVD1BWP30P140LVT U7475 ( .I(i_data_bus[506]), .ZN(n9628) );
  INVD1BWP30P140LVT U7476 ( .I(i_data_bus[410]), .ZN(n9627) );
  OAI22D1BWP30P140LVT U7477 ( .A1(n9628), .A2(n7524), .B1(n9627), .B2(n7411), 
        .ZN(n6998) );
  AOI22D1BWP30P140LVT U7478 ( .A1(i_data_bus[602]), .A2(n7531), .B1(
        i_data_bus[954]), .B2(n7528), .ZN(n6996) );
  AOI22D1BWP30P140LVT U7479 ( .A1(i_data_bus[986]), .A2(n7525), .B1(
        i_data_bus[922]), .B2(n7527), .ZN(n6995) );
  AOI22D1BWP30P140LVT U7480 ( .A1(i_data_bus[1018]), .A2(n7532), .B1(
        i_data_bus[570]), .B2(n7526), .ZN(n6994) );
  AOI22D1BWP30P140LVT U7481 ( .A1(i_data_bus[538]), .A2(n7530), .B1(
        i_data_bus[634]), .B2(n7529), .ZN(n6993) );
  ND4D1BWP30P140LVT U7482 ( .A1(n6996), .A2(n6995), .A3(n6994), .A4(n6993), 
        .ZN(n6997) );
  NR4D0BWP30P140LVT U7483 ( .A1(n7000), .A2(n6999), .A3(n6998), .A4(n6997), 
        .ZN(n7001) );
  ND4D4BWP30P140LVT U7484 ( .A1(n7004), .A2(n7003), .A3(n7002), .A4(n7001), 
        .ZN(o_data_bus[90]) );
  AOI22D1BWP30P140LVT U7485 ( .A1(i_data_bus[377]), .A2(n7495), .B1(
        i_data_bus[473]), .B2(n7472), .ZN(n7024) );
  AOI22D1BWP30P140LVT U7486 ( .A1(i_data_bus[345]), .A2(n7493), .B1(
        i_data_bus[313]), .B2(n7494), .ZN(n7023) );
  AOI22D1BWP30P140LVT U7487 ( .A1(i_data_bus[921]), .A2(n7527), .B1(
        i_data_bus[985]), .B2(n7525), .ZN(n7008) );
  AOI22D1BWP30P140LVT U7488 ( .A1(i_data_bus[537]), .A2(n7530), .B1(
        i_data_bus[953]), .B2(n7528), .ZN(n7007) );
  AOI22D1BWP30P140LVT U7489 ( .A1(i_data_bus[1017]), .A2(n7532), .B1(
        i_data_bus[633]), .B2(n7529), .ZN(n7006) );
  AOI22D1BWP30P140LVT U7490 ( .A1(i_data_bus[569]), .A2(n7526), .B1(
        i_data_bus[601]), .B2(n7531), .ZN(n7005) );
  AN4D0BWP30P140LVT U7491 ( .A1(n7008), .A2(n7007), .A3(n7006), .A4(n7005), 
        .Z(n7022) );
  INVD1BWP30P140LVT U7492 ( .I(i_data_bus[409]), .ZN(n8581) );
  MOAI22D1BWP30P140LVT U7493 ( .A1(n8581), .A2(n7411), .B1(i_data_bus[281]), 
        .B2(n7436), .ZN(n7020) );
  INVD1BWP30P140LVT U7494 ( .I(i_data_bus[505]), .ZN(n8761) );
  MOAI22D1BWP30P140LVT U7495 ( .A1(n8761), .A2(n7524), .B1(i_data_bus[441]), 
        .B2(n7523), .ZN(n7019) );
  AOI22D1BWP30P140LVT U7496 ( .A1(i_data_bus[121]), .A2(n7512), .B1(
        i_data_bus[249]), .B2(n7501), .ZN(n7012) );
  AOI22D1BWP30P140LVT U7497 ( .A1(i_data_bus[57]), .A2(n7514), .B1(
        i_data_bus[857]), .B2(n7498), .ZN(n7011) );
  AOI22D1BWP30P140LVT U7498 ( .A1(i_data_bus[153]), .A2(n7503), .B1(
        i_data_bus[889]), .B2(n7497), .ZN(n7010) );
  AOI22D1BWP30P140LVT U7499 ( .A1(i_data_bus[89]), .A2(n7511), .B1(
        i_data_bus[217]), .B2(n7502), .ZN(n7009) );
  ND4D1BWP30P140LVT U7500 ( .A1(n7012), .A2(n7011), .A3(n7010), .A4(n7009), 
        .ZN(n7018) );
  AOI22D1BWP30P140LVT U7501 ( .A1(i_data_bus[729]), .A2(n7510), .B1(
        i_data_bus[793]), .B2(n7516), .ZN(n7016) );
  AOI22D1BWP30P140LVT U7502 ( .A1(i_data_bus[697]), .A2(n7509), .B1(
        i_data_bus[185]), .B2(n7515), .ZN(n7015) );
  AOI22D1BWP30P140LVT U7503 ( .A1(i_data_bus[25]), .A2(n7500), .B1(
        i_data_bus[825]), .B2(n7513), .ZN(n7014) );
  AOI22D1BWP30P140LVT U7504 ( .A1(i_data_bus[665]), .A2(n7499), .B1(
        i_data_bus[761]), .B2(n7504), .ZN(n7013) );
  ND4D1BWP30P140LVT U7505 ( .A1(n7016), .A2(n7015), .A3(n7014), .A4(n7013), 
        .ZN(n7017) );
  NR4D0BWP30P140LVT U7506 ( .A1(n7020), .A2(n7019), .A3(n7018), .A4(n7017), 
        .ZN(n7021) );
  ND4D4BWP30P140LVT U7507 ( .A1(n7024), .A2(n7023), .A3(n7022), .A4(n7021), 
        .ZN(o_data_bus[89]) );
  AOI22D1BWP30P140LVT U7508 ( .A1(i_data_bus[344]), .A2(n7493), .B1(
        i_data_bus[408]), .B2(n7496), .ZN(n7044) );
  AOI22D1BWP30P140LVT U7509 ( .A1(i_data_bus[440]), .A2(n7523), .B1(
        i_data_bus[472]), .B2(n7472), .ZN(n7043) );
  AOI22D1BWP30P140LVT U7510 ( .A1(i_data_bus[696]), .A2(n7509), .B1(
        i_data_bus[760]), .B2(n7504), .ZN(n7028) );
  AOI22D1BWP30P140LVT U7511 ( .A1(i_data_bus[248]), .A2(n7501), .B1(
        i_data_bus[888]), .B2(n7497), .ZN(n7027) );
  AOI22D1BWP30P140LVT U7512 ( .A1(i_data_bus[88]), .A2(n7511), .B1(
        i_data_bus[216]), .B2(n7502), .ZN(n7026) );
  AOI22D1BWP30P140LVT U7513 ( .A1(i_data_bus[824]), .A2(n7513), .B1(
        i_data_bus[184]), .B2(n7515), .ZN(n7025) );
  AN4D0BWP30P140LVT U7514 ( .A1(n7028), .A2(n7027), .A3(n7026), .A4(n7025), 
        .Z(n7042) );
  AOI22D1BWP30P140LVT U7515 ( .A1(i_data_bus[24]), .A2(n7500), .B1(
        i_data_bus[728]), .B2(n7510), .ZN(n7032) );
  AOI22D1BWP30P140LVT U7516 ( .A1(i_data_bus[856]), .A2(n7498), .B1(
        i_data_bus[664]), .B2(n7499), .ZN(n7031) );
  AOI22D1BWP30P140LVT U7517 ( .A1(i_data_bus[120]), .A2(n7512), .B1(
        i_data_bus[56]), .B2(n7514), .ZN(n7030) );
  AOI22D1BWP30P140LVT U7518 ( .A1(i_data_bus[792]), .A2(n7516), .B1(
        i_data_bus[152]), .B2(n7503), .ZN(n7029) );
  ND4D1BWP30P140LVT U7519 ( .A1(n7032), .A2(n7031), .A3(n7030), .A4(n7029), 
        .ZN(n7040) );
  INVD1BWP30P140LVT U7520 ( .I(i_data_bus[504]), .ZN(n8046) );
  MOAI22D1BWP30P140LVT U7521 ( .A1(n8046), .A2(n7524), .B1(i_data_bus[376]), 
        .B2(n7495), .ZN(n7039) );
  INVD1BWP30P140LVT U7522 ( .I(i_data_bus[280]), .ZN(n7857) );
  INVD1BWP30P140LVT U7523 ( .I(i_data_bus[312]), .ZN(n8782) );
  OAI22D1BWP30P140LVT U7524 ( .A1(n7857), .A2(n7521), .B1(n8782), .B2(n7394), 
        .ZN(n7038) );
  AOI22D1BWP30P140LVT U7525 ( .A1(i_data_bus[984]), .A2(n7525), .B1(
        i_data_bus[568]), .B2(n7526), .ZN(n7036) );
  AOI22D1BWP30P140LVT U7526 ( .A1(i_data_bus[1016]), .A2(n7532), .B1(
        i_data_bus[920]), .B2(n7527), .ZN(n7035) );
  AOI22D1BWP30P140LVT U7527 ( .A1(i_data_bus[632]), .A2(n7529), .B1(
        i_data_bus[536]), .B2(n7530), .ZN(n7034) );
  AOI22D1BWP30P140LVT U7528 ( .A1(i_data_bus[600]), .A2(n7531), .B1(
        i_data_bus[952]), .B2(n7528), .ZN(n7033) );
  ND4D1BWP30P140LVT U7529 ( .A1(n7036), .A2(n7035), .A3(n7034), .A4(n7033), 
        .ZN(n7037) );
  NR4D0BWP30P140LVT U7530 ( .A1(n7040), .A2(n7039), .A3(n7038), .A4(n7037), 
        .ZN(n7041) );
  ND4D4BWP30P140LVT U7531 ( .A1(n7044), .A2(n7043), .A3(n7042), .A4(n7041), 
        .ZN(o_data_bus[88]) );
  AOI22D1BWP30P140LVT U7532 ( .A1(i_data_bus[503]), .A2(n7459), .B1(
        i_data_bus[343]), .B2(n7493), .ZN(n7064) );
  AOI22D1BWP30P140LVT U7533 ( .A1(i_data_bus[311]), .A2(n7494), .B1(
        i_data_bus[407]), .B2(n7496), .ZN(n7063) );
  AOI22D1BWP30P140LVT U7534 ( .A1(i_data_bus[183]), .A2(n7515), .B1(
        i_data_bus[151]), .B2(n7503), .ZN(n7048) );
  AOI22D1BWP30P140LVT U7535 ( .A1(i_data_bus[55]), .A2(n7514), .B1(
        i_data_bus[727]), .B2(n7510), .ZN(n7047) );
  AOI22D1BWP30P140LVT U7536 ( .A1(i_data_bus[759]), .A2(n7504), .B1(
        i_data_bus[663]), .B2(n7499), .ZN(n7046) );
  AOI22D1BWP30P140LVT U7537 ( .A1(i_data_bus[23]), .A2(n7500), .B1(
        i_data_bus[823]), .B2(n7513), .ZN(n7045) );
  AN4D0BWP30P140LVT U7538 ( .A1(n7048), .A2(n7047), .A3(n7046), .A4(n7045), 
        .Z(n7062) );
  AOI22D1BWP30P140LVT U7539 ( .A1(i_data_bus[87]), .A2(n7511), .B1(
        i_data_bus[119]), .B2(n7512), .ZN(n7052) );
  AOI22D1BWP30P140LVT U7540 ( .A1(i_data_bus[695]), .A2(n7509), .B1(
        i_data_bus[791]), .B2(n7516), .ZN(n7051) );
  AOI22D1BWP30P140LVT U7541 ( .A1(i_data_bus[247]), .A2(n7501), .B1(
        i_data_bus[215]), .B2(n7502), .ZN(n7050) );
  AOI22D1BWP30P140LVT U7542 ( .A1(i_data_bus[887]), .A2(n7497), .B1(
        i_data_bus[855]), .B2(n7498), .ZN(n7049) );
  ND4D1BWP30P140LVT U7543 ( .A1(n7052), .A2(n7051), .A3(n7050), .A4(n7049), 
        .ZN(n7060) );
  INVD1BWP30P140LVT U7544 ( .I(i_data_bus[471]), .ZN(n8950) );
  INVD1BWP30P140LVT U7545 ( .I(i_data_bus[375]), .ZN(n9290) );
  OAI22D1BWP30P140LVT U7546 ( .A1(n8950), .A2(n7522), .B1(n9290), .B2(n7369), 
        .ZN(n7059) );
  INVD1BWP30P140LVT U7547 ( .I(i_data_bus[439]), .ZN(n9291) );
  MOAI22D1BWP30P140LVT U7548 ( .A1(n9291), .A2(n7437), .B1(i_data_bus[279]), 
        .B2(n7436), .ZN(n7058) );
  AOI22D1BWP30P140LVT U7549 ( .A1(i_data_bus[1015]), .A2(n7532), .B1(
        i_data_bus[567]), .B2(n7526), .ZN(n7056) );
  AOI22D1BWP30P140LVT U7550 ( .A1(i_data_bus[631]), .A2(n7529), .B1(
        i_data_bus[919]), .B2(n7527), .ZN(n7055) );
  AOI22D1BWP30P140LVT U7551 ( .A1(i_data_bus[983]), .A2(n7525), .B1(
        i_data_bus[535]), .B2(n7530), .ZN(n7054) );
  AOI22D1BWP30P140LVT U7552 ( .A1(i_data_bus[599]), .A2(n7531), .B1(
        i_data_bus[951]), .B2(n7528), .ZN(n7053) );
  ND4D1BWP30P140LVT U7553 ( .A1(n7056), .A2(n7055), .A3(n7054), .A4(n7053), 
        .ZN(n7057) );
  NR4D0BWP30P140LVT U7554 ( .A1(n7060), .A2(n7059), .A3(n7058), .A4(n7057), 
        .ZN(n7061) );
  ND4D4BWP30P140LVT U7555 ( .A1(n7064), .A2(n7063), .A3(n7062), .A4(n7061), 
        .ZN(o_data_bus[87]) );
  AOI22D1BWP30P140LVT U7556 ( .A1(i_data_bus[438]), .A2(n7523), .B1(
        i_data_bus[502]), .B2(n7459), .ZN(n7084) );
  AOI22D1BWP30P140LVT U7557 ( .A1(i_data_bus[310]), .A2(n7494), .B1(
        i_data_bus[278]), .B2(n7436), .ZN(n7083) );
  AOI22D1BWP30P140LVT U7558 ( .A1(i_data_bus[822]), .A2(n7513), .B1(
        i_data_bus[246]), .B2(n7501), .ZN(n7068) );
  AOI22D1BWP30P140LVT U7559 ( .A1(i_data_bus[118]), .A2(n7512), .B1(
        i_data_bus[86]), .B2(n7511), .ZN(n7067) );
  AOI22D1BWP30P140LVT U7560 ( .A1(i_data_bus[758]), .A2(n7504), .B1(
        i_data_bus[886]), .B2(n7497), .ZN(n7066) );
  AOI22D1BWP30P140LVT U7561 ( .A1(i_data_bus[182]), .A2(n7515), .B1(
        i_data_bus[214]), .B2(n7502), .ZN(n7065) );
  AN4D0BWP30P140LVT U7562 ( .A1(n7068), .A2(n7067), .A3(n7066), .A4(n7065), 
        .Z(n7082) );
  AOI22D1BWP30P140LVT U7563 ( .A1(i_data_bus[22]), .A2(n7500), .B1(
        i_data_bus[662]), .B2(n7499), .ZN(n7072) );
  AOI22D1BWP30P140LVT U7564 ( .A1(i_data_bus[54]), .A2(n7514), .B1(
        i_data_bus[150]), .B2(n7503), .ZN(n7071) );
  AOI22D1BWP30P140LVT U7565 ( .A1(i_data_bus[694]), .A2(n7509), .B1(
        i_data_bus[726]), .B2(n7510), .ZN(n7070) );
  AOI22D1BWP30P140LVT U7566 ( .A1(i_data_bus[790]), .A2(n7516), .B1(
        i_data_bus[854]), .B2(n7498), .ZN(n7069) );
  ND4D1BWP30P140LVT U7567 ( .A1(n7072), .A2(n7071), .A3(n7070), .A4(n7069), 
        .ZN(n7080) );
  INVD1BWP30P140LVT U7568 ( .I(i_data_bus[470]), .ZN(n8804) );
  MOAI22D1BWP30P140LVT U7569 ( .A1(n8804), .A2(n7522), .B1(i_data_bus[374]), 
        .B2(n7495), .ZN(n7079) );
  INVD1BWP30P140LVT U7570 ( .I(i_data_bus[342]), .ZN(n8803) );
  MOAI22D1BWP30P140LVT U7571 ( .A1(n8803), .A2(n7458), .B1(i_data_bus[406]), 
        .B2(n7496), .ZN(n7078) );
  AOI22D1BWP30P140LVT U7572 ( .A1(i_data_bus[534]), .A2(n7530), .B1(
        i_data_bus[918]), .B2(n7527), .ZN(n7076) );
  AOI22D1BWP30P140LVT U7573 ( .A1(i_data_bus[566]), .A2(n7526), .B1(
        i_data_bus[982]), .B2(n7525), .ZN(n7075) );
  AOI22D1BWP30P140LVT U7574 ( .A1(i_data_bus[1014]), .A2(n7532), .B1(
        i_data_bus[598]), .B2(n7531), .ZN(n7074) );
  AOI22D1BWP30P140LVT U7575 ( .A1(i_data_bus[950]), .A2(n7528), .B1(
        i_data_bus[630]), .B2(n7529), .ZN(n7073) );
  ND4D1BWP30P140LVT U7576 ( .A1(n7076), .A2(n7075), .A3(n7074), .A4(n7073), 
        .ZN(n7077) );
  NR4D0BWP30P140LVT U7577 ( .A1(n7080), .A2(n7079), .A3(n7078), .A4(n7077), 
        .ZN(n7081) );
  ND4D4BWP30P140LVT U7578 ( .A1(n7084), .A2(n7083), .A3(n7082), .A4(n7081), 
        .ZN(o_data_bus[86]) );
  AOI22D1BWP30P140LVT U7579 ( .A1(i_data_bus[339]), .A2(n7493), .B1(
        i_data_bus[435]), .B2(n7523), .ZN(n7104) );
  AOI22D1BWP30P140LVT U7580 ( .A1(i_data_bus[371]), .A2(n7495), .B1(
        i_data_bus[403]), .B2(n7496), .ZN(n7103) );
  AOI22D1BWP30P140LVT U7581 ( .A1(i_data_bus[243]), .A2(n7501), .B1(
        i_data_bus[659]), .B2(n7499), .ZN(n7088) );
  AOI22D1BWP30P140LVT U7582 ( .A1(i_data_bus[19]), .A2(n7500), .B1(
        i_data_bus[883]), .B2(n7497), .ZN(n7087) );
  AOI22D1BWP30P140LVT U7583 ( .A1(i_data_bus[179]), .A2(n7515), .B1(
        i_data_bus[851]), .B2(n7498), .ZN(n7086) );
  AOI22D1BWP30P140LVT U7584 ( .A1(i_data_bus[211]), .A2(n7502), .B1(
        i_data_bus[787]), .B2(n7516), .ZN(n7085) );
  AN4D0BWP30P140LVT U7585 ( .A1(n7088), .A2(n7087), .A3(n7086), .A4(n7085), 
        .Z(n7102) );
  AOI22D1BWP30P140LVT U7586 ( .A1(i_data_bus[83]), .A2(n7511), .B1(
        i_data_bus[691]), .B2(n7509), .ZN(n7092) );
  AOI22D1BWP30P140LVT U7587 ( .A1(i_data_bus[115]), .A2(n7512), .B1(
        i_data_bus[755]), .B2(n7504), .ZN(n7091) );
  AOI22D1BWP30P140LVT U7588 ( .A1(i_data_bus[147]), .A2(n7503), .B1(
        i_data_bus[819]), .B2(n7513), .ZN(n7090) );
  AOI22D1BWP30P140LVT U7589 ( .A1(i_data_bus[51]), .A2(n7514), .B1(
        i_data_bus[723]), .B2(n7510), .ZN(n7089) );
  ND4D1BWP30P140LVT U7590 ( .A1(n7092), .A2(n7091), .A3(n7090), .A4(n7089), 
        .ZN(n7100) );
  INVD1BWP30P140LVT U7591 ( .I(i_data_bus[499]), .ZN(n7878) );
  MOAI22D1BWP30P140LVT U7592 ( .A1(n7878), .A2(n7524), .B1(i_data_bus[275]), 
        .B2(n7436), .ZN(n7099) );
  INVD1BWP30P140LVT U7593 ( .I(i_data_bus[307]), .ZN(n8433) );
  MOAI22D1BWP30P140LVT U7594 ( .A1(n8433), .A2(n7394), .B1(i_data_bus[467]), 
        .B2(n7472), .ZN(n7098) );
  AOI22D1BWP30P140LVT U7595 ( .A1(i_data_bus[627]), .A2(n7529), .B1(
        i_data_bus[595]), .B2(n7531), .ZN(n7096) );
  AOI22D1BWP30P140LVT U7596 ( .A1(i_data_bus[531]), .A2(n7530), .B1(
        i_data_bus[947]), .B2(n7528), .ZN(n7095) );
  AOI22D1BWP30P140LVT U7597 ( .A1(i_data_bus[979]), .A2(n7525), .B1(
        i_data_bus[1011]), .B2(n7532), .ZN(n7094) );
  AOI22D1BWP30P140LVT U7598 ( .A1(i_data_bus[563]), .A2(n7526), .B1(
        i_data_bus[915]), .B2(n7527), .ZN(n7093) );
  ND4D1BWP30P140LVT U7599 ( .A1(n7096), .A2(n7095), .A3(n7094), .A4(n7093), 
        .ZN(n7097) );
  NR4D0BWP30P140LVT U7600 ( .A1(n7100), .A2(n7099), .A3(n7098), .A4(n7097), 
        .ZN(n7101) );
  ND4D4BWP30P140LVT U7601 ( .A1(n7104), .A2(n7103), .A3(n7102), .A4(n7101), 
        .ZN(o_data_bus[83]) );
  AOI22D1BWP30P140LVT U7602 ( .A1(i_data_bus[498]), .A2(n7459), .B1(
        i_data_bus[306]), .B2(n7494), .ZN(n7124) );
  AOI22D1BWP30P140LVT U7603 ( .A1(i_data_bus[274]), .A2(n7436), .B1(
        i_data_bus[434]), .B2(n7523), .ZN(n7123) );
  AOI22D1BWP30P140LVT U7604 ( .A1(i_data_bus[18]), .A2(n7500), .B1(
        i_data_bus[690]), .B2(n7509), .ZN(n7108) );
  AOI22D1BWP30P140LVT U7605 ( .A1(i_data_bus[50]), .A2(n7514), .B1(
        i_data_bus[850]), .B2(n7498), .ZN(n7107) );
  AOI22D1BWP30P140LVT U7606 ( .A1(i_data_bus[82]), .A2(n7511), .B1(
        i_data_bus[754]), .B2(n7504), .ZN(n7106) );
  AOI22D1BWP30P140LVT U7607 ( .A1(i_data_bus[146]), .A2(n7503), .B1(
        i_data_bus[786]), .B2(n7516), .ZN(n7105) );
  AN4D0BWP30P140LVT U7608 ( .A1(n7108), .A2(n7107), .A3(n7106), .A4(n7105), 
        .Z(n7122) );
  AOI22D1BWP30P140LVT U7609 ( .A1(i_data_bus[402]), .A2(n7496), .B1(
        i_data_bus[370]), .B2(n7495), .ZN(n7120) );
  AO22D1BWP30P140LVT U7610 ( .A1(i_data_bus[466]), .A2(n7472), .B1(
        i_data_bus[338]), .B2(n7493), .Z(n7119) );
  AOI22D1BWP30P140LVT U7611 ( .A1(i_data_bus[242]), .A2(n7501), .B1(
        i_data_bus[178]), .B2(n7515), .ZN(n7112) );
  AOI22D1BWP30P140LVT U7612 ( .A1(i_data_bus[722]), .A2(n7510), .B1(
        i_data_bus[210]), .B2(n7502), .ZN(n7111) );
  AOI22D1BWP30P140LVT U7613 ( .A1(i_data_bus[818]), .A2(n7513), .B1(
        i_data_bus[658]), .B2(n7499), .ZN(n7110) );
  AOI22D1BWP30P140LVT U7614 ( .A1(i_data_bus[114]), .A2(n7512), .B1(
        i_data_bus[882]), .B2(n7497), .ZN(n7109) );
  ND4D1BWP30P140LVT U7615 ( .A1(n7112), .A2(n7111), .A3(n7110), .A4(n7109), 
        .ZN(n7118) );
  AOI22D1BWP30P140LVT U7616 ( .A1(i_data_bus[594]), .A2(n7531), .B1(
        i_data_bus[530]), .B2(n7530), .ZN(n7116) );
  AOI22D1BWP30P140LVT U7617 ( .A1(i_data_bus[562]), .A2(n7526), .B1(
        i_data_bus[946]), .B2(n7528), .ZN(n7115) );
  AOI22D1BWP30P140LVT U7618 ( .A1(i_data_bus[626]), .A2(n7529), .B1(
        i_data_bus[978]), .B2(n7525), .ZN(n7114) );
  AOI22D1BWP30P140LVT U7619 ( .A1(i_data_bus[1010]), .A2(n7532), .B1(
        i_data_bus[914]), .B2(n7527), .ZN(n7113) );
  ND4D1BWP30P140LVT U7620 ( .A1(n7116), .A2(n7115), .A3(n7114), .A4(n7113), 
        .ZN(n7117) );
  INR4D0BWP30P140LVT U7621 ( .A1(n7120), .B1(n7119), .B2(n7118), .B3(n7117), 
        .ZN(n7121) );
  ND4D4BWP30P140LVT U7622 ( .A1(n7124), .A2(n7123), .A3(n7122), .A4(n7121), 
        .ZN(o_data_bus[82]) );
  AOI22D1BWP30P140LVT U7623 ( .A1(i_data_bus[462]), .A2(n7472), .B1(
        i_data_bus[334]), .B2(n7493), .ZN(n7144) );
  AOI22D1BWP30P140LVT U7624 ( .A1(i_data_bus[270]), .A2(n7436), .B1(
        i_data_bus[302]), .B2(n7494), .ZN(n7143) );
  AOI22D1BWP30P140LVT U7625 ( .A1(i_data_bus[206]), .A2(n7502), .B1(
        i_data_bus[814]), .B2(n7513), .ZN(n7128) );
  AOI22D1BWP30P140LVT U7626 ( .A1(i_data_bus[238]), .A2(n7501), .B1(
        i_data_bus[654]), .B2(n7499), .ZN(n7127) );
  AOI22D1BWP30P140LVT U7627 ( .A1(i_data_bus[46]), .A2(n7514), .B1(
        i_data_bus[782]), .B2(n7516), .ZN(n7126) );
  AOI22D1BWP30P140LVT U7628 ( .A1(i_data_bus[14]), .A2(n7500), .B1(
        i_data_bus[718]), .B2(n7510), .ZN(n7125) );
  AN4D0BWP30P140LVT U7629 ( .A1(n7128), .A2(n7127), .A3(n7126), .A4(n7125), 
        .Z(n7142) );
  AOI22D1BWP30P140LVT U7630 ( .A1(i_data_bus[110]), .A2(n7512), .B1(
        i_data_bus[174]), .B2(n7515), .ZN(n7132) );
  AOI22D1BWP30P140LVT U7631 ( .A1(i_data_bus[78]), .A2(n7511), .B1(
        i_data_bus[750]), .B2(n7504), .ZN(n7131) );
  AOI22D1BWP30P140LVT U7632 ( .A1(i_data_bus[142]), .A2(n7503), .B1(
        i_data_bus[846]), .B2(n7498), .ZN(n7130) );
  AOI22D1BWP30P140LVT U7633 ( .A1(i_data_bus[878]), .A2(n7497), .B1(
        i_data_bus[686]), .B2(n7509), .ZN(n7129) );
  ND4D1BWP30P140LVT U7634 ( .A1(n7132), .A2(n7131), .A3(n7130), .A4(n7129), 
        .ZN(n7140) );
  INVD1BWP30P140LVT U7635 ( .I(i_data_bus[398]), .ZN(n8251) );
  MOAI22D1BWP30P140LVT U7636 ( .A1(n8251), .A2(n7411), .B1(i_data_bus[430]), 
        .B2(n7523), .ZN(n7139) );
  INVD1BWP30P140LVT U7637 ( .I(i_data_bus[494]), .ZN(n9398) );
  MOAI22D1BWP30P140LVT U7638 ( .A1(n9398), .A2(n7524), .B1(i_data_bus[366]), 
        .B2(n7495), .ZN(n7138) );
  AOI22D1BWP30P140LVT U7639 ( .A1(i_data_bus[974]), .A2(n7525), .B1(
        i_data_bus[942]), .B2(n7528), .ZN(n7136) );
  AOI22D1BWP30P140LVT U7640 ( .A1(i_data_bus[1006]), .A2(n7532), .B1(
        i_data_bus[558]), .B2(n7526), .ZN(n7135) );
  AOI22D1BWP30P140LVT U7641 ( .A1(i_data_bus[910]), .A2(n7527), .B1(
        i_data_bus[590]), .B2(n7531), .ZN(n7134) );
  AOI22D1BWP30P140LVT U7642 ( .A1(i_data_bus[622]), .A2(n7529), .B1(
        i_data_bus[526]), .B2(n7530), .ZN(n7133) );
  ND4D1BWP30P140LVT U7643 ( .A1(n7136), .A2(n7135), .A3(n7134), .A4(n7133), 
        .ZN(n7137) );
  NR4D0BWP30P140LVT U7644 ( .A1(n7140), .A2(n7139), .A3(n7138), .A4(n7137), 
        .ZN(n7141) );
  ND4D4BWP30P140LVT U7645 ( .A1(n7144), .A2(n7143), .A3(n7142), .A4(n7141), 
        .ZN(o_data_bus[78]) );
  AOI22D1BWP30P140LVT U7646 ( .A1(i_data_bus[268]), .A2(n7436), .B1(
        i_data_bus[332]), .B2(n7493), .ZN(n7164) );
  AOI22D1BWP30P140LVT U7647 ( .A1(i_data_bus[300]), .A2(n7494), .B1(
        i_data_bus[396]), .B2(n7496), .ZN(n7163) );
  AOI22D1BWP30P140LVT U7648 ( .A1(i_data_bus[76]), .A2(n7511), .B1(
        i_data_bus[844]), .B2(n7498), .ZN(n7148) );
  AOI22D1BWP30P140LVT U7649 ( .A1(i_data_bus[716]), .A2(n7510), .B1(
        i_data_bus[204]), .B2(n7502), .ZN(n7147) );
  AOI22D1BWP30P140LVT U7650 ( .A1(i_data_bus[684]), .A2(n7509), .B1(
        i_data_bus[236]), .B2(n7501), .ZN(n7146) );
  AOI22D1BWP30P140LVT U7651 ( .A1(i_data_bus[12]), .A2(n7500), .B1(
        i_data_bus[172]), .B2(n7515), .ZN(n7145) );
  AN4D0BWP30P140LVT U7652 ( .A1(n7148), .A2(n7147), .A3(n7146), .A4(n7145), 
        .Z(n7162) );
  AOI22D1BWP30P140LVT U7653 ( .A1(i_data_bus[364]), .A2(n7495), .B1(
        i_data_bus[428]), .B2(n7523), .ZN(n7160) );
  AOI22D1BWP30P140LVT U7654 ( .A1(i_data_bus[44]), .A2(n7514), .B1(
        i_data_bus[108]), .B2(n7512), .ZN(n7152) );
  AOI22D1BWP30P140LVT U7655 ( .A1(i_data_bus[812]), .A2(n7513), .B1(
        i_data_bus[876]), .B2(n7497), .ZN(n7151) );
  AOI22D1BWP30P140LVT U7656 ( .A1(i_data_bus[780]), .A2(n7516), .B1(
        i_data_bus[748]), .B2(n7504), .ZN(n7150) );
  AOI22D1BWP30P140LVT U7657 ( .A1(i_data_bus[140]), .A2(n7503), .B1(
        i_data_bus[652]), .B2(n7499), .ZN(n7149) );
  ND4D1BWP30P140LVT U7658 ( .A1(n7152), .A2(n7151), .A3(n7150), .A4(n7149), 
        .ZN(n7159) );
  INVD1BWP30P140LVT U7659 ( .I(i_data_bus[460]), .ZN(n8972) );
  INVD1BWP30P140LVT U7660 ( .I(i_data_bus[492]), .ZN(n8971) );
  OAI22D1BWP30P140LVT U7661 ( .A1(n8972), .A2(n7522), .B1(n8971), .B2(n7524), 
        .ZN(n7158) );
  AOI22D1BWP30P140LVT U7662 ( .A1(i_data_bus[940]), .A2(n7528), .B1(
        i_data_bus[972]), .B2(n7525), .ZN(n7156) );
  AOI22D1BWP30P140LVT U7663 ( .A1(i_data_bus[620]), .A2(n7529), .B1(
        i_data_bus[588]), .B2(n7531), .ZN(n7155) );
  AOI22D1BWP30P140LVT U7664 ( .A1(i_data_bus[908]), .A2(n7527), .B1(
        i_data_bus[1004]), .B2(n7532), .ZN(n7154) );
  AOI22D1BWP30P140LVT U7665 ( .A1(i_data_bus[556]), .A2(n7526), .B1(
        i_data_bus[524]), .B2(n7530), .ZN(n7153) );
  ND4D1BWP30P140LVT U7666 ( .A1(n7156), .A2(n7155), .A3(n7154), .A4(n7153), 
        .ZN(n7157) );
  INR4D0BWP30P140LVT U7667 ( .A1(n7160), .B1(n7159), .B2(n7158), .B3(n7157), 
        .ZN(n7161) );
  ND4D4BWP30P140LVT U7668 ( .A1(n7164), .A2(n7163), .A3(n7162), .A4(n7161), 
        .ZN(o_data_bus[76]) );
  AOI22D1BWP30P140LVT U7669 ( .A1(i_data_bus[437]), .A2(n7523), .B1(
        i_data_bus[501]), .B2(n7459), .ZN(n7184) );
  AOI22D1BWP30P140LVT U7670 ( .A1(i_data_bus[341]), .A2(n7493), .B1(
        i_data_bus[277]), .B2(n7436), .ZN(n7183) );
  AOI22D1BWP30P140LVT U7671 ( .A1(i_data_bus[981]), .A2(n7525), .B1(
        i_data_bus[1013]), .B2(n7532), .ZN(n7168) );
  AOI22D1BWP30P140LVT U7672 ( .A1(i_data_bus[949]), .A2(n7528), .B1(
        i_data_bus[917]), .B2(n7527), .ZN(n7167) );
  AOI22D1BWP30P140LVT U7673 ( .A1(i_data_bus[629]), .A2(n7529), .B1(
        i_data_bus[565]), .B2(n7526), .ZN(n7166) );
  AOI22D1BWP30P140LVT U7674 ( .A1(i_data_bus[597]), .A2(n7531), .B1(
        i_data_bus[533]), .B2(n7530), .ZN(n7165) );
  AN4D0BWP30P140LVT U7675 ( .A1(n7168), .A2(n7167), .A3(n7166), .A4(n7165), 
        .Z(n7182) );
  INVD1BWP30P140LVT U7676 ( .I(i_data_bus[373]), .ZN(n9312) );
  MOAI22D1BWP30P140LVT U7677 ( .A1(n9312), .A2(n7369), .B1(i_data_bus[469]), 
        .B2(n7472), .ZN(n7180) );
  INVD1BWP30P140LVT U7678 ( .I(i_data_bus[309]), .ZN(n8412) );
  INVD1BWP30P140LVT U7679 ( .I(i_data_bus[405]), .ZN(n8107) );
  OAI22D1BWP30P140LVT U7680 ( .A1(n8412), .A2(n7394), .B1(n8107), .B2(n7411), 
        .ZN(n7179) );
  AOI22D1BWP30P140LVT U7681 ( .A1(i_data_bus[821]), .A2(n7513), .B1(
        i_data_bus[725]), .B2(n7510), .ZN(n7172) );
  AOI22D1BWP30P140LVT U7682 ( .A1(i_data_bus[181]), .A2(n7515), .B1(
        i_data_bus[213]), .B2(n7502), .ZN(n7171) );
  AOI22D1BWP30P140LVT U7683 ( .A1(i_data_bus[21]), .A2(n7500), .B1(
        i_data_bus[149]), .B2(n7503), .ZN(n7170) );
  AOI22D1BWP30P140LVT U7684 ( .A1(i_data_bus[853]), .A2(n7498), .B1(
        i_data_bus[789]), .B2(n7516), .ZN(n7169) );
  ND4D1BWP30P140LVT U7685 ( .A1(n7172), .A2(n7171), .A3(n7170), .A4(n7169), 
        .ZN(n7178) );
  AOI22D1BWP30P140LVT U7686 ( .A1(i_data_bus[117]), .A2(n7512), .B1(
        i_data_bus[693]), .B2(n7509), .ZN(n7176) );
  AOI22D1BWP30P140LVT U7687 ( .A1(i_data_bus[757]), .A2(n7504), .B1(
        i_data_bus[885]), .B2(n7497), .ZN(n7175) );
  AOI22D1BWP30P140LVT U7688 ( .A1(i_data_bus[85]), .A2(n7511), .B1(
        i_data_bus[661]), .B2(n7499), .ZN(n7174) );
  AOI22D1BWP30P140LVT U7689 ( .A1(i_data_bus[53]), .A2(n7514), .B1(
        i_data_bus[245]), .B2(n7501), .ZN(n7173) );
  ND4D1BWP30P140LVT U7690 ( .A1(n7176), .A2(n7175), .A3(n7174), .A4(n7173), 
        .ZN(n7177) );
  NR4D0BWP30P140LVT U7691 ( .A1(n7180), .A2(n7179), .A3(n7178), .A4(n7177), 
        .ZN(n7181) );
  ND4D4BWP30P140LVT U7692 ( .A1(n7184), .A2(n7183), .A3(n7182), .A4(n7181), 
        .ZN(o_data_bus[85]) );
  AOI22D1BWP30P140LVT U7693 ( .A1(i_data_bus[304]), .A2(n7494), .B1(
        i_data_bus[368]), .B2(n7495), .ZN(n7204) );
  AOI22D1BWP30P140LVT U7694 ( .A1(i_data_bus[336]), .A2(n7493), .B1(
        i_data_bus[464]), .B2(n7472), .ZN(n7203) );
  AOI22D1BWP30P140LVT U7695 ( .A1(i_data_bus[528]), .A2(n7530), .B1(
        i_data_bus[912]), .B2(n7527), .ZN(n7188) );
  AOI22D1BWP30P140LVT U7696 ( .A1(i_data_bus[624]), .A2(n7529), .B1(
        i_data_bus[976]), .B2(n7525), .ZN(n7187) );
  AOI22D1BWP30P140LVT U7697 ( .A1(i_data_bus[944]), .A2(n7528), .B1(
        i_data_bus[592]), .B2(n7531), .ZN(n7186) );
  AOI22D1BWP30P140LVT U7698 ( .A1(i_data_bus[560]), .A2(n7526), .B1(
        i_data_bus[1008]), .B2(n7532), .ZN(n7185) );
  AN4D0BWP30P140LVT U7699 ( .A1(n7188), .A2(n7187), .A3(n7186), .A4(n7185), 
        .Z(n7202) );
  INVD1BWP30P140LVT U7700 ( .I(i_data_bus[496]), .ZN(n8209) );
  MOAI22D1BWP30P140LVT U7701 ( .A1(n8209), .A2(n7524), .B1(i_data_bus[272]), 
        .B2(n7436), .ZN(n7200) );
  INVD1BWP30P140LVT U7702 ( .I(i_data_bus[400]), .ZN(n7899) );
  MOAI22D1BWP30P140LVT U7703 ( .A1(n7899), .A2(n7411), .B1(i_data_bus[432]), 
        .B2(n7523), .ZN(n7199) );
  AOI22D1BWP30P140LVT U7704 ( .A1(i_data_bus[16]), .A2(n7500), .B1(
        i_data_bus[144]), .B2(n7503), .ZN(n7192) );
  AOI22D1BWP30P140LVT U7705 ( .A1(i_data_bus[752]), .A2(n7504), .B1(
        i_data_bus[816]), .B2(n7513), .ZN(n7191) );
  AOI22D1BWP30P140LVT U7706 ( .A1(i_data_bus[784]), .A2(n7516), .B1(
        i_data_bus[656]), .B2(n7499), .ZN(n7190) );
  AOI22D1BWP30P140LVT U7707 ( .A1(i_data_bus[880]), .A2(n7497), .B1(
        i_data_bus[688]), .B2(n7509), .ZN(n7189) );
  ND4D1BWP30P140LVT U7708 ( .A1(n7192), .A2(n7191), .A3(n7190), .A4(n7189), 
        .ZN(n7198) );
  AOI22D1BWP30P140LVT U7709 ( .A1(i_data_bus[80]), .A2(n7511), .B1(
        i_data_bus[848]), .B2(n7498), .ZN(n7196) );
  AOI22D1BWP30P140LVT U7710 ( .A1(i_data_bus[112]), .A2(n7512), .B1(
        i_data_bus[176]), .B2(n7515), .ZN(n7195) );
  AOI22D1BWP30P140LVT U7711 ( .A1(i_data_bus[48]), .A2(n7514), .B1(
        i_data_bus[720]), .B2(n7510), .ZN(n7194) );
  AOI22D1BWP30P140LVT U7712 ( .A1(i_data_bus[208]), .A2(n7502), .B1(
        i_data_bus[240]), .B2(n7501), .ZN(n7193) );
  ND4D1BWP30P140LVT U7713 ( .A1(n7196), .A2(n7195), .A3(n7194), .A4(n7193), 
        .ZN(n7197) );
  NR4D0BWP30P140LVT U7714 ( .A1(n7200), .A2(n7199), .A3(n7198), .A4(n7197), 
        .ZN(n7201) );
  ND4D4BWP30P140LVT U7715 ( .A1(n7204), .A2(n7203), .A3(n7202), .A4(n7201), 
        .ZN(o_data_bus[80]) );
  AOI22D1BWP30P140LVT U7716 ( .A1(i_data_bus[491]), .A2(n7459), .B1(
        i_data_bus[427]), .B2(n7523), .ZN(n7224) );
  AOI22D1BWP30P140LVT U7717 ( .A1(i_data_bus[363]), .A2(n7495), .B1(
        i_data_bus[299]), .B2(n7494), .ZN(n7223) );
  AOI22D1BWP30P140LVT U7718 ( .A1(i_data_bus[139]), .A2(n7503), .B1(
        i_data_bus[683]), .B2(n7509), .ZN(n7208) );
  AOI22D1BWP30P140LVT U7719 ( .A1(i_data_bus[75]), .A2(n7511), .B1(
        i_data_bus[171]), .B2(n7515), .ZN(n7207) );
  AOI22D1BWP30P140LVT U7720 ( .A1(i_data_bus[747]), .A2(n7504), .B1(
        i_data_bus[779]), .B2(n7516), .ZN(n7206) );
  AOI22D1BWP30P140LVT U7721 ( .A1(i_data_bus[11]), .A2(n7500), .B1(
        i_data_bus[107]), .B2(n7512), .ZN(n7205) );
  AN4D0BWP30P140LVT U7722 ( .A1(n7208), .A2(n7207), .A3(n7206), .A4(n7205), 
        .Z(n7222) );
  AOI22D1BWP30P140LVT U7723 ( .A1(i_data_bus[395]), .A2(n7496), .B1(
        i_data_bus[267]), .B2(n7436), .ZN(n7220) );
  AOI22D1BWP30P140LVT U7724 ( .A1(i_data_bus[651]), .A2(n7499), .B1(
        i_data_bus[715]), .B2(n7510), .ZN(n7212) );
  AOI22D1BWP30P140LVT U7725 ( .A1(i_data_bus[203]), .A2(n7502), .B1(
        i_data_bus[875]), .B2(n7497), .ZN(n7211) );
  AOI22D1BWP30P140LVT U7726 ( .A1(i_data_bus[43]), .A2(n7514), .B1(
        i_data_bus[811]), .B2(n7513), .ZN(n7210) );
  AOI22D1BWP30P140LVT U7727 ( .A1(i_data_bus[843]), .A2(n7498), .B1(
        i_data_bus[235]), .B2(n7501), .ZN(n7209) );
  ND4D1BWP30P140LVT U7728 ( .A1(n7212), .A2(n7211), .A3(n7210), .A4(n7209), 
        .ZN(n7219) );
  INVD1BWP30P140LVT U7729 ( .I(i_data_bus[459]), .ZN(n9650) );
  INVD1BWP30P140LVT U7730 ( .I(i_data_bus[331]), .ZN(n8514) );
  OAI22D1BWP30P140LVT U7731 ( .A1(n9650), .A2(n7522), .B1(n8514), .B2(n7458), 
        .ZN(n7218) );
  AOI22D1BWP30P140LVT U7732 ( .A1(i_data_bus[907]), .A2(n7527), .B1(
        i_data_bus[619]), .B2(n7529), .ZN(n7216) );
  AOI22D1BWP30P140LVT U7733 ( .A1(i_data_bus[523]), .A2(n7530), .B1(
        i_data_bus[555]), .B2(n7526), .ZN(n7215) );
  AOI22D1BWP30P140LVT U7734 ( .A1(i_data_bus[1003]), .A2(n7532), .B1(
        i_data_bus[587]), .B2(n7531), .ZN(n7214) );
  AOI22D1BWP30P140LVT U7735 ( .A1(i_data_bus[939]), .A2(n7528), .B1(
        i_data_bus[971]), .B2(n7525), .ZN(n7213) );
  ND4D1BWP30P140LVT U7736 ( .A1(n7216), .A2(n7215), .A3(n7214), .A4(n7213), 
        .ZN(n7217) );
  INR4D0BWP30P140LVT U7737 ( .A1(n7220), .B1(n7219), .B2(n7218), .B3(n7217), 
        .ZN(n7221) );
  ND4D4BWP30P140LVT U7738 ( .A1(n7224), .A2(n7223), .A3(n7222), .A4(n7221), 
        .ZN(o_data_bus[75]) );
  AOI22D1BWP30P140LVT U7739 ( .A1(i_data_bus[489]), .A2(n7459), .B1(
        i_data_bus[329]), .B2(n7493), .ZN(n7244) );
  AOI22D1BWP30P140LVT U7740 ( .A1(i_data_bus[265]), .A2(n7436), .B1(
        i_data_bus[457]), .B2(n7472), .ZN(n7243) );
  AOI22D1BWP30P140LVT U7741 ( .A1(i_data_bus[41]), .A2(n7514), .B1(
        i_data_bus[745]), .B2(n7504), .ZN(n7228) );
  AOI22D1BWP30P140LVT U7742 ( .A1(i_data_bus[73]), .A2(n7511), .B1(
        i_data_bus[841]), .B2(n7498), .ZN(n7227) );
  AOI22D1BWP30P140LVT U7743 ( .A1(i_data_bus[873]), .A2(n7497), .B1(
        i_data_bus[809]), .B2(n7513), .ZN(n7226) );
  AOI22D1BWP30P140LVT U7744 ( .A1(i_data_bus[681]), .A2(n7509), .B1(
        i_data_bus[777]), .B2(n7516), .ZN(n7225) );
  AN4D0BWP30P140LVT U7745 ( .A1(n7228), .A2(n7227), .A3(n7226), .A4(n7225), 
        .Z(n7242) );
  AOI22D1BWP30P140LVT U7746 ( .A1(i_data_bus[425]), .A2(n7523), .B1(
        i_data_bus[361]), .B2(n7495), .ZN(n7240) );
  AOI22D1BWP30P140LVT U7747 ( .A1(i_data_bus[201]), .A2(n7502), .B1(
        i_data_bus[233]), .B2(n7501), .ZN(n7232) );
  AOI22D1BWP30P140LVT U7748 ( .A1(i_data_bus[169]), .A2(n7515), .B1(
        i_data_bus[649]), .B2(n7499), .ZN(n7231) );
  AOI22D1BWP30P140LVT U7749 ( .A1(i_data_bus[9]), .A2(n7500), .B1(
        i_data_bus[137]), .B2(n7503), .ZN(n7230) );
  AOI22D1BWP30P140LVT U7750 ( .A1(i_data_bus[105]), .A2(n7512), .B1(
        i_data_bus[713]), .B2(n7510), .ZN(n7229) );
  ND4D1BWP30P140LVT U7751 ( .A1(n7232), .A2(n7231), .A3(n7230), .A4(n7229), 
        .ZN(n7239) );
  INVD1BWP30P140LVT U7752 ( .I(i_data_bus[297]), .ZN(n9688) );
  INVD1BWP30P140LVT U7753 ( .I(i_data_bus[393]), .ZN(n8313) );
  OAI22D1BWP30P140LVT U7754 ( .A1(n9688), .A2(n7394), .B1(n8313), .B2(n7411), 
        .ZN(n7238) );
  AOI22D1BWP30P140LVT U7755 ( .A1(i_data_bus[585]), .A2(n7531), .B1(
        i_data_bus[617]), .B2(n7529), .ZN(n7236) );
  AOI22D1BWP30P140LVT U7756 ( .A1(i_data_bus[521]), .A2(n7530), .B1(
        i_data_bus[969]), .B2(n7525), .ZN(n7235) );
  AOI22D1BWP30P140LVT U7757 ( .A1(i_data_bus[1001]), .A2(n7532), .B1(
        i_data_bus[937]), .B2(n7528), .ZN(n7234) );
  AOI22D1BWP30P140LVT U7758 ( .A1(i_data_bus[905]), .A2(n7527), .B1(
        i_data_bus[553]), .B2(n7526), .ZN(n7233) );
  ND4D1BWP30P140LVT U7759 ( .A1(n7236), .A2(n7235), .A3(n7234), .A4(n7233), 
        .ZN(n7237) );
  INR4D0BWP30P140LVT U7760 ( .A1(n7240), .B1(n7239), .B2(n7238), .B3(n7237), 
        .ZN(n7241) );
  ND4D4BWP30P140LVT U7761 ( .A1(n7244), .A2(n7243), .A3(n7242), .A4(n7241), 
        .ZN(o_data_bus[73]) );
  AOI22D1BWP30P140LVT U7762 ( .A1(i_data_bus[488]), .A2(n7459), .B1(
        i_data_bus[360]), .B2(n7495), .ZN(n7264) );
  AOI22D1BWP30P140LVT U7763 ( .A1(i_data_bus[264]), .A2(n7436), .B1(
        i_data_bus[424]), .B2(n7523), .ZN(n7263) );
  AOI22D1BWP30P140LVT U7764 ( .A1(i_data_bus[840]), .A2(n7498), .B1(
        i_data_bus[776]), .B2(n7516), .ZN(n7248) );
  AOI22D1BWP30P140LVT U7765 ( .A1(i_data_bus[72]), .A2(n7511), .B1(
        i_data_bus[744]), .B2(n7504), .ZN(n7247) );
  AOI22D1BWP30P140LVT U7766 ( .A1(i_data_bus[808]), .A2(n7513), .B1(
        i_data_bus[648]), .B2(n7499), .ZN(n7246) );
  AOI22D1BWP30P140LVT U7767 ( .A1(i_data_bus[680]), .A2(n7509), .B1(
        i_data_bus[136]), .B2(n7503), .ZN(n7245) );
  AN4D0BWP30P140LVT U7768 ( .A1(n7248), .A2(n7247), .A3(n7246), .A4(n7245), 
        .Z(n7262) );
  AOI22D1BWP30P140LVT U7769 ( .A1(i_data_bus[456]), .A2(n7472), .B1(
        i_data_bus[328]), .B2(n7493), .ZN(n7260) );
  AOI22D1BWP30P140LVT U7770 ( .A1(i_data_bus[872]), .A2(n7497), .B1(
        i_data_bus[232]), .B2(n7501), .ZN(n7252) );
  AOI22D1BWP30P140LVT U7771 ( .A1(i_data_bus[8]), .A2(n7500), .B1(
        i_data_bus[200]), .B2(n7502), .ZN(n7251) );
  AOI22D1BWP30P140LVT U7772 ( .A1(i_data_bus[40]), .A2(n7514), .B1(
        i_data_bus[712]), .B2(n7510), .ZN(n7250) );
  AOI22D1BWP30P140LVT U7773 ( .A1(i_data_bus[104]), .A2(n7512), .B1(
        i_data_bus[168]), .B2(n7515), .ZN(n7249) );
  ND4D1BWP30P140LVT U7774 ( .A1(n7252), .A2(n7251), .A3(n7250), .A4(n7249), 
        .ZN(n7259) );
  INVD1BWP30P140LVT U7775 ( .I(i_data_bus[296]), .ZN(n9462) );
  MOAI22D1BWP30P140LVT U7776 ( .A1(n9462), .A2(n7394), .B1(i_data_bus[392]), 
        .B2(n7496), .ZN(n7258) );
  AOI22D1BWP30P140LVT U7777 ( .A1(i_data_bus[1000]), .A2(n7532), .B1(
        i_data_bus[584]), .B2(n7531), .ZN(n7256) );
  AOI22D1BWP30P140LVT U7778 ( .A1(i_data_bus[616]), .A2(n7529), .B1(
        i_data_bus[520]), .B2(n7530), .ZN(n7255) );
  AOI22D1BWP30P140LVT U7779 ( .A1(i_data_bus[968]), .A2(n7525), .B1(
        i_data_bus[936]), .B2(n7528), .ZN(n7254) );
  AOI22D1BWP30P140LVT U7780 ( .A1(i_data_bus[552]), .A2(n7526), .B1(
        i_data_bus[904]), .B2(n7527), .ZN(n7253) );
  ND4D1BWP30P140LVT U7781 ( .A1(n7256), .A2(n7255), .A3(n7254), .A4(n7253), 
        .ZN(n7257) );
  INR4D0BWP30P140LVT U7782 ( .A1(n7260), .B1(n7259), .B2(n7258), .B3(n7257), 
        .ZN(n7261) );
  ND4D4BWP30P140LVT U7783 ( .A1(n7264), .A2(n7263), .A3(n7262), .A4(n7261), 
        .ZN(o_data_bus[72]) );
  AOI22D1BWP30P140LVT U7784 ( .A1(i_data_bus[404]), .A2(n7496), .B1(
        i_data_bus[500]), .B2(n7459), .ZN(n7284) );
  AOI22D1BWP30P140LVT U7785 ( .A1(i_data_bus[340]), .A2(n7493), .B1(
        i_data_bus[276]), .B2(n7436), .ZN(n7283) );
  AOI22D1BWP30P140LVT U7786 ( .A1(i_data_bus[948]), .A2(n7528), .B1(
        i_data_bus[916]), .B2(n7527), .ZN(n7268) );
  AOI22D1BWP30P140LVT U7787 ( .A1(i_data_bus[1012]), .A2(n7532), .B1(
        i_data_bus[564]), .B2(n7526), .ZN(n7267) );
  AOI22D1BWP30P140LVT U7788 ( .A1(i_data_bus[596]), .A2(n7531), .B1(
        i_data_bus[532]), .B2(n7530), .ZN(n7266) );
  AOI22D1BWP30P140LVT U7789 ( .A1(i_data_bus[980]), .A2(n7525), .B1(
        i_data_bus[628]), .B2(n7529), .ZN(n7265) );
  AN4D0BWP30P140LVT U7790 ( .A1(n7268), .A2(n7267), .A3(n7266), .A4(n7265), 
        .Z(n7282) );
  INVD1BWP30P140LVT U7791 ( .I(i_data_bus[468]), .ZN(n8128) );
  MOAI22D1BWP30P140LVT U7792 ( .A1(n8128), .A2(n7522), .B1(i_data_bus[372]), 
        .B2(n7495), .ZN(n7280) );
  INVD1BWP30P140LVT U7793 ( .I(i_data_bus[308]), .ZN(n9354) );
  MOAI22D1BWP30P140LVT U7794 ( .A1(n9354), .A2(n7394), .B1(i_data_bus[436]), 
        .B2(n7523), .ZN(n7279) );
  AOI22D1BWP30P140LVT U7795 ( .A1(i_data_bus[212]), .A2(n7502), .B1(
        i_data_bus[180]), .B2(n7515), .ZN(n7272) );
  AOI22D1BWP30P140LVT U7796 ( .A1(i_data_bus[52]), .A2(n7514), .B1(
        i_data_bus[788]), .B2(n7516), .ZN(n7271) );
  AOI22D1BWP30P140LVT U7797 ( .A1(i_data_bus[852]), .A2(n7498), .B1(
        i_data_bus[148]), .B2(n7503), .ZN(n7270) );
  AOI22D1BWP30P140LVT U7798 ( .A1(i_data_bus[884]), .A2(n7497), .B1(
        i_data_bus[660]), .B2(n7499), .ZN(n7269) );
  ND4D1BWP30P140LVT U7799 ( .A1(n7272), .A2(n7271), .A3(n7270), .A4(n7269), 
        .ZN(n7278) );
  AOI22D1BWP30P140LVT U7800 ( .A1(i_data_bus[20]), .A2(n7500), .B1(
        i_data_bus[724]), .B2(n7510), .ZN(n7276) );
  AOI22D1BWP30P140LVT U7801 ( .A1(i_data_bus[244]), .A2(n7501), .B1(
        i_data_bus[756]), .B2(n7504), .ZN(n7275) );
  AOI22D1BWP30P140LVT U7802 ( .A1(i_data_bus[116]), .A2(n7512), .B1(
        i_data_bus[820]), .B2(n7513), .ZN(n7274) );
  AOI22D1BWP30P140LVT U7803 ( .A1(i_data_bus[84]), .A2(n7511), .B1(
        i_data_bus[692]), .B2(n7509), .ZN(n7273) );
  ND4D1BWP30P140LVT U7804 ( .A1(n7276), .A2(n7275), .A3(n7274), .A4(n7273), 
        .ZN(n7277) );
  NR4D0BWP30P140LVT U7805 ( .A1(n7280), .A2(n7279), .A3(n7278), .A4(n7277), 
        .ZN(n7281) );
  ND4D4BWP30P140LVT U7806 ( .A1(n7284), .A2(n7283), .A3(n7282), .A4(n7281), 
        .ZN(o_data_bus[84]) );
  AOI22D1BWP30P140LVT U7807 ( .A1(i_data_bus[433]), .A2(n7523), .B1(
        i_data_bus[401]), .B2(n7496), .ZN(n7304) );
  AOI22D1BWP30P140LVT U7808 ( .A1(i_data_bus[465]), .A2(n7472), .B1(
        i_data_bus[497]), .B2(n7459), .ZN(n7303) );
  AOI22D1BWP30P140LVT U7809 ( .A1(i_data_bus[881]), .A2(n7497), .B1(
        i_data_bus[145]), .B2(n7503), .ZN(n7288) );
  AOI22D1BWP30P140LVT U7810 ( .A1(i_data_bus[657]), .A2(n7499), .B1(
        i_data_bus[753]), .B2(n7504), .ZN(n7287) );
  AOI22D1BWP30P140LVT U7811 ( .A1(i_data_bus[849]), .A2(n7498), .B1(
        i_data_bus[817]), .B2(n7513), .ZN(n7286) );
  AOI22D1BWP30P140LVT U7812 ( .A1(i_data_bus[785]), .A2(n7516), .B1(
        i_data_bus[721]), .B2(n7510), .ZN(n7285) );
  AN4D0BWP30P140LVT U7813 ( .A1(n7288), .A2(n7287), .A3(n7286), .A4(n7285), 
        .Z(n7302) );
  AOI22D1BWP30P140LVT U7814 ( .A1(i_data_bus[337]), .A2(n7493), .B1(
        i_data_bus[273]), .B2(n7436), .ZN(n7300) );
  AOI22D1BWP30P140LVT U7815 ( .A1(i_data_bus[17]), .A2(n7500), .B1(
        i_data_bus[49]), .B2(n7514), .ZN(n7292) );
  AOI22D1BWP30P140LVT U7816 ( .A1(i_data_bus[241]), .A2(n7501), .B1(
        i_data_bus[209]), .B2(n7502), .ZN(n7291) );
  AOI22D1BWP30P140LVT U7817 ( .A1(i_data_bus[81]), .A2(n7511), .B1(
        i_data_bus[689]), .B2(n7509), .ZN(n7290) );
  AOI22D1BWP30P140LVT U7818 ( .A1(i_data_bus[113]), .A2(n7512), .B1(
        i_data_bus[177]), .B2(n7515), .ZN(n7289) );
  ND4D1BWP30P140LVT U7819 ( .A1(n7292), .A2(n7291), .A3(n7290), .A4(n7289), 
        .ZN(n7299) );
  INVD1BWP30P140LVT U7820 ( .I(i_data_bus[369]), .ZN(n9376) );
  MOAI22D1BWP30P140LVT U7821 ( .A1(n9376), .A2(n7369), .B1(i_data_bus[305]), 
        .B2(n7494), .ZN(n7298) );
  AOI22D1BWP30P140LVT U7822 ( .A1(i_data_bus[625]), .A2(n7529), .B1(
        i_data_bus[1009]), .B2(n7532), .ZN(n7296) );
  AOI22D1BWP30P140LVT U7823 ( .A1(i_data_bus[593]), .A2(n7531), .B1(
        i_data_bus[529]), .B2(n7530), .ZN(n7295) );
  AOI22D1BWP30P140LVT U7824 ( .A1(i_data_bus[945]), .A2(n7528), .B1(
        i_data_bus[977]), .B2(n7525), .ZN(n7294) );
  AOI22D1BWP30P140LVT U7825 ( .A1(i_data_bus[913]), .A2(n7527), .B1(
        i_data_bus[561]), .B2(n7526), .ZN(n7293) );
  ND4D1BWP30P140LVT U7826 ( .A1(n7296), .A2(n7295), .A3(n7294), .A4(n7293), 
        .ZN(n7297) );
  INR4D0BWP30P140LVT U7827 ( .A1(n7300), .B1(n7299), .B2(n7298), .B3(n7297), 
        .ZN(n7301) );
  ND4D4BWP30P140LVT U7828 ( .A1(n7304), .A2(n7303), .A3(n7302), .A4(n7301), 
        .ZN(o_data_bus[81]) );
  AOI22D1BWP30P140LVT U7829 ( .A1(i_data_bus[271]), .A2(n7436), .B1(
        i_data_bus[303]), .B2(n7494), .ZN(n7324) );
  AOI22D1BWP30P140LVT U7830 ( .A1(i_data_bus[431]), .A2(n7523), .B1(
        i_data_bus[335]), .B2(n7493), .ZN(n7323) );
  AOI22D1BWP30P140LVT U7831 ( .A1(i_data_bus[911]), .A2(n7527), .B1(
        i_data_bus[623]), .B2(n7529), .ZN(n7308) );
  AOI22D1BWP30P140LVT U7832 ( .A1(i_data_bus[975]), .A2(n7525), .B1(
        i_data_bus[527]), .B2(n7530), .ZN(n7307) );
  AOI22D1BWP30P140LVT U7833 ( .A1(i_data_bus[1007]), .A2(n7532), .B1(
        i_data_bus[943]), .B2(n7528), .ZN(n7306) );
  AOI22D1BWP30P140LVT U7834 ( .A1(i_data_bus[591]), .A2(n7531), .B1(
        i_data_bus[559]), .B2(n7526), .ZN(n7305) );
  AN4D0BWP30P140LVT U7835 ( .A1(n7308), .A2(n7307), .A3(n7306), .A4(n7305), 
        .Z(n7322) );
  INVD1BWP30P140LVT U7836 ( .I(i_data_bus[463]), .ZN(n8230) );
  MOAI22D1BWP30P140LVT U7837 ( .A1(n8230), .A2(n7522), .B1(i_data_bus[495]), 
        .B2(n7459), .ZN(n7320) );
  INVD1BWP30P140LVT U7838 ( .I(i_data_bus[399]), .ZN(n8845) );
  INVD1BWP30P140LVT U7839 ( .I(i_data_bus[367]), .ZN(n7920) );
  OAI22D1BWP30P140LVT U7840 ( .A1(n8845), .A2(n7411), .B1(n7920), .B2(n7369), 
        .ZN(n7319) );
  AOI22D1BWP30P140LVT U7841 ( .A1(i_data_bus[143]), .A2(n7503), .B1(
        i_data_bus[655]), .B2(n7499), .ZN(n7312) );
  AOI22D1BWP30P140LVT U7842 ( .A1(i_data_bus[47]), .A2(n7514), .B1(
        i_data_bus[687]), .B2(n7509), .ZN(n7311) );
  AOI22D1BWP30P140LVT U7843 ( .A1(i_data_bus[15]), .A2(n7500), .B1(
        i_data_bus[239]), .B2(n7501), .ZN(n7310) );
  AOI22D1BWP30P140LVT U7844 ( .A1(i_data_bus[207]), .A2(n7502), .B1(
        i_data_bus[879]), .B2(n7497), .ZN(n7309) );
  ND4D1BWP30P140LVT U7845 ( .A1(n7312), .A2(n7311), .A3(n7310), .A4(n7309), 
        .ZN(n7318) );
  AOI22D1BWP30P140LVT U7846 ( .A1(i_data_bus[79]), .A2(n7511), .B1(
        i_data_bus[175]), .B2(n7515), .ZN(n7316) );
  AOI22D1BWP30P140LVT U7847 ( .A1(i_data_bus[719]), .A2(n7510), .B1(
        i_data_bus[783]), .B2(n7516), .ZN(n7315) );
  AOI22D1BWP30P140LVT U7848 ( .A1(i_data_bus[111]), .A2(n7512), .B1(
        i_data_bus[751]), .B2(n7504), .ZN(n7314) );
  AOI22D1BWP30P140LVT U7849 ( .A1(i_data_bus[847]), .A2(n7498), .B1(
        i_data_bus[815]), .B2(n7513), .ZN(n7313) );
  ND4D1BWP30P140LVT U7850 ( .A1(n7316), .A2(n7315), .A3(n7314), .A4(n7313), 
        .ZN(n7317) );
  NR4D0BWP30P140LVT U7851 ( .A1(n7320), .A2(n7319), .A3(n7318), .A4(n7317), 
        .ZN(n7321) );
  ND4D4BWP30P140LVT U7852 ( .A1(n7324), .A2(n7323), .A3(n7322), .A4(n7321), 
        .ZN(o_data_bus[79]) );
  AOI22D1BWP30P140LVT U7853 ( .A1(i_data_bus[298]), .A2(n7494), .B1(
        i_data_bus[426]), .B2(n7523), .ZN(n7344) );
  AOI22D1BWP30P140LVT U7854 ( .A1(i_data_bus[458]), .A2(n7472), .B1(
        i_data_bus[266]), .B2(n7436), .ZN(n7343) );
  AOI22D1BWP30P140LVT U7855 ( .A1(i_data_bus[234]), .A2(n7501), .B1(
        i_data_bus[874]), .B2(n7497), .ZN(n7328) );
  AOI22D1BWP30P140LVT U7856 ( .A1(i_data_bus[106]), .A2(n7512), .B1(
        i_data_bus[170]), .B2(n7515), .ZN(n7327) );
  AOI22D1BWP30P140LVT U7857 ( .A1(i_data_bus[42]), .A2(n7514), .B1(
        i_data_bus[74]), .B2(n7511), .ZN(n7326) );
  AOI22D1BWP30P140LVT U7858 ( .A1(i_data_bus[714]), .A2(n7510), .B1(
        i_data_bus[682]), .B2(n7509), .ZN(n7325) );
  AN4D0BWP30P140LVT U7859 ( .A1(n7328), .A2(n7327), .A3(n7326), .A4(n7325), 
        .Z(n7342) );
  AOI22D1BWP30P140LVT U7860 ( .A1(i_data_bus[650]), .A2(n7499), .B1(
        i_data_bus[746]), .B2(n7504), .ZN(n7332) );
  AOI22D1BWP30P140LVT U7861 ( .A1(i_data_bus[10]), .A2(n7500), .B1(
        i_data_bus[778]), .B2(n7516), .ZN(n7331) );
  AOI22D1BWP30P140LVT U7862 ( .A1(i_data_bus[202]), .A2(n7502), .B1(
        i_data_bus[810]), .B2(n7513), .ZN(n7330) );
  AOI22D1BWP30P140LVT U7863 ( .A1(i_data_bus[842]), .A2(n7498), .B1(
        i_data_bus[138]), .B2(n7503), .ZN(n7329) );
  ND4D1BWP30P140LVT U7864 ( .A1(n7332), .A2(n7331), .A3(n7330), .A4(n7329), 
        .ZN(n7340) );
  INVD1BWP30P140LVT U7865 ( .I(i_data_bus[490]), .ZN(n8887) );
  MOAI22D1BWP30P140LVT U7866 ( .A1(n8887), .A2(n7524), .B1(i_data_bus[362]), 
        .B2(n7495), .ZN(n7339) );
  INVD1BWP30P140LVT U7867 ( .I(i_data_bus[394]), .ZN(n8535) );
  MOAI22D1BWP30P140LVT U7868 ( .A1(n8535), .A2(n7411), .B1(i_data_bus[330]), 
        .B2(n7493), .ZN(n7338) );
  AOI22D1BWP30P140LVT U7869 ( .A1(i_data_bus[970]), .A2(n7525), .B1(
        i_data_bus[522]), .B2(n7530), .ZN(n7336) );
  AOI22D1BWP30P140LVT U7870 ( .A1(i_data_bus[618]), .A2(n7529), .B1(
        i_data_bus[938]), .B2(n7528), .ZN(n7335) );
  AOI22D1BWP30P140LVT U7871 ( .A1(i_data_bus[554]), .A2(n7526), .B1(
        i_data_bus[586]), .B2(n7531), .ZN(n7334) );
  AOI22D1BWP30P140LVT U7872 ( .A1(i_data_bus[1002]), .A2(n7532), .B1(
        i_data_bus[906]), .B2(n7527), .ZN(n7333) );
  ND4D1BWP30P140LVT U7873 ( .A1(n7336), .A2(n7335), .A3(n7334), .A4(n7333), 
        .ZN(n7337) );
  NR4D0BWP30P140LVT U7874 ( .A1(n7340), .A2(n7339), .A3(n7338), .A4(n7337), 
        .ZN(n7341) );
  ND4D4BWP30P140LVT U7875 ( .A1(n7344), .A2(n7343), .A3(n7342), .A4(n7341), 
        .ZN(o_data_bus[74]) );
  AOI22D1BWP30P140LVT U7876 ( .A1(i_data_bus[358]), .A2(n7495), .B1(
        i_data_bus[262]), .B2(n7436), .ZN(n7364) );
  AOI22D1BWP30P140LVT U7877 ( .A1(i_data_bus[294]), .A2(n7494), .B1(
        i_data_bus[326]), .B2(n7493), .ZN(n7363) );
  AOI22D1BWP30P140LVT U7878 ( .A1(i_data_bus[582]), .A2(n7531), .B1(
        i_data_bus[998]), .B2(n7532), .ZN(n7348) );
  AOI22D1BWP30P140LVT U7879 ( .A1(i_data_bus[614]), .A2(n7529), .B1(
        i_data_bus[934]), .B2(n7528), .ZN(n7347) );
  AOI22D1BWP30P140LVT U7880 ( .A1(i_data_bus[966]), .A2(n7525), .B1(
        i_data_bus[518]), .B2(n7530), .ZN(n7346) );
  AOI22D1BWP30P140LVT U7881 ( .A1(i_data_bus[550]), .A2(n7526), .B1(
        i_data_bus[902]), .B2(n7527), .ZN(n7345) );
  AN4D0BWP30P140LVT U7882 ( .A1(n7348), .A2(n7347), .A3(n7346), .A4(n7345), 
        .Z(n7362) );
  AOI22D1BWP30P140LVT U7883 ( .A1(i_data_bus[486]), .A2(n7459), .B1(
        i_data_bus[422]), .B2(n7523), .ZN(n7360) );
  INVD1BWP30P140LVT U7884 ( .I(i_data_bus[390]), .ZN(n8993) );
  INVD1BWP30P140LVT U7885 ( .I(i_data_bus[454]), .ZN(n9505) );
  OAI22D1BWP30P140LVT U7886 ( .A1(n8993), .A2(n7411), .B1(n9505), .B2(n7522), 
        .ZN(n7359) );
  AOI22D1BWP30P140LVT U7887 ( .A1(i_data_bus[38]), .A2(n7514), .B1(
        i_data_bus[806]), .B2(n7513), .ZN(n7352) );
  AOI22D1BWP30P140LVT U7888 ( .A1(i_data_bus[198]), .A2(n7502), .B1(
        i_data_bus[678]), .B2(n7509), .ZN(n7351) );
  AOI22D1BWP30P140LVT U7889 ( .A1(i_data_bus[646]), .A2(n7499), .B1(
        i_data_bus[774]), .B2(n7516), .ZN(n7350) );
  AOI22D1BWP30P140LVT U7890 ( .A1(i_data_bus[6]), .A2(n7500), .B1(
        i_data_bus[230]), .B2(n7501), .ZN(n7349) );
  ND4D1BWP30P140LVT U7891 ( .A1(n7352), .A2(n7351), .A3(n7350), .A4(n7349), 
        .ZN(n7358) );
  AOI22D1BWP30P140LVT U7892 ( .A1(i_data_bus[742]), .A2(n7504), .B1(
        i_data_bus[710]), .B2(n7510), .ZN(n7356) );
  AOI22D1BWP30P140LVT U7893 ( .A1(i_data_bus[70]), .A2(n7511), .B1(
        i_data_bus[870]), .B2(n7497), .ZN(n7355) );
  AOI22D1BWP30P140LVT U7894 ( .A1(i_data_bus[102]), .A2(n7512), .B1(
        i_data_bus[134]), .B2(n7503), .ZN(n7354) );
  AOI22D1BWP30P140LVT U7895 ( .A1(i_data_bus[838]), .A2(n7498), .B1(
        i_data_bus[166]), .B2(n7515), .ZN(n7353) );
  ND4D1BWP30P140LVT U7896 ( .A1(n7356), .A2(n7355), .A3(n7354), .A4(n7353), 
        .ZN(n7357) );
  INR4D0BWP30P140LVT U7897 ( .A1(n7360), .B1(n7359), .B2(n7358), .B3(n7357), 
        .ZN(n7361) );
  ND4D4BWP30P140LVT U7898 ( .A1(n7364), .A2(n7363), .A3(n7362), .A4(n7361), 
        .ZN(o_data_bus[70]) );
  AOI22D1BWP30P140LVT U7899 ( .A1(i_data_bus[455]), .A2(n7472), .B1(
        i_data_bus[423]), .B2(n7523), .ZN(n7385) );
  AOI22D1BWP30P140LVT U7900 ( .A1(i_data_bus[263]), .A2(n7436), .B1(
        i_data_bus[391]), .B2(n7496), .ZN(n7384) );
  AOI22D1BWP30P140LVT U7901 ( .A1(i_data_bus[903]), .A2(n7527), .B1(
        i_data_bus[967]), .B2(n7525), .ZN(n7368) );
  AOI22D1BWP30P140LVT U7902 ( .A1(i_data_bus[519]), .A2(n7530), .B1(
        i_data_bus[551]), .B2(n7526), .ZN(n7367) );
  AOI22D1BWP30P140LVT U7903 ( .A1(i_data_bus[615]), .A2(n7529), .B1(
        i_data_bus[583]), .B2(n7531), .ZN(n7366) );
  AOI22D1BWP30P140LVT U7904 ( .A1(i_data_bus[999]), .A2(n7532), .B1(
        i_data_bus[935]), .B2(n7528), .ZN(n7365) );
  AN4D0BWP30P140LVT U7905 ( .A1(n7368), .A2(n7367), .A3(n7366), .A4(n7365), 
        .Z(n7383) );
  INVD1BWP30P140LVT U7906 ( .I(i_data_bus[359]), .ZN(n8908) );
  MOAI22D1BWP30P140LVT U7907 ( .A1(n8908), .A2(n7369), .B1(i_data_bus[295]), 
        .B2(n7494), .ZN(n7381) );
  INVD1BWP30P140LVT U7908 ( .I(i_data_bus[487]), .ZN(n8625) );
  MOAI22D1BWP30P140LVT U7909 ( .A1(n8625), .A2(n7524), .B1(i_data_bus[327]), 
        .B2(n7493), .ZN(n7380) );
  AOI22D1BWP30P140LVT U7910 ( .A1(i_data_bus[743]), .A2(n7504), .B1(
        i_data_bus[167]), .B2(n7515), .ZN(n7373) );
  AOI22D1BWP30P140LVT U7911 ( .A1(i_data_bus[679]), .A2(n7509), .B1(
        i_data_bus[647]), .B2(n7499), .ZN(n7372) );
  AOI22D1BWP30P140LVT U7912 ( .A1(i_data_bus[71]), .A2(n7511), .B1(
        i_data_bus[231]), .B2(n7501), .ZN(n7371) );
  AOI22D1BWP30P140LVT U7913 ( .A1(i_data_bus[39]), .A2(n7514), .B1(
        i_data_bus[7]), .B2(n7500), .ZN(n7370) );
  ND4D1BWP30P140LVT U7914 ( .A1(n7373), .A2(n7372), .A3(n7371), .A4(n7370), 
        .ZN(n7379) );
  AOI22D1BWP30P140LVT U7915 ( .A1(i_data_bus[839]), .A2(n7498), .B1(
        i_data_bus[775]), .B2(n7516), .ZN(n7377) );
  AOI22D1BWP30P140LVT U7916 ( .A1(i_data_bus[135]), .A2(n7503), .B1(
        i_data_bus[199]), .B2(n7502), .ZN(n7376) );
  AOI22D1BWP30P140LVT U7917 ( .A1(i_data_bus[871]), .A2(n7497), .B1(
        i_data_bus[711]), .B2(n7510), .ZN(n7375) );
  AOI22D1BWP30P140LVT U7918 ( .A1(i_data_bus[103]), .A2(n7512), .B1(
        i_data_bus[807]), .B2(n7513), .ZN(n7374) );
  ND4D1BWP30P140LVT U7919 ( .A1(n7377), .A2(n7376), .A3(n7375), .A4(n7374), 
        .ZN(n7378) );
  NR4D0BWP30P140LVT U7920 ( .A1(n7381), .A2(n7380), .A3(n7379), .A4(n7378), 
        .ZN(n7382) );
  ND4D4BWP30P140LVT U7921 ( .A1(n7385), .A2(n7384), .A3(n7383), .A4(n7382), 
        .ZN(o_data_bus[71]) );
  AOI22D1BWP30P140LVT U7922 ( .A1(i_data_bus[421]), .A2(n7523), .B1(
        i_data_bus[261]), .B2(n7436), .ZN(n7406) );
  AOI22D1BWP30P140LVT U7923 ( .A1(i_data_bus[453]), .A2(n7472), .B1(
        i_data_bus[325]), .B2(n7493), .ZN(n7405) );
  AOI22D1BWP30P140LVT U7924 ( .A1(i_data_bus[677]), .A2(n7509), .B1(
        i_data_bus[741]), .B2(n7504), .ZN(n7389) );
  AOI22D1BWP30P140LVT U7925 ( .A1(i_data_bus[37]), .A2(n7514), .B1(
        i_data_bus[709]), .B2(n7510), .ZN(n7388) );
  AOI22D1BWP30P140LVT U7926 ( .A1(i_data_bus[645]), .A2(n7499), .B1(
        i_data_bus[805]), .B2(n7513), .ZN(n7387) );
  AOI22D1BWP30P140LVT U7927 ( .A1(i_data_bus[101]), .A2(n7512), .B1(
        i_data_bus[69]), .B2(n7511), .ZN(n7386) );
  AN4D0BWP30P140LVT U7928 ( .A1(n7389), .A2(n7388), .A3(n7387), .A4(n7386), 
        .Z(n7404) );
  AOI22D1BWP30P140LVT U7929 ( .A1(i_data_bus[357]), .A2(n7495), .B1(
        i_data_bus[389]), .B2(n7496), .ZN(n7402) );
  AOI22D1BWP30P140LVT U7930 ( .A1(i_data_bus[773]), .A2(n7516), .B1(
        i_data_bus[837]), .B2(n7498), .ZN(n7393) );
  AOI22D1BWP30P140LVT U7931 ( .A1(i_data_bus[197]), .A2(n7502), .B1(
        i_data_bus[869]), .B2(n7497), .ZN(n7392) );
  AOI22D1BWP30P140LVT U7932 ( .A1(i_data_bus[165]), .A2(n7515), .B1(
        i_data_bus[229]), .B2(n7501), .ZN(n7391) );
  AOI22D1BWP30P140LVT U7933 ( .A1(i_data_bus[5]), .A2(n7500), .B1(
        i_data_bus[133]), .B2(n7503), .ZN(n7390) );
  ND4D1BWP30P140LVT U7934 ( .A1(n7393), .A2(n7392), .A3(n7391), .A4(n7390), 
        .ZN(n7401) );
  INVD1BWP30P140LVT U7935 ( .I(i_data_bus[293]), .ZN(n9333) );
  MOAI22D1BWP30P140LVT U7936 ( .A1(n9333), .A2(n7394), .B1(i_data_bus[485]), 
        .B2(n7459), .ZN(n7400) );
  AOI22D1BWP30P140LVT U7937 ( .A1(i_data_bus[581]), .A2(n7531), .B1(
        i_data_bus[933]), .B2(n7528), .ZN(n7398) );
  AOI22D1BWP30P140LVT U7938 ( .A1(i_data_bus[901]), .A2(n7527), .B1(
        i_data_bus[549]), .B2(n7526), .ZN(n7397) );
  AOI22D1BWP30P140LVT U7939 ( .A1(i_data_bus[517]), .A2(n7530), .B1(
        i_data_bus[965]), .B2(n7525), .ZN(n7396) );
  AOI22D1BWP30P140LVT U7940 ( .A1(i_data_bus[613]), .A2(n7529), .B1(
        i_data_bus[997]), .B2(n7532), .ZN(n7395) );
  ND4D1BWP30P140LVT U7941 ( .A1(n7398), .A2(n7397), .A3(n7396), .A4(n7395), 
        .ZN(n7399) );
  INR4D0BWP30P140LVT U7942 ( .A1(n7402), .B1(n7401), .B2(n7400), .B3(n7399), 
        .ZN(n7403) );
  ND4D4BWP30P140LVT U7943 ( .A1(n7406), .A2(n7405), .A3(n7404), .A4(n7403), 
        .ZN(o_data_bus[69]) );
  AOI22D1BWP30P140LVT U7944 ( .A1(i_data_bus[420]), .A2(n7523), .B1(
        i_data_bus[292]), .B2(n7494), .ZN(n7427) );
  AOI22D1BWP30P140LVT U7945 ( .A1(i_data_bus[356]), .A2(n7495), .B1(
        i_data_bus[260]), .B2(n7436), .ZN(n7426) );
  AOI22D1BWP30P140LVT U7946 ( .A1(i_data_bus[612]), .A2(n7529), .B1(
        i_data_bus[900]), .B2(n7527), .ZN(n7410) );
  AOI22D1BWP30P140LVT U7947 ( .A1(i_data_bus[548]), .A2(n7526), .B1(
        i_data_bus[932]), .B2(n7528), .ZN(n7409) );
  AOI22D1BWP30P140LVT U7948 ( .A1(i_data_bus[964]), .A2(n7525), .B1(
        i_data_bus[580]), .B2(n7531), .ZN(n7408) );
  AOI22D1BWP30P140LVT U7949 ( .A1(i_data_bus[516]), .A2(n7530), .B1(
        i_data_bus[996]), .B2(n7532), .ZN(n7407) );
  AN4D0BWP30P140LVT U7950 ( .A1(n7410), .A2(n7409), .A3(n7408), .A4(n7407), 
        .Z(n7425) );
  INVD1BWP30P140LVT U7951 ( .I(i_data_bus[388]), .ZN(n8648) );
  MOAI22D1BWP30P140LVT U7952 ( .A1(n8648), .A2(n7411), .B1(i_data_bus[484]), 
        .B2(n7459), .ZN(n7423) );
  INVD1BWP30P140LVT U7953 ( .I(i_data_bus[452]), .ZN(n9527) );
  INVD1BWP30P140LVT U7954 ( .I(i_data_bus[324]), .ZN(n9116) );
  OAI22D1BWP30P140LVT U7955 ( .A1(n9527), .A2(n7522), .B1(n9116), .B2(n7458), 
        .ZN(n7422) );
  AOI22D1BWP30P140LVT U7956 ( .A1(i_data_bus[228]), .A2(n7501), .B1(
        i_data_bus[868]), .B2(n7497), .ZN(n7415) );
  AOI22D1BWP30P140LVT U7957 ( .A1(i_data_bus[708]), .A2(n7510), .B1(
        i_data_bus[644]), .B2(n7499), .ZN(n7414) );
  AOI22D1BWP30P140LVT U7958 ( .A1(i_data_bus[4]), .A2(n7500), .B1(
        i_data_bus[740]), .B2(n7504), .ZN(n7413) );
  AOI22D1BWP30P140LVT U7959 ( .A1(i_data_bus[132]), .A2(n7503), .B1(
        i_data_bus[804]), .B2(n7513), .ZN(n7412) );
  ND4D1BWP30P140LVT U7960 ( .A1(n7415), .A2(n7414), .A3(n7413), .A4(n7412), 
        .ZN(n7421) );
  AOI22D1BWP30P140LVT U7961 ( .A1(i_data_bus[100]), .A2(n7512), .B1(
        i_data_bus[68]), .B2(n7511), .ZN(n7419) );
  AOI22D1BWP30P140LVT U7962 ( .A1(i_data_bus[196]), .A2(n7502), .B1(
        i_data_bus[772]), .B2(n7516), .ZN(n7418) );
  AOI22D1BWP30P140LVT U7963 ( .A1(i_data_bus[36]), .A2(n7514), .B1(
        i_data_bus[836]), .B2(n7498), .ZN(n7417) );
  AOI22D1BWP30P140LVT U7964 ( .A1(i_data_bus[676]), .A2(n7509), .B1(
        i_data_bus[164]), .B2(n7515), .ZN(n7416) );
  ND4D1BWP30P140LVT U7965 ( .A1(n7419), .A2(n7418), .A3(n7417), .A4(n7416), 
        .ZN(n7420) );
  NR4D0BWP30P140LVT U7966 ( .A1(n7423), .A2(n7422), .A3(n7421), .A4(n7420), 
        .ZN(n7424) );
  ND4D4BWP30P140LVT U7967 ( .A1(n7427), .A2(n7426), .A3(n7425), .A4(n7424), 
        .ZN(o_data_bus[68]) );
  AOI22D1BWP30P140LVT U7968 ( .A1(i_data_bus[323]), .A2(n7493), .B1(
        i_data_bus[291]), .B2(n7494), .ZN(n7449) );
  AOI22D1BWP30P140LVT U7969 ( .A1(i_data_bus[387]), .A2(n7496), .B1(
        i_data_bus[483]), .B2(n7459), .ZN(n7448) );
  AOI22D1BWP30P140LVT U7970 ( .A1(i_data_bus[227]), .A2(n7501), .B1(
        i_data_bus[195]), .B2(n7502), .ZN(n7431) );
  AOI22D1BWP30P140LVT U7971 ( .A1(i_data_bus[643]), .A2(n7499), .B1(
        i_data_bus[867]), .B2(n7497), .ZN(n7430) );
  AOI22D1BWP30P140LVT U7972 ( .A1(i_data_bus[35]), .A2(n7514), .B1(
        i_data_bus[835]), .B2(n7498), .ZN(n7429) );
  AOI22D1BWP30P140LVT U7973 ( .A1(i_data_bus[3]), .A2(n7500), .B1(
        i_data_bus[99]), .B2(n7512), .ZN(n7428) );
  AN4D0BWP30P140LVT U7974 ( .A1(n7431), .A2(n7430), .A3(n7429), .A4(n7428), 
        .Z(n7447) );
  AOI22D1BWP30P140LVT U7975 ( .A1(i_data_bus[163]), .A2(n7515), .B1(
        i_data_bus[803]), .B2(n7513), .ZN(n7435) );
  AOI22D1BWP30P140LVT U7976 ( .A1(i_data_bus[131]), .A2(n7503), .B1(
        i_data_bus[675]), .B2(n7509), .ZN(n7434) );
  AOI22D1BWP30P140LVT U7977 ( .A1(i_data_bus[771]), .A2(n7516), .B1(
        i_data_bus[739]), .B2(n7504), .ZN(n7433) );
  AOI22D1BWP30P140LVT U7978 ( .A1(i_data_bus[67]), .A2(n7511), .B1(
        i_data_bus[707]), .B2(n7510), .ZN(n7432) );
  ND4D1BWP30P140LVT U7979 ( .A1(n7435), .A2(n7434), .A3(n7433), .A4(n7432), 
        .ZN(n7445) );
  INVD1BWP30P140LVT U7980 ( .I(i_data_bus[451]), .ZN(n8669) );
  MOAI22D1BWP30P140LVT U7981 ( .A1(n8669), .A2(n7522), .B1(i_data_bus[355]), 
        .B2(n7495), .ZN(n7444) );
  INVD1BWP30P140LVT U7982 ( .I(i_data_bus[419]), .ZN(n9567) );
  MOAI22D1BWP30P140LVT U7983 ( .A1(n9567), .A2(n7437), .B1(i_data_bus[259]), 
        .B2(n7436), .ZN(n7443) );
  AOI22D1BWP30P140LVT U7984 ( .A1(i_data_bus[515]), .A2(n7530), .B1(
        i_data_bus[995]), .B2(n7532), .ZN(n7441) );
  AOI22D1BWP30P140LVT U7985 ( .A1(i_data_bus[899]), .A2(n7527), .B1(
        i_data_bus[611]), .B2(n7529), .ZN(n7440) );
  AOI22D1BWP30P140LVT U7986 ( .A1(i_data_bus[963]), .A2(n7525), .B1(
        i_data_bus[931]), .B2(n7528), .ZN(n7439) );
  AOI22D1BWP30P140LVT U7987 ( .A1(i_data_bus[579]), .A2(n7531), .B1(
        i_data_bus[547]), .B2(n7526), .ZN(n7438) );
  ND4D1BWP30P140LVT U7988 ( .A1(n7441), .A2(n7440), .A3(n7439), .A4(n7438), 
        .ZN(n7442) );
  NR4D0BWP30P140LVT U7989 ( .A1(n7445), .A2(n7444), .A3(n7443), .A4(n7442), 
        .ZN(n7446) );
  ND4D4BWP30P140LVT U7990 ( .A1(n7449), .A2(n7448), .A3(n7447), .A4(n7446), 
        .ZN(o_data_bus[67]) );
  AOI22D1BWP30P140LVT U7991 ( .A1(i_data_bus[386]), .A2(n7496), .B1(
        i_data_bus[354]), .B2(n7495), .ZN(n7471) );
  AOI22D1BWP30P140LVT U7992 ( .A1(i_data_bus[290]), .A2(n7494), .B1(
        i_data_bus[418]), .B2(n7523), .ZN(n7470) );
  AOI22D1BWP30P140LVT U7993 ( .A1(i_data_bus[162]), .A2(n7515), .B1(
        i_data_bus[130]), .B2(n7503), .ZN(n7453) );
  AOI22D1BWP30P140LVT U7994 ( .A1(i_data_bus[738]), .A2(n7504), .B1(
        i_data_bus[706]), .B2(n7510), .ZN(n7452) );
  AOI22D1BWP30P140LVT U7995 ( .A1(i_data_bus[34]), .A2(n7514), .B1(
        i_data_bus[194]), .B2(n7502), .ZN(n7451) );
  AOI22D1BWP30P140LVT U7996 ( .A1(i_data_bus[866]), .A2(n7497), .B1(
        i_data_bus[834]), .B2(n7498), .ZN(n7450) );
  AN4D0BWP30P140LVT U7997 ( .A1(n7453), .A2(n7452), .A3(n7451), .A4(n7450), 
        .Z(n7469) );
  AOI22D1BWP30P140LVT U7998 ( .A1(i_data_bus[98]), .A2(n7512), .B1(
        i_data_bus[226]), .B2(n7501), .ZN(n7457) );
  AOI22D1BWP30P140LVT U7999 ( .A1(i_data_bus[2]), .A2(n7500), .B1(
        i_data_bus[642]), .B2(n7499), .ZN(n7456) );
  AOI22D1BWP30P140LVT U8000 ( .A1(i_data_bus[802]), .A2(n7513), .B1(
        i_data_bus[770]), .B2(n7516), .ZN(n7455) );
  AOI22D1BWP30P140LVT U8001 ( .A1(i_data_bus[66]), .A2(n7511), .B1(
        i_data_bus[674]), .B2(n7509), .ZN(n7454) );
  ND4D1BWP30P140LVT U8002 ( .A1(n7457), .A2(n7456), .A3(n7455), .A4(n7454), 
        .ZN(n7467) );
  INVD1BWP30P140LVT U8003 ( .I(i_data_bus[450]), .ZN(n7633) );
  INVD1BWP30P140LVT U8004 ( .I(i_data_bus[322]), .ZN(n9138) );
  OAI22D1BWP30P140LVT U8005 ( .A1(n7633), .A2(n7522), .B1(n9138), .B2(n7458), 
        .ZN(n7466) );
  INVD1BWP30P140LVT U8006 ( .I(i_data_bus[258]), .ZN(n9139) );
  MOAI22D1BWP30P140LVT U8007 ( .A1(n9139), .A2(n7521), .B1(i_data_bus[482]), 
        .B2(n7459), .ZN(n7465) );
  AOI22D1BWP30P140LVT U8008 ( .A1(i_data_bus[578]), .A2(n7531), .B1(
        i_data_bus[610]), .B2(n7529), .ZN(n7463) );
  AOI22D1BWP30P140LVT U8009 ( .A1(i_data_bus[546]), .A2(n7526), .B1(
        i_data_bus[898]), .B2(n7527), .ZN(n7462) );
  AOI22D1BWP30P140LVT U8010 ( .A1(i_data_bus[962]), .A2(n7525), .B1(
        i_data_bus[514]), .B2(n7530), .ZN(n7461) );
  AOI22D1BWP30P140LVT U8011 ( .A1(i_data_bus[994]), .A2(n7532), .B1(
        i_data_bus[930]), .B2(n7528), .ZN(n7460) );
  ND4D1BWP30P140LVT U8012 ( .A1(n7463), .A2(n7462), .A3(n7461), .A4(n7460), 
        .ZN(n7464) );
  NR4D0BWP30P140LVT U8013 ( .A1(n7467), .A2(n7466), .A3(n7465), .A4(n7464), 
        .ZN(n7468) );
  ND4D4BWP30P140LVT U8014 ( .A1(n7471), .A2(n7470), .A3(n7469), .A4(n7468), 
        .ZN(o_data_bus[66]) );
  AOI22D1BWP30P140LVT U8015 ( .A1(i_data_bus[449]), .A2(n7472), .B1(
        i_data_bus[417]), .B2(n7523), .ZN(n7492) );
  AOI22D1BWP30P140LVT U8016 ( .A1(i_data_bus[353]), .A2(n7495), .B1(
        i_data_bus[321]), .B2(n7493), .ZN(n7491) );
  AOI22D1BWP30P140LVT U8017 ( .A1(i_data_bus[97]), .A2(n7512), .B1(
        i_data_bus[705]), .B2(n7510), .ZN(n7476) );
  AOI22D1BWP30P140LVT U8018 ( .A1(i_data_bus[129]), .A2(n7503), .B1(
        i_data_bus[833]), .B2(n7498), .ZN(n7475) );
  AOI22D1BWP30P140LVT U8019 ( .A1(i_data_bus[161]), .A2(n7515), .B1(
        i_data_bus[225]), .B2(n7501), .ZN(n7474) );
  AOI22D1BWP30P140LVT U8020 ( .A1(i_data_bus[65]), .A2(n7511), .B1(
        i_data_bus[801]), .B2(n7513), .ZN(n7473) );
  AN4D0BWP30P140LVT U8021 ( .A1(n7476), .A2(n7475), .A3(n7474), .A4(n7473), 
        .Z(n7490) );
  AOI22D1BWP30P140LVT U8022 ( .A1(i_data_bus[769]), .A2(n7516), .B1(
        i_data_bus[673]), .B2(n7509), .ZN(n7480) );
  AOI22D1BWP30P140LVT U8023 ( .A1(i_data_bus[737]), .A2(n7504), .B1(
        i_data_bus[193]), .B2(n7502), .ZN(n7479) );
  AOI22D1BWP30P140LVT U8024 ( .A1(i_data_bus[1]), .A2(n7500), .B1(
        i_data_bus[865]), .B2(n7497), .ZN(n7478) );
  AOI22D1BWP30P140LVT U8025 ( .A1(i_data_bus[33]), .A2(n7514), .B1(
        i_data_bus[641]), .B2(n7499), .ZN(n7477) );
  ND4D1BWP30P140LVT U8026 ( .A1(n7480), .A2(n7479), .A3(n7478), .A4(n7477), 
        .ZN(n7488) );
  INVD1BWP30P140LVT U8027 ( .I(i_data_bus[257]), .ZN(n9054) );
  MOAI22D1BWP30P140LVT U8028 ( .A1(n9054), .A2(n7521), .B1(i_data_bus[289]), 
        .B2(n7494), .ZN(n7487) );
  INVD1BWP30P140LVT U8029 ( .I(i_data_bus[481]), .ZN(n8556) );
  MOAI22D1BWP30P140LVT U8030 ( .A1(n8556), .A2(n7524), .B1(i_data_bus[385]), 
        .B2(n7496), .ZN(n7486) );
  AOI22D1BWP30P140LVT U8031 ( .A1(i_data_bus[577]), .A2(n7531), .B1(
        i_data_bus[993]), .B2(n7532), .ZN(n7484) );
  AOI22D1BWP30P140LVT U8032 ( .A1(i_data_bus[897]), .A2(n7527), .B1(
        i_data_bus[513]), .B2(n7530), .ZN(n7483) );
  AOI22D1BWP30P140LVT U8033 ( .A1(i_data_bus[961]), .A2(n7525), .B1(
        i_data_bus[609]), .B2(n7529), .ZN(n7482) );
  AOI22D1BWP30P140LVT U8034 ( .A1(i_data_bus[545]), .A2(n7526), .B1(
        i_data_bus[929]), .B2(n7528), .ZN(n7481) );
  ND4D1BWP30P140LVT U8035 ( .A1(n7484), .A2(n7483), .A3(n7482), .A4(n7481), 
        .ZN(n7485) );
  NR4D0BWP30P140LVT U8036 ( .A1(n7488), .A2(n7487), .A3(n7486), .A4(n7485), 
        .ZN(n7489) );
  ND4D4BWP30P140LVT U8037 ( .A1(n7492), .A2(n7491), .A3(n7490), .A4(n7489), 
        .ZN(o_data_bus[65]) );
  AOI22D1BWP30P140LVT U8038 ( .A1(i_data_bus[288]), .A2(n7494), .B1(
        i_data_bus[320]), .B2(n7493), .ZN(n7544) );
  AOI22D1BWP30P140LVT U8039 ( .A1(i_data_bus[384]), .A2(n7496), .B1(
        i_data_bus[352]), .B2(n7495), .ZN(n7543) );
  AOI22D1BWP30P140LVT U8040 ( .A1(i_data_bus[832]), .A2(n7498), .B1(
        i_data_bus[864]), .B2(n7497), .ZN(n7508) );
  AOI22D1BWP30P140LVT U8041 ( .A1(i_data_bus[0]), .A2(n7500), .B1(
        i_data_bus[640]), .B2(n7499), .ZN(n7507) );
  AOI22D1BWP30P140LVT U8042 ( .A1(i_data_bus[192]), .A2(n7502), .B1(
        i_data_bus[224]), .B2(n7501), .ZN(n7506) );
  AOI22D1BWP30P140LVT U8043 ( .A1(i_data_bus[736]), .A2(n7504), .B1(
        i_data_bus[128]), .B2(n7503), .ZN(n7505) );
  AN4D0BWP30P140LVT U8044 ( .A1(n7508), .A2(n7507), .A3(n7506), .A4(n7505), 
        .Z(n7542) );
  AOI22D1BWP30P140LVT U8045 ( .A1(i_data_bus[704]), .A2(n7510), .B1(
        i_data_bus[672]), .B2(n7509), .ZN(n7520) );
  AOI22D1BWP30P140LVT U8046 ( .A1(i_data_bus[96]), .A2(n7512), .B1(
        i_data_bus[64]), .B2(n7511), .ZN(n7519) );
  AOI22D1BWP30P140LVT U8047 ( .A1(i_data_bus[32]), .A2(n7514), .B1(
        i_data_bus[800]), .B2(n7513), .ZN(n7518) );
  AOI22D1BWP30P140LVT U8048 ( .A1(i_data_bus[768]), .A2(n7516), .B1(
        i_data_bus[160]), .B2(n7515), .ZN(n7517) );
  ND4D1BWP30P140LVT U8049 ( .A1(n7520), .A2(n7519), .A3(n7518), .A4(n7517), 
        .ZN(n7540) );
  INVD1BWP30P140LVT U8050 ( .I(i_data_bus[448]), .ZN(n8715) );
  INVD1BWP30P140LVT U8051 ( .I(i_data_bus[256]), .ZN(n9182) );
  OAI22D1BWP30P140LVT U8052 ( .A1(n8715), .A2(n7522), .B1(n9182), .B2(n7521), 
        .ZN(n7539) );
  INVD1BWP30P140LVT U8053 ( .I(i_data_bus[480]), .ZN(n7691) );
  MOAI22D1BWP30P140LVT U8054 ( .A1(n7691), .A2(n7524), .B1(i_data_bus[416]), 
        .B2(n7523), .ZN(n7538) );
  AOI22D1BWP30P140LVT U8055 ( .A1(i_data_bus[544]), .A2(n7526), .B1(
        i_data_bus[960]), .B2(n7525), .ZN(n7536) );
  AOI22D1BWP30P140LVT U8056 ( .A1(i_data_bus[928]), .A2(n7528), .B1(
        i_data_bus[896]), .B2(n7527), .ZN(n7535) );
  AOI22D1BWP30P140LVT U8057 ( .A1(i_data_bus[512]), .A2(n7530), .B1(
        i_data_bus[608]), .B2(n7529), .ZN(n7534) );
  AOI22D1BWP30P140LVT U8058 ( .A1(i_data_bus[992]), .A2(n7532), .B1(
        i_data_bus[576]), .B2(n7531), .ZN(n7533) );
  ND4D1BWP30P140LVT U8059 ( .A1(n7536), .A2(n7535), .A3(n7534), .A4(n7533), 
        .ZN(n7537) );
  NR4D0BWP30P140LVT U8060 ( .A1(n7540), .A2(n7539), .A3(n7538), .A4(n7537), 
        .ZN(n7541) );
  ND4D4BWP30P140LVT U8061 ( .A1(n7544), .A2(n7543), .A3(n7542), .A4(n7541), 
        .ZN(o_data_bus[64]) );
  NR3D0P7BWP30P140LVT U8062 ( .A1(n11717), .A2(n7545), .A3(n7555), .ZN(n8702)
         );
  INR3D0BWP30P140LVT U8063 ( .A1(i_cmd[213]), .B1(n11745), .B2(n7558), .ZN(
        n8690) );
  AOI22D1BWP30P140LVT U8064 ( .A1(i_data_bus[1021]), .A2(n8702), .B1(
        i_data_bus[861]), .B2(n8690), .ZN(n7584) );
  NR3D0P7BWP30P140LVT U8065 ( .A1(n11740), .A2(n7546), .A3(n7555), .ZN(n8704)
         );
  INVD1BWP30P140LVT U8066 ( .I(i_cmd[197]), .ZN(n7547) );
  NR3D0P7BWP30P140LVT U8067 ( .A1(n11754), .A2(n7547), .A3(n7558), .ZN(n8707)
         );
  AOI22D1BWP30P140LVT U8068 ( .A1(i_data_bus[957]), .A2(n8704), .B1(
        i_data_bus[797]), .B2(n8707), .ZN(n7583) );
  ND3D1BWP30P140LVT U8069 ( .A1(i_valid[14]), .A2(i_cmd[117]), .A3(n7568), 
        .ZN(n8714) );
  INVD1BWP30P140LVT U8070 ( .I(n8714), .ZN(n8626) );
  ND3D1BWP30P140LVT U8071 ( .A1(i_valid[6]), .A2(i_cmd[53]), .A3(n7571), .ZN(
        n8623) );
  INVD1BWP30P140LVT U8072 ( .I(n8623), .ZN(n8713) );
  AOI22D1BWP30P140LVT U8073 ( .A1(i_data_bus[477]), .A2(n8626), .B1(
        i_data_bus[221]), .B2(n8713), .ZN(n7582) );
  INR3D0BWP30P140LVT U8074 ( .A1(i_cmd[29]), .B1(n11726), .B2(n7557), .ZN(
        n8692) );
  INR3D0BWP30P140LVT U8075 ( .A1(i_cmd[221]), .B1(n11749), .B2(n7558), .ZN(
        n8706) );
  AOI22D1BWP30P140LVT U8076 ( .A1(i_data_bus[125]), .A2(n8692), .B1(
        i_data_bus[893]), .B2(n8706), .ZN(n7553) );
  INVD1BWP30P140LVT U8077 ( .I(i_cmd[5]), .ZN(n7548) );
  NR3D0P7BWP30P140LVT U8078 ( .A1(n11703), .A2(n7548), .A3(n7557), .ZN(n8683)
         );
  INVD1BWP30P140LVT U8079 ( .I(i_valid[9]), .ZN(n11711) );
  INR3D0BWP30P140LVT U8080 ( .A1(i_cmd[77]), .B1(n11711), .B2(n7560), .ZN(
        n8705) );
  AOI22D1BWP30P140LVT U8081 ( .A1(i_data_bus[29]), .A2(n8683), .B1(
        i_data_bus[317]), .B2(n8705), .ZN(n7552) );
  NR3D0P7BWP30P140LVT U8082 ( .A1(n11715), .A2(n7549), .A3(n7555), .ZN(n8708)
         );
  INVD1BWP30P140LVT U8083 ( .I(i_valid[11]), .ZN(n11731) );
  INR3D0BWP30P140LVT U8084 ( .A1(i_cmd[93]), .B1(n11731), .B2(n7560), .ZN(
        n8701) );
  AOI22D1BWP30P140LVT U8085 ( .A1(i_data_bus[989]), .A2(n8708), .B1(
        i_data_bus[381]), .B2(n8701), .ZN(n7551) );
  INR3D0BWP30P140LVT U8086 ( .A1(i_cmd[173]), .B1(n11756), .B2(n7559), .ZN(
        n8689) );
  INR3D0BWP30P140LVT U8087 ( .A1(i_cmd[181]), .B1(n11748), .B2(n7559), .ZN(
        n8703) );
  AOI22D1BWP30P140LVT U8088 ( .A1(i_data_bus[701]), .A2(n8689), .B1(
        i_data_bus[733]), .B2(n8703), .ZN(n7550) );
  ND4D1BWP30P140LVT U8089 ( .A1(n7553), .A2(n7552), .A3(n7551), .A4(n7550), 
        .ZN(n7580) );
  INR3D0BWP30P140LVT U8090 ( .A1(i_cmd[13]), .B1(n11737), .B2(n7557), .ZN(
        n8684) );
  INVD1BWP30P140LVT U8091 ( .I(i_cmd[165]), .ZN(n7554) );
  NR3D0P7BWP30P140LVT U8092 ( .A1(n11747), .A2(n7554), .A3(n7559), .ZN(n8693)
         );
  AOI22D1BWP30P140LVT U8093 ( .A1(i_data_bus[61]), .A2(n8684), .B1(
        i_data_bus[669]), .B2(n8693), .ZN(n7565) );
  NR3D0P7BWP30P140LVT U8094 ( .A1(n11735), .A2(n7556), .A3(n7555), .ZN(n8686)
         );
  INVD1BWP30P140LVT U8095 ( .I(i_valid[10]), .ZN(n11700) );
  INR3D0BWP30P140LVT U8096 ( .A1(i_cmd[85]), .B1(n11700), .B2(n7560), .ZN(
        n8685) );
  AOI22D1BWP30P140LVT U8097 ( .A1(i_data_bus[925]), .A2(n8686), .B1(
        i_data_bus[349]), .B2(n8685), .ZN(n7564) );
  INR3D0BWP30P140LVT U8098 ( .A1(i_cmd[21]), .B1(n11699), .B2(n7557), .ZN(
        n8694) );
  INR3D0BWP30P140LVT U8099 ( .A1(i_cmd[205]), .B1(n11751), .B2(n7558), .ZN(
        n8695) );
  AOI22D1BWP30P140LVT U8100 ( .A1(i_data_bus[93]), .A2(n8694), .B1(
        i_data_bus[829]), .B2(n8695), .ZN(n7563) );
  INR3D0BWP30P140LVT U8101 ( .A1(i_cmd[189]), .B1(n11750), .B2(n7559), .ZN(
        n8696) );
  INVD1BWP30P140LVT U8102 ( .I(i_valid[8]), .ZN(n11728) );
  NR3D0P7BWP30P140LVT U8103 ( .A1(n11728), .A2(n7561), .A3(n7560), .ZN(n8691)
         );
  AOI22D1BWP30P140LVT U8104 ( .A1(i_data_bus[765]), .A2(n8696), .B1(
        i_data_bus[285]), .B2(n8691), .ZN(n7562) );
  ND4D1BWP30P140LVT U8105 ( .A1(n7565), .A2(n7564), .A3(n7563), .A4(n7562), 
        .ZN(n7579) );
  ND3D1BWP30P140LVT U8106 ( .A1(i_valid[15]), .A2(i_cmd[125]), .A3(n7568), 
        .ZN(n8624) );
  INR3D0BWP30P140LVT U8107 ( .A1(n7568), .B1(n7566), .B2(n11705), .ZN(n8719)
         );
  MOAI22D1BWP30P140LVT U8108 ( .A1(n7567), .A2(n8624), .B1(i_data_bus[413]), 
        .B2(n8719), .ZN(n7578) );
  AN3D1BWP30P140LVT U8109 ( .A1(i_valid[13]), .A2(i_cmd[109]), .A3(n7568), .Z(
        n8717) );
  ND3D1BWP30P140LVT U8110 ( .A1(i_valid[5]), .A2(i_cmd[45]), .A3(n7571), .ZN(
        n8602) );
  INVD1BWP30P140LVT U8111 ( .I(n8602), .ZN(n8716) );
  AOI22D1BWP30P140LVT U8112 ( .A1(i_data_bus[445]), .A2(n8717), .B1(
        i_data_bus[189]), .B2(n8716), .ZN(n7576) );
  INVD1BWP30P140LVT U8113 ( .I(i_cmd[37]), .ZN(n7570) );
  NR3D0P7BWP30P140LVT U8114 ( .A1(n11721), .A2(n7570), .A3(n7569), .ZN(n8688)
         );
  AN3D1BWP30P140LVT U8115 ( .A1(i_cmd[61]), .A2(i_valid[7]), .A3(n7571), .Z(
        n8687) );
  AOI22D1BWP30P140LVT U8116 ( .A1(i_data_bus[157]), .A2(n8688), .B1(
        i_data_bus[253]), .B2(n8687), .ZN(n7575) );
  INR3D0BWP30P140LVT U8117 ( .A1(i_cmd[141]), .B1(n11701), .B2(n7572), .ZN(
        n8723) );
  NR3D0P7BWP30P140LVT U8118 ( .A1(n11713), .A2(n6492), .A3(n7572), .ZN(n8721)
         );
  AOI22D1BWP30P140LVT U8119 ( .A1(i_data_bus[573]), .A2(n8723), .B1(
        i_data_bus[541]), .B2(n8721), .ZN(n7574) );
  INR3D0BWP30P140LVT U8120 ( .A1(i_cmd[157]), .B1(n11697), .B2(n7572), .ZN(
        n8720) );
  INR3D0BWP30P140LVT U8121 ( .A1(i_cmd[149]), .B1(n11733), .B2(n7572), .ZN(
        n8722) );
  AOI22D1BWP30P140LVT U8122 ( .A1(i_data_bus[637]), .A2(n8720), .B1(
        i_data_bus[605]), .B2(n8722), .ZN(n7573) );
  ND4D1BWP30P140LVT U8123 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), 
        .ZN(n7577) );
  NR4D0BWP30P140LVT U8124 ( .A1(n7580), .A2(n7579), .A3(n7578), .A4(n7577), 
        .ZN(n7581) );
  ND4D4BWP30P140LVT U8125 ( .A1(n7584), .A2(n7583), .A3(n7582), .A4(n7581), 
        .ZN(o_data_bus[189]) );
  AOI22D1BWP30P140LVT U8126 ( .A1(i_data_bus[936]), .A2(n8704), .B1(
        i_data_bus[808]), .B2(n8695), .ZN(n7604) );
  AOI22D1BWP30P140LVT U8127 ( .A1(i_data_bus[904]), .A2(n8686), .B1(
        i_data_bus[40]), .B2(n8684), .ZN(n7603) );
  INVD1BWP30P140LVT U8128 ( .I(n8624), .ZN(n8718) );
  AOI22D1BWP30P140LVT U8129 ( .A1(i_data_bus[456]), .A2(n8626), .B1(
        i_data_bus[488]), .B2(n8718), .ZN(n7602) );
  AOI22D1BWP30P140LVT U8130 ( .A1(i_data_bus[200]), .A2(n8713), .B1(
        i_data_bus[136]), .B2(n8688), .ZN(n7600) );
  AOI22D1BWP30P140LVT U8131 ( .A1(i_data_bus[104]), .A2(n8692), .B1(
        i_data_bus[1000]), .B2(n8702), .ZN(n7588) );
  AOI22D1BWP30P140LVT U8132 ( .A1(i_data_bus[72]), .A2(n8694), .B1(
        i_data_bus[712]), .B2(n8703), .ZN(n7587) );
  AOI22D1BWP30P140LVT U8133 ( .A1(i_data_bus[840]), .A2(n8690), .B1(
        i_data_bus[648]), .B2(n8693), .ZN(n7586) );
  AOI22D1BWP30P140LVT U8134 ( .A1(i_data_bus[968]), .A2(n8708), .B1(
        i_data_bus[328]), .B2(n8685), .ZN(n7585) );
  ND4D1BWP30P140LVT U8135 ( .A1(n7588), .A2(n7587), .A3(n7586), .A4(n7585), 
        .ZN(n7599) );
  AOI22D1BWP30P140LVT U8136 ( .A1(i_data_bus[8]), .A2(n8683), .B1(
        i_data_bus[776]), .B2(n8707), .ZN(n7592) );
  AOI22D1BWP30P140LVT U8137 ( .A1(i_data_bus[744]), .A2(n8696), .B1(
        i_data_bus[680]), .B2(n8689), .ZN(n7591) );
  AOI22D1BWP30P140LVT U8138 ( .A1(i_data_bus[264]), .A2(n8691), .B1(
        i_data_bus[872]), .B2(n8706), .ZN(n7590) );
  AOI22D1BWP30P140LVT U8139 ( .A1(i_data_bus[296]), .A2(n8705), .B1(
        i_data_bus[360]), .B2(n8701), .ZN(n7589) );
  ND4D1BWP30P140LVT U8140 ( .A1(n7592), .A2(n7591), .A3(n7590), .A4(n7589), 
        .ZN(n7598) );
  AOI22D1BWP30P140LVT U8141 ( .A1(i_data_bus[424]), .A2(n8717), .B1(
        i_data_bus[392]), .B2(n8719), .ZN(n7596) );
  AOI22D1BWP30P140LVT U8142 ( .A1(i_data_bus[168]), .A2(n8716), .B1(
        i_data_bus[232]), .B2(n8687), .ZN(n7595) );
  AOI22D1BWP30P140LVT U8143 ( .A1(i_data_bus[616]), .A2(n8720), .B1(
        i_data_bus[552]), .B2(n8723), .ZN(n7594) );
  AOI22D1BWP30P140LVT U8144 ( .A1(i_data_bus[584]), .A2(n8722), .B1(
        i_data_bus[520]), .B2(n8721), .ZN(n7593) );
  ND4D1BWP30P140LVT U8145 ( .A1(n7596), .A2(n7595), .A3(n7594), .A4(n7593), 
        .ZN(n7597) );
  INR4D0BWP30P140LVT U8146 ( .A1(n7600), .B1(n7599), .B2(n7598), .B3(n7597), 
        .ZN(n7601) );
  ND4D4BWP30P140LVT U8147 ( .A1(n7604), .A2(n7603), .A3(n7602), .A4(n7601), 
        .ZN(o_data_bus[168]) );
  AOI22D1BWP30P140LVT U8148 ( .A1(i_data_bus[731]), .A2(n8703), .B1(
        i_data_bus[827]), .B2(n8695), .ZN(n7624) );
  AOI22D1BWP30P140LVT U8149 ( .A1(i_data_bus[91]), .A2(n8694), .B1(
        i_data_bus[347]), .B2(n8685), .ZN(n7623) );
  AOI22D1BWP30P140LVT U8150 ( .A1(i_data_bus[507]), .A2(n8718), .B1(
        i_data_bus[251]), .B2(n8687), .ZN(n7622) );
  AOI22D1BWP30P140LVT U8151 ( .A1(i_data_bus[315]), .A2(n8705), .B1(
        i_data_bus[795]), .B2(n8707), .ZN(n7608) );
  AOI22D1BWP30P140LVT U8152 ( .A1(i_data_bus[987]), .A2(n8708), .B1(
        i_data_bus[1019]), .B2(n8702), .ZN(n7607) );
  AOI22D1BWP30P140LVT U8153 ( .A1(i_data_bus[667]), .A2(n8693), .B1(
        i_data_bus[699]), .B2(n8689), .ZN(n7606) );
  AOI22D1BWP30P140LVT U8154 ( .A1(i_data_bus[379]), .A2(n8701), .B1(
        i_data_bus[859]), .B2(n8690), .ZN(n7605) );
  ND4D1BWP30P140LVT U8155 ( .A1(n7608), .A2(n7607), .A3(n7606), .A4(n7605), 
        .ZN(n7620) );
  AOI22D1BWP30P140LVT U8156 ( .A1(i_data_bus[123]), .A2(n8692), .B1(
        i_data_bus[283]), .B2(n8691), .ZN(n7612) );
  AOI22D1BWP30P140LVT U8157 ( .A1(i_data_bus[923]), .A2(n8686), .B1(
        i_data_bus[59]), .B2(n8684), .ZN(n7611) );
  AOI22D1BWP30P140LVT U8158 ( .A1(i_data_bus[955]), .A2(n8704), .B1(
        i_data_bus[891]), .B2(n8706), .ZN(n7610) );
  AOI22D1BWP30P140LVT U8159 ( .A1(i_data_bus[27]), .A2(n8683), .B1(
        i_data_bus[763]), .B2(n8696), .ZN(n7609) );
  ND4D1BWP30P140LVT U8160 ( .A1(n7612), .A2(n7611), .A3(n7610), .A4(n7609), 
        .ZN(n7619) );
  INVD1BWP30P140LVT U8161 ( .I(i_data_bus[187]), .ZN(n7712) );
  MOAI22D1BWP30P140LVT U8162 ( .A1(n7712), .A2(n8602), .B1(i_data_bus[219]), 
        .B2(n8713), .ZN(n7618) );
  AOI22D1BWP30P140LVT U8163 ( .A1(i_data_bus[411]), .A2(n8719), .B1(
        i_data_bus[443]), .B2(n8717), .ZN(n7616) );
  AOI22D1BWP30P140LVT U8164 ( .A1(i_data_bus[155]), .A2(n8688), .B1(
        i_data_bus[475]), .B2(n8626), .ZN(n7615) );
  AOI22D1BWP30P140LVT U8165 ( .A1(i_data_bus[539]), .A2(n8721), .B1(
        i_data_bus[635]), .B2(n8720), .ZN(n7614) );
  AOI22D1BWP30P140LVT U8166 ( .A1(i_data_bus[571]), .A2(n8723), .B1(
        i_data_bus[603]), .B2(n8722), .ZN(n7613) );
  ND4D1BWP30P140LVT U8167 ( .A1(n7616), .A2(n7615), .A3(n7614), .A4(n7613), 
        .ZN(n7617) );
  NR4D0BWP30P140LVT U8168 ( .A1(n7620), .A2(n7619), .A3(n7618), .A4(n7617), 
        .ZN(n7621) );
  ND4D4BWP30P140LVT U8169 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), 
        .ZN(o_data_bus[187]) );
  AOI22D1BWP30P140LVT U8170 ( .A1(i_data_bus[962]), .A2(n8708), .B1(
        i_data_bus[258]), .B2(n8691), .ZN(n7645) );
  AOI22D1BWP30P140LVT U8171 ( .A1(i_data_bus[898]), .A2(n8686), .B1(
        i_data_bus[2]), .B2(n8683), .ZN(n7644) );
  AOI22D1BWP30P140LVT U8172 ( .A1(i_data_bus[482]), .A2(n8718), .B1(
        i_data_bus[418]), .B2(n8717), .ZN(n7643) );
  AOI22D1BWP30P140LVT U8173 ( .A1(i_data_bus[994]), .A2(n8702), .B1(
        i_data_bus[706]), .B2(n8703), .ZN(n7628) );
  AOI22D1BWP30P140LVT U8174 ( .A1(i_data_bus[98]), .A2(n8692), .B1(
        i_data_bus[674]), .B2(n8689), .ZN(n7627) );
  AOI22D1BWP30P140LVT U8175 ( .A1(i_data_bus[66]), .A2(n8694), .B1(
        i_data_bus[322]), .B2(n8685), .ZN(n7626) );
  AOI22D1BWP30P140LVT U8176 ( .A1(i_data_bus[290]), .A2(n8705), .B1(
        i_data_bus[642]), .B2(n8693), .ZN(n7625) );
  ND4D1BWP30P140LVT U8177 ( .A1(n7628), .A2(n7627), .A3(n7626), .A4(n7625), 
        .ZN(n7641) );
  AOI22D1BWP30P140LVT U8178 ( .A1(i_data_bus[930]), .A2(n8704), .B1(
        i_data_bus[770]), .B2(n8707), .ZN(n7632) );
  AOI22D1BWP30P140LVT U8179 ( .A1(i_data_bus[834]), .A2(n8690), .B1(
        i_data_bus[738]), .B2(n8696), .ZN(n7631) );
  AOI22D1BWP30P140LVT U8180 ( .A1(i_data_bus[802]), .A2(n8695), .B1(
        i_data_bus[354]), .B2(n8701), .ZN(n7630) );
  AOI22D1BWP30P140LVT U8181 ( .A1(i_data_bus[34]), .A2(n8684), .B1(
        i_data_bus[866]), .B2(n8706), .ZN(n7629) );
  ND4D1BWP30P140LVT U8182 ( .A1(n7632), .A2(n7631), .A3(n7630), .A4(n7629), 
        .ZN(n7640) );
  INVD1BWP30P140LVT U8183 ( .I(i_data_bus[194]), .ZN(n8391) );
  OAI22D1BWP30P140LVT U8184 ( .A1(n8391), .A2(n8623), .B1(n7633), .B2(n8714), 
        .ZN(n7639) );
  AOI22D1BWP30P140LVT U8185 ( .A1(i_data_bus[226]), .A2(n8687), .B1(
        i_data_bus[130]), .B2(n8688), .ZN(n7637) );
  AOI22D1BWP30P140LVT U8186 ( .A1(i_data_bus[162]), .A2(n8716), .B1(
        i_data_bus[386]), .B2(n8719), .ZN(n7636) );
  AOI22D1BWP30P140LVT U8187 ( .A1(i_data_bus[546]), .A2(n8723), .B1(
        i_data_bus[610]), .B2(n8720), .ZN(n7635) );
  AOI22D1BWP30P140LVT U8188 ( .A1(i_data_bus[578]), .A2(n8722), .B1(
        i_data_bus[514]), .B2(n8721), .ZN(n7634) );
  ND4D1BWP30P140LVT U8189 ( .A1(n7637), .A2(n7636), .A3(n7635), .A4(n7634), 
        .ZN(n7638) );
  NR4D0BWP30P140LVT U8190 ( .A1(n7641), .A2(n7640), .A3(n7639), .A4(n7638), 
        .ZN(n7642) );
  ND4D4BWP30P140LVT U8191 ( .A1(n7645), .A2(n7644), .A3(n7643), .A4(n7642), 
        .ZN(o_data_bus[162]) );
  INR3D0BWP30P140LVT U8192 ( .A1(i_cmd[191]), .B1(n11750), .B2(n7651), .ZN(
        n9546) );
  INR3D0BWP30P140LVT U8193 ( .A1(i_cmd[223]), .B1(n11749), .B2(n7650), .ZN(
        n9556) );
  AOI22D1BWP30P140LVT U8194 ( .A1(i_data_bus[761]), .A2(n9546), .B1(
        i_data_bus[889]), .B2(n9556), .ZN(n7686) );
  NR3D0P7BWP30P140LVT U8195 ( .A1(n7654), .A2(n11737), .A3(n7646), .ZN(n9548)
         );
  NR3D0P7BWP30P140LVT U8196 ( .A1(n7654), .A2(n7647), .A3(n11726), .ZN(n9555)
         );
  AOI22D1BWP30P140LVT U8197 ( .A1(i_data_bus[57]), .A2(n9548), .B1(
        i_data_bus[121]), .B2(n9555), .ZN(n7685) );
  ND3D1BWP30P140LVT U8198 ( .A1(i_valid[11]), .A2(i_cmd[95]), .A3(n7669), .ZN(
        n9375) );
  INVD1BWP30P140LVT U8199 ( .I(n9375), .ZN(n9569) );
  ND3D1BWP30P140LVT U8200 ( .A1(i_valid[9]), .A2(i_cmd[79]), .A3(n7669), .ZN(
        n9461) );
  INVD1BWP30P140LVT U8201 ( .I(n9461), .ZN(n9584) );
  AOI22D1BWP30P140LVT U8202 ( .A1(i_data_bus[377]), .A2(n9569), .B1(
        i_data_bus[313]), .B2(n9584), .ZN(n7684) );
  INVD1BWP30P140LVT U8203 ( .I(i_cmd[167]), .ZN(n7648) );
  NR3D0P7BWP30P140LVT U8204 ( .A1(n11747), .A2(n7648), .A3(n7651), .ZN(n9558)
         );
  NR3D0P7BWP30P140LVT U8205 ( .A1(n11754), .A2(n7649), .A3(n7650), .ZN(n9547)
         );
  AOI22D1BWP30P140LVT U8206 ( .A1(i_data_bus[665]), .A2(n9558), .B1(
        i_data_bus[793]), .B2(n9547), .ZN(n7658) );
  INR3D0BWP30P140LVT U8207 ( .A1(i_cmd[207]), .B1(n11751), .B2(n7650), .ZN(
        n9552) );
  INR3D0BWP30P140LVT U8208 ( .A1(i_cmd[215]), .B1(n11745), .B2(n7650), .ZN(
        n9557) );
  AOI22D1BWP30P140LVT U8209 ( .A1(i_data_bus[825]), .A2(n9552), .B1(
        i_data_bus[857]), .B2(n9557), .ZN(n7657) );
  INR3D0BWP30P140LVT U8210 ( .A1(i_cmd[183]), .B1(n11748), .B2(n7651), .ZN(
        n9554) );
  INR3D0BWP30P140LVT U8211 ( .A1(i_cmd[175]), .B1(n11756), .B2(n7651), .ZN(
        n9559) );
  AOI22D1BWP30P140LVT U8212 ( .A1(i_data_bus[729]), .A2(n9554), .B1(
        i_data_bus[697]), .B2(n9559), .ZN(n7656) );
  NR3D0P7BWP30P140LVT U8213 ( .A1(n7654), .A2(n11703), .A3(n7652), .ZN(n9553)
         );
  NR3D0P7BWP30P140LVT U8214 ( .A1(n7654), .A2(n7653), .A3(n11699), .ZN(n9549)
         );
  AOI22D1BWP30P140LVT U8215 ( .A1(i_data_bus[25]), .A2(n9553), .B1(
        i_data_bus[89]), .B2(n9549), .ZN(n7655) );
  ND4D1BWP30P140LVT U8216 ( .A1(n7658), .A2(n7657), .A3(n7656), .A4(n7655), 
        .ZN(n7682) );
  INVD1BWP30P140LVT U8217 ( .I(i_cmd[103]), .ZN(n7660) );
  NR3D0P7BWP30P140LVT U8218 ( .A1(n11705), .A2(n7660), .A3(n7659), .ZN(n9585)
         );
  INVD1BWP30P140LVT U8219 ( .I(n9585), .ZN(n9245) );
  INR3D0BWP30P140LVT U8220 ( .A1(i_cmd[255]), .B1(n11717), .B2(n7673), .ZN(
        n9571) );
  MOAI22D1BWP30P140LVT U8221 ( .A1(n8581), .A2(n9245), .B1(i_data_bus[1017]), 
        .B2(n9571), .ZN(n7681) );
  NR3D0P7BWP30P140LVT U8222 ( .A1(n11735), .A2(n7661), .A3(n7673), .ZN(n9581)
         );
  INR3D0BWP30P140LVT U8223 ( .A1(i_cmd[247]), .B1(n11715), .B2(n7673), .ZN(
        n9551) );
  AOI22D1BWP30P140LVT U8224 ( .A1(i_data_bus[921]), .A2(n9581), .B1(
        i_data_bus[985]), .B2(n9551), .ZN(n7668) );
  NR3D0P7BWP30P140LVT U8225 ( .A1(n11721), .A2(n7662), .A3(n7674), .ZN(n9533)
         );
  INR3D0BWP30P140LVT U8226 ( .A1(i_cmd[55]), .B1(n7674), .B2(n11030), .ZN(
        n9550) );
  AOI22D1BWP30P140LVT U8227 ( .A1(i_data_bus[153]), .A2(n9533), .B1(
        i_data_bus[217]), .B2(n9550), .ZN(n7667) );
  INR3D0BWP30P140LVT U8228 ( .A1(i_cmd[143]), .B1(n11701), .B2(n7664), .ZN(
        n9575) );
  INVD1BWP30P140LVT U8229 ( .I(i_cmd[135]), .ZN(n7663) );
  NR3D0P7BWP30P140LVT U8230 ( .A1(n11713), .A2(n7663), .A3(n7664), .ZN(n9573)
         );
  AOI22D1BWP30P140LVT U8231 ( .A1(i_data_bus[569]), .A2(n9575), .B1(
        i_data_bus[537]), .B2(n9573), .ZN(n7666) );
  INR3D0BWP30P140LVT U8232 ( .A1(i_cmd[159]), .B1(n11697), .B2(n7664), .ZN(
        n9574) );
  INR3D0BWP30P140LVT U8233 ( .A1(i_cmd[151]), .B1(n11733), .B2(n7664), .ZN(
        n9572) );
  AOI22D1BWP30P140LVT U8234 ( .A1(i_data_bus[633]), .A2(n9574), .B1(
        i_data_bus[601]), .B2(n9572), .ZN(n7665) );
  ND4D1BWP30P140LVT U8235 ( .A1(n7668), .A2(n7667), .A3(n7666), .A4(n7665), 
        .ZN(n7680) );
  ND3D1BWP30P140LVT U8236 ( .A1(i_valid[10]), .A2(i_cmd[87]), .A3(n7669), .ZN(
        n9247) );
  INVD1BWP30P140LVT U8237 ( .I(n9247), .ZN(n9570) );
  INVD1BWP30P140LVT U8238 ( .I(i_cmd[71]), .ZN(n7671) );
  NR3D0P7BWP30P140LVT U8239 ( .A1(n11728), .A2(n7671), .A3(n7670), .ZN(n9586)
         );
  AOI22D1BWP30P140LVT U8240 ( .A1(i_data_bus[345]), .A2(n9570), .B1(
        i_data_bus[281]), .B2(n9586), .ZN(n7678) );
  INR3D0BWP30P140LVT U8241 ( .A1(i_cmd[47]), .B1(n7674), .B2(n11023), .ZN(
        n9583) );
  ND3D1BWP30P140LVT U8242 ( .A1(i_valid[13]), .A2(i_cmd[111]), .A3(n7672), 
        .ZN(n9566) );
  INVD1BWP30P140LVT U8243 ( .I(n9566), .ZN(n9532) );
  AOI22D1BWP30P140LVT U8244 ( .A1(i_data_bus[185]), .A2(n9583), .B1(
        i_data_bus[441]), .B2(n9532), .ZN(n7677) );
  ND3D1BWP30P140LVT U8245 ( .A1(i_valid[14]), .A2(i_cmd[119]), .A3(n7672), 
        .ZN(n9526) );
  INVD1BWP30P140LVT U8246 ( .I(n9526), .ZN(n9582) );
  ND3D1BWP30P140LVT U8247 ( .A1(i_valid[15]), .A2(i_cmd[127]), .A3(n7672), 
        .ZN(n9397) );
  INVD1BWP30P140LVT U8248 ( .I(n9397), .ZN(n9580) );
  AOI22D1BWP30P140LVT U8249 ( .A1(i_data_bus[473]), .A2(n9582), .B1(
        i_data_bus[505]), .B2(n9580), .ZN(n7676) );
  INR3D0BWP30P140LVT U8250 ( .A1(i_cmd[239]), .B1(n11740), .B2(n7673), .ZN(
        n9587) );
  INR3D0BWP30P140LVT U8251 ( .A1(i_cmd[63]), .B1(n11032), .B2(n7674), .ZN(
        n9568) );
  AOI22D1BWP30P140LVT U8252 ( .A1(i_data_bus[953]), .A2(n9587), .B1(
        i_data_bus[249]), .B2(n9568), .ZN(n7675) );
  ND4D1BWP30P140LVT U8253 ( .A1(n7678), .A2(n7677), .A3(n7676), .A4(n7675), 
        .ZN(n7679) );
  NR4D0BWP30P140LVT U8254 ( .A1(n7682), .A2(n7681), .A3(n7680), .A4(n7679), 
        .ZN(n7683) );
  ND4D4BWP30P140LVT U8255 ( .A1(n7686), .A2(n7685), .A3(n7684), .A4(n7683), 
        .ZN(o_data_bus[249]) );
  AOI22D1BWP30P140LVT U8256 ( .A1(i_data_bus[32]), .A2(n9548), .B1(
        i_data_bus[768]), .B2(n9547), .ZN(n7707) );
  AOI22D1BWP30P140LVT U8257 ( .A1(i_data_bus[96]), .A2(n9555), .B1(
        i_data_bus[704]), .B2(n9554), .ZN(n7706) );
  AOI22D1BWP30P140LVT U8258 ( .A1(i_data_bus[352]), .A2(n9569), .B1(
        i_data_bus[320]), .B2(n9570), .ZN(n7705) );
  AOI22D1BWP30P140LVT U8259 ( .A1(i_data_bus[0]), .A2(n9553), .B1(
        i_data_bus[64]), .B2(n9549), .ZN(n7690) );
  AOI22D1BWP30P140LVT U8260 ( .A1(i_data_bus[640]), .A2(n9558), .B1(
        i_data_bus[864]), .B2(n9556), .ZN(n7689) );
  AOI22D1BWP30P140LVT U8261 ( .A1(i_data_bus[736]), .A2(n9546), .B1(
        i_data_bus[800]), .B2(n9552), .ZN(n7688) );
  AOI22D1BWP30P140LVT U8262 ( .A1(i_data_bus[832]), .A2(n9557), .B1(
        i_data_bus[672]), .B2(n9559), .ZN(n7687) );
  ND4D1BWP30P140LVT U8263 ( .A1(n7690), .A2(n7689), .A3(n7688), .A4(n7687), 
        .ZN(n7703) );
  MOAI22D1BWP30P140LVT U8264 ( .A1(n7691), .A2(n9397), .B1(i_data_bus[288]), 
        .B2(n9584), .ZN(n7702) );
  AOI22D1BWP30P140LVT U8265 ( .A1(i_data_bus[992]), .A2(n9571), .B1(
        i_data_bus[224]), .B2(n9568), .ZN(n7695) );
  AOI22D1BWP30P140LVT U8266 ( .A1(i_data_bus[896]), .A2(n9581), .B1(
        i_data_bus[384]), .B2(n9585), .ZN(n7694) );
  AOI22D1BWP30P140LVT U8267 ( .A1(i_data_bus[512]), .A2(n9573), .B1(
        i_data_bus[608]), .B2(n9574), .ZN(n7693) );
  AOI22D1BWP30P140LVT U8268 ( .A1(i_data_bus[544]), .A2(n9575), .B1(
        i_data_bus[576]), .B2(n9572), .ZN(n7692) );
  ND4D1BWP30P140LVT U8269 ( .A1(n7695), .A2(n7694), .A3(n7693), .A4(n7692), 
        .ZN(n7701) );
  AOI22D1BWP30P140LVT U8270 ( .A1(i_data_bus[928]), .A2(n9587), .B1(
        i_data_bus[160]), .B2(n9583), .ZN(n7699) );
  AOI22D1BWP30P140LVT U8271 ( .A1(i_data_bus[960]), .A2(n9551), .B1(
        i_data_bus[416]), .B2(n9532), .ZN(n7698) );
  AOI22D1BWP30P140LVT U8272 ( .A1(i_data_bus[448]), .A2(n9582), .B1(
        i_data_bus[128]), .B2(n9533), .ZN(n7697) );
  AOI22D1BWP30P140LVT U8273 ( .A1(i_data_bus[192]), .A2(n9550), .B1(
        i_data_bus[256]), .B2(n9586), .ZN(n7696) );
  ND4D1BWP30P140LVT U8274 ( .A1(n7699), .A2(n7698), .A3(n7697), .A4(n7696), 
        .ZN(n7700) );
  NR4D0BWP30P140LVT U8275 ( .A1(n7703), .A2(n7702), .A3(n7701), .A4(n7700), 
        .ZN(n7704) );
  ND4D4BWP30P140LVT U8276 ( .A1(n7707), .A2(n7706), .A3(n7705), .A4(n7704), 
        .ZN(o_data_bus[224]) );
  AOI22D1BWP30P140LVT U8277 ( .A1(i_data_bus[59]), .A2(n9548), .B1(
        i_data_bus[827]), .B2(n9552), .ZN(n7729) );
  AOI22D1BWP30P140LVT U8278 ( .A1(i_data_bus[123]), .A2(n9555), .B1(
        i_data_bus[859]), .B2(n9557), .ZN(n7728) );
  AOI22D1BWP30P140LVT U8279 ( .A1(i_data_bus[507]), .A2(n9580), .B1(
        i_data_bus[155]), .B2(n9533), .ZN(n7727) );
  AOI22D1BWP30P140LVT U8280 ( .A1(i_data_bus[91]), .A2(n9549), .B1(
        i_data_bus[731]), .B2(n9554), .ZN(n7711) );
  AOI22D1BWP30P140LVT U8281 ( .A1(i_data_bus[667]), .A2(n9558), .B1(
        i_data_bus[699]), .B2(n9559), .ZN(n7710) );
  AOI22D1BWP30P140LVT U8282 ( .A1(i_data_bus[27]), .A2(n9553), .B1(
        i_data_bus[795]), .B2(n9547), .ZN(n7709) );
  AOI22D1BWP30P140LVT U8283 ( .A1(i_data_bus[891]), .A2(n9556), .B1(
        i_data_bus[763]), .B2(n9546), .ZN(n7708) );
  ND4D1BWP30P140LVT U8284 ( .A1(n7711), .A2(n7710), .A3(n7709), .A4(n7708), 
        .ZN(n7725) );
  INVD1BWP30P140LVT U8285 ( .I(n9583), .ZN(n9419) );
  OAI22D1BWP30P140LVT U8286 ( .A1(n7713), .A2(n9247), .B1(n7712), .B2(n9419), 
        .ZN(n7724) );
  AOI22D1BWP30P140LVT U8287 ( .A1(i_data_bus[219]), .A2(n9550), .B1(
        i_data_bus[283]), .B2(n9586), .ZN(n7717) );
  AOI22D1BWP30P140LVT U8288 ( .A1(i_data_bus[1019]), .A2(n9571), .B1(
        i_data_bus[379]), .B2(n9569), .ZN(n7716) );
  AOI22D1BWP30P140LVT U8289 ( .A1(i_data_bus[571]), .A2(n9575), .B1(
        i_data_bus[539]), .B2(n9573), .ZN(n7715) );
  AOI22D1BWP30P140LVT U8290 ( .A1(i_data_bus[603]), .A2(n9572), .B1(
        i_data_bus[635]), .B2(n9574), .ZN(n7714) );
  ND4D1BWP30P140LVT U8291 ( .A1(n7717), .A2(n7716), .A3(n7715), .A4(n7714), 
        .ZN(n7723) );
  AOI22D1BWP30P140LVT U8292 ( .A1(i_data_bus[315]), .A2(n9584), .B1(
        i_data_bus[475]), .B2(n9582), .ZN(n7721) );
  AOI22D1BWP30P140LVT U8293 ( .A1(i_data_bus[987]), .A2(n9551), .B1(
        i_data_bus[443]), .B2(n9532), .ZN(n7720) );
  AOI22D1BWP30P140LVT U8294 ( .A1(i_data_bus[411]), .A2(n9585), .B1(
        i_data_bus[251]), .B2(n9568), .ZN(n7719) );
  AOI22D1BWP30P140LVT U8295 ( .A1(i_data_bus[923]), .A2(n9581), .B1(
        i_data_bus[955]), .B2(n9587), .ZN(n7718) );
  ND4D1BWP30P140LVT U8296 ( .A1(n7721), .A2(n7720), .A3(n7719), .A4(n7718), 
        .ZN(n7722) );
  NR4D0BWP30P140LVT U8297 ( .A1(n7725), .A2(n7724), .A3(n7723), .A4(n7722), 
        .ZN(n7726) );
  ND4D4BWP30P140LVT U8298 ( .A1(n7729), .A2(n7728), .A3(n7727), .A4(n7726), 
        .ZN(o_data_bus[251]) );
  AOI22D1BWP30P140LVT U8299 ( .A1(i_data_bus[874]), .A2(n8706), .B1(
        i_data_bus[714]), .B2(n8703), .ZN(n7749) );
  AOI22D1BWP30P140LVT U8300 ( .A1(i_data_bus[362]), .A2(n8701), .B1(
        i_data_bus[810]), .B2(n8695), .ZN(n7748) );
  AOI22D1BWP30P140LVT U8301 ( .A1(i_data_bus[490]), .A2(n8718), .B1(
        i_data_bus[138]), .B2(n8688), .ZN(n7747) );
  AOI22D1BWP30P140LVT U8302 ( .A1(i_data_bus[106]), .A2(n8692), .B1(
        i_data_bus[74]), .B2(n8694), .ZN(n7733) );
  AOI22D1BWP30P140LVT U8303 ( .A1(i_data_bus[970]), .A2(n8708), .B1(
        i_data_bus[266]), .B2(n8691), .ZN(n7732) );
  AOI22D1BWP30P140LVT U8304 ( .A1(i_data_bus[778]), .A2(n8707), .B1(
        i_data_bus[842]), .B2(n8690), .ZN(n7731) );
  AOI22D1BWP30P140LVT U8305 ( .A1(i_data_bus[1002]), .A2(n8702), .B1(
        i_data_bus[42]), .B2(n8684), .ZN(n7730) );
  ND4D1BWP30P140LVT U8306 ( .A1(n7733), .A2(n7732), .A3(n7731), .A4(n7730), 
        .ZN(n7745) );
  AOI22D1BWP30P140LVT U8307 ( .A1(i_data_bus[938]), .A2(n8704), .B1(
        i_data_bus[330]), .B2(n8685), .ZN(n7737) );
  AOI22D1BWP30P140LVT U8308 ( .A1(i_data_bus[650]), .A2(n8693), .B1(
        i_data_bus[298]), .B2(n8705), .ZN(n7736) );
  AOI22D1BWP30P140LVT U8309 ( .A1(i_data_bus[10]), .A2(n8683), .B1(
        i_data_bus[746]), .B2(n8696), .ZN(n7735) );
  AOI22D1BWP30P140LVT U8310 ( .A1(i_data_bus[906]), .A2(n8686), .B1(
        i_data_bus[682]), .B2(n8689), .ZN(n7734) );
  ND4D1BWP30P140LVT U8311 ( .A1(n7737), .A2(n7736), .A3(n7735), .A4(n7734), 
        .ZN(n7744) );
  INVD1BWP30P140LVT U8312 ( .I(n8719), .ZN(n8647) );
  MOAI22D1BWP30P140LVT U8313 ( .A1(n8535), .A2(n8647), .B1(i_data_bus[202]), 
        .B2(n8713), .ZN(n7743) );
  AOI22D1BWP30P140LVT U8314 ( .A1(i_data_bus[170]), .A2(n8716), .B1(
        i_data_bus[426]), .B2(n8717), .ZN(n7741) );
  AOI22D1BWP30P140LVT U8315 ( .A1(i_data_bus[234]), .A2(n8687), .B1(
        i_data_bus[458]), .B2(n8626), .ZN(n7740) );
  AOI22D1BWP30P140LVT U8316 ( .A1(i_data_bus[554]), .A2(n8723), .B1(
        i_data_bus[522]), .B2(n8721), .ZN(n7739) );
  AOI22D1BWP30P140LVT U8317 ( .A1(i_data_bus[618]), .A2(n8720), .B1(
        i_data_bus[586]), .B2(n8722), .ZN(n7738) );
  ND4D1BWP30P140LVT U8318 ( .A1(n7741), .A2(n7740), .A3(n7739), .A4(n7738), 
        .ZN(n7742) );
  NR4D0BWP30P140LVT U8319 ( .A1(n7745), .A2(n7744), .A3(n7743), .A4(n7742), 
        .ZN(n7746) );
  ND4D4BWP30P140LVT U8320 ( .A1(n7749), .A2(n7748), .A3(n7747), .A4(n7746), 
        .ZN(o_data_bus[170]) );
  INR3D0BWP30P140LVT U8321 ( .A1(i_cmd[16]), .B1(n11699), .B2(n7759), .ZN(
        n9672) );
  NR3D0P7BWP30P140LVT U8322 ( .A1(n11735), .A2(n7750), .A3(n7756), .ZN(n9682)
         );
  AOI22D1BWP30P140LVT U8323 ( .A1(i_data_bus[95]), .A2(n9672), .B1(
        i_data_bus[927]), .B2(n9682), .ZN(n7791) );
  NR3D0P7BWP30P140LVT U8324 ( .A1(n11715), .A2(n7751), .A3(n7756), .ZN(n9678)
         );
  INR3D0BWP30P140LVT U8325 ( .A1(i_cmd[40]), .B1(n11023), .B2(n7760), .ZN(
        n9675) );
  AOI22D1BWP30P140LVT U8326 ( .A1(i_data_bus[991]), .A2(n9678), .B1(
        i_data_bus[191]), .B2(n9675), .ZN(n7790) );
  INVD1BWP30P140LVT U8327 ( .I(n7752), .ZN(n7753) );
  ND3D1BWP30P140LVT U8328 ( .A1(i_valid[8]), .A2(n7753), .A3(n7778), .ZN(n9181) );
  INVD1BWP30P140LVT U8329 ( .I(n9181), .ZN(n9694) );
  AN3D1BWP30P140LVT U8330 ( .A1(i_valid[21]), .A2(i_cmd[168]), .A3(n7776), .Z(
        n9705) );
  AOI22D1BWP30P140LVT U8331 ( .A1(i_data_bus[287]), .A2(n9694), .B1(
        i_data_bus[703]), .B2(n9705), .ZN(n7789) );
  NR3D0P7BWP30P140LVT U8332 ( .A1(n11717), .A2(n7754), .A3(n7756), .ZN(n9677)
         );
  INR3D0BWP30P140LVT U8333 ( .A1(i_cmd[8]), .B1(n11737), .B2(n7759), .ZN(n9670) );
  AOI22D1BWP30P140LVT U8334 ( .A1(i_data_bus[1023]), .A2(n9677), .B1(
        i_data_bus[63]), .B2(n9670), .ZN(n7764) );
  NR3D0P7BWP30P140LVT U8335 ( .A1(n11703), .A2(n7755), .A3(n7759), .ZN(n9676)
         );
  NR3D0P7BWP30P140LVT U8336 ( .A1(n11740), .A2(n7757), .A3(n7756), .ZN(n9669)
         );
  AOI22D1BWP30P140LVT U8337 ( .A1(i_data_bus[31]), .A2(n9676), .B1(
        i_data_bus[959]), .B2(n9669), .ZN(n7763) );
  INR3D0BWP30P140LVT U8338 ( .A1(i_cmd[48]), .B1(n11030), .B2(n7760), .ZN(
        n9679) );
  INVD1BWP30P140LVT U8339 ( .I(i_cmd[32]), .ZN(n7758) );
  NR3D0P7BWP30P140LVT U8340 ( .A1(n11721), .A2(n7758), .A3(n7760), .ZN(n9681)
         );
  AOI22D1BWP30P140LVT U8341 ( .A1(i_data_bus[223]), .A2(n9679), .B1(
        i_data_bus[159]), .B2(n9681), .ZN(n7762) );
  INR3D0BWP30P140LVT U8342 ( .A1(i_cmd[24]), .B1(n11726), .B2(n7759), .ZN(
        n9680) );
  INR3D0BWP30P140LVT U8343 ( .A1(i_cmd[56]), .B1(n11032), .B2(n7760), .ZN(
        n9671) );
  AOI22D1BWP30P140LVT U8344 ( .A1(i_data_bus[127]), .A2(n9680), .B1(
        i_data_bus[255]), .B2(n9671), .ZN(n7761) );
  ND4D1BWP30P140LVT U8345 ( .A1(n7764), .A2(n7763), .A3(n7762), .A4(n7761), 
        .ZN(n7787) );
  INVD1BWP30P140LVT U8346 ( .I(i_valid[14]), .ZN(n11706) );
  INR3D0BWP30P140LVT U8347 ( .A1(i_cmd[112]), .B1(n7774), .B2(n11706), .ZN(
        n9703) );
  INVD1BWP30P140LVT U8348 ( .I(n9703), .ZN(n9649) );
  NR3D0P7BWP30P140LVT U8349 ( .A1(n11754), .A2(n7765), .A3(n7779), .ZN(n9673)
         );
  MOAI22D1BWP30P140LVT U8350 ( .A1(n7766), .A2(n9649), .B1(i_data_bus[799]), 
        .B2(n9673), .ZN(n7786) );
  NR3D0P7BWP30P140LVT U8351 ( .A1(n11705), .A2(n7767), .A3(n7774), .ZN(n9708)
         );
  INR3D0BWP30P140LVT U8352 ( .A1(i_cmd[216]), .B1(n11749), .B2(n7779), .ZN(
        n9710) );
  AOI22D1BWP30P140LVT U8353 ( .A1(i_data_bus[415]), .A2(n9708), .B1(
        i_data_bus[895]), .B2(n9710), .ZN(n7773) );
  INVD1BWP30P140LVT U8354 ( .I(i_valid[13]), .ZN(n11698) );
  INR3D0BWP30P140LVT U8355 ( .A1(i_cmd[104]), .B1(n11698), .B2(n7774), .ZN(
        n9709) );
  AN3D1BWP30P140LVT U8356 ( .A1(i_valid[23]), .A2(i_cmd[184]), .A3(n7776), .Z(
        n9706) );
  AOI22D1BWP30P140LVT U8357 ( .A1(i_data_bus[447]), .A2(n9709), .B1(
        i_data_bus[767]), .B2(n9706), .ZN(n7772) );
  INR3D0BWP30P140LVT U8358 ( .A1(i_cmd[144]), .B1(n11733), .B2(n7769), .ZN(
        n9697) );
  INVD1BWP30P140LVT U8359 ( .I(i_cmd[128]), .ZN(n7768) );
  NR3D0P7BWP30P140LVT U8360 ( .A1(n11713), .A2(n7768), .A3(n7769), .ZN(n9698)
         );
  AOI22D1BWP30P140LVT U8361 ( .A1(i_data_bus[607]), .A2(n9697), .B1(
        i_data_bus[543]), .B2(n9698), .ZN(n7771) );
  INR3D0BWP30P140LVT U8362 ( .A1(i_cmd[136]), .B1(n11701), .B2(n7769), .ZN(
        n9695) );
  INR3D0BWP30P140LVT U8363 ( .A1(i_cmd[152]), .B1(n11697), .B2(n7769), .ZN(
        n9696) );
  AOI22D1BWP30P140LVT U8364 ( .A1(i_data_bus[575]), .A2(n9695), .B1(
        i_data_bus[639]), .B2(n9696), .ZN(n7770) );
  ND4D1BWP30P140LVT U8365 ( .A1(n7773), .A2(n7772), .A3(n7771), .A4(n7770), 
        .ZN(n7785) );
  INVD1BWP30P140LVT U8366 ( .I(i_valid[15]), .ZN(n11719) );
  INR3D0BWP30P140LVT U8367 ( .A1(i_cmd[120]), .B1(n7774), .B2(n11719), .ZN(
        n9656) );
  ND3D1BWP30P140LVT U8368 ( .A1(i_valid[10]), .A2(i_cmd[80]), .A3(n7778), .ZN(
        n9137) );
  INVD1BWP30P140LVT U8369 ( .I(n9137), .ZN(n9692) );
  AOI22D1BWP30P140LVT U8370 ( .A1(i_data_bus[511]), .A2(n9656), .B1(
        i_data_bus[351]), .B2(n9692), .ZN(n7783) );
  AN3D1BWP30P140LVT U8371 ( .A1(i_valid[22]), .A2(i_cmd[176]), .A3(n7776), .Z(
        n9704) );
  ND3D1BWP30P140LVT U8372 ( .A1(i_valid[11]), .A2(i_cmd[88]), .A3(n7778), .ZN(
        n9604) );
  INVD1BWP30P140LVT U8373 ( .I(n9604), .ZN(n9691) );
  AOI22D1BWP30P140LVT U8374 ( .A1(i_data_bus[735]), .A2(n9704), .B1(
        i_data_bus[383]), .B2(n9691), .ZN(n7782) );
  INVD1BWP30P140LVT U8375 ( .I(n7775), .ZN(n7777) );
  AN3D1BWP30P140LVT U8376 ( .A1(i_valid[20]), .A2(n7777), .A3(n7776), .Z(n9707) );
  INR3D0BWP30P140LVT U8377 ( .A1(i_cmd[208]), .B1(n11745), .B2(n7779), .ZN(
        n9693) );
  AOI22D1BWP30P140LVT U8378 ( .A1(i_data_bus[671]), .A2(n9707), .B1(
        i_data_bus[863]), .B2(n9693), .ZN(n7781) );
  ND3D1BWP30P140LVT U8379 ( .A1(i_valid[9]), .A2(i_cmd[72]), .A3(n7778), .ZN(
        n9687) );
  INVD1BWP30P140LVT U8380 ( .I(n9687), .ZN(n9655) );
  INR3D0BWP30P140LVT U8381 ( .A1(i_cmd[200]), .B1(n11751), .B2(n7779), .ZN(
        n9674) );
  AOI22D1BWP30P140LVT U8382 ( .A1(i_data_bus[319]), .A2(n9655), .B1(
        i_data_bus[831]), .B2(n9674), .ZN(n7780) );
  ND4D1BWP30P140LVT U8383 ( .A1(n7783), .A2(n7782), .A3(n7781), .A4(n7780), 
        .ZN(n7784) );
  NR4D0BWP30P140LVT U8384 ( .A1(n7787), .A2(n7786), .A3(n7785), .A4(n7784), 
        .ZN(n7788) );
  ND4D4BWP30P140LVT U8385 ( .A1(n7791), .A2(n7790), .A3(n7789), .A4(n7788), 
        .ZN(o_data_bus[31]) );
  AOI22D1BWP30P140LVT U8386 ( .A1(i_data_bus[62]), .A2(n9670), .B1(
        i_data_bus[190]), .B2(n9675), .ZN(n7811) );
  AOI22D1BWP30P140LVT U8387 ( .A1(i_data_bus[126]), .A2(n9680), .B1(
        i_data_bus[1022]), .B2(n9677), .ZN(n7810) );
  AOI22D1BWP30P140LVT U8388 ( .A1(i_data_bus[318]), .A2(n9655), .B1(
        i_data_bus[414]), .B2(n9708), .ZN(n7809) );
  AOI22D1BWP30P140LVT U8389 ( .A1(i_data_bus[446]), .A2(n9709), .B1(
        i_data_bus[702]), .B2(n9705), .ZN(n7807) );
  AOI22D1BWP30P140LVT U8390 ( .A1(i_data_bus[926]), .A2(n9682), .B1(
        i_data_bus[990]), .B2(n9678), .ZN(n7795) );
  AOI22D1BWP30P140LVT U8391 ( .A1(i_data_bus[30]), .A2(n9676), .B1(
        i_data_bus[94]), .B2(n9672), .ZN(n7794) );
  AOI22D1BWP30P140LVT U8392 ( .A1(i_data_bus[958]), .A2(n9669), .B1(
        i_data_bus[222]), .B2(n9679), .ZN(n7793) );
  AOI22D1BWP30P140LVT U8393 ( .A1(i_data_bus[254]), .A2(n9671), .B1(
        i_data_bus[158]), .B2(n9681), .ZN(n7792) );
  ND4D1BWP30P140LVT U8394 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), 
        .ZN(n7806) );
  AOI22D1BWP30P140LVT U8395 ( .A1(i_data_bus[350]), .A2(n9692), .B1(
        i_data_bus[766]), .B2(n9706), .ZN(n7799) );
  AOI22D1BWP30P140LVT U8396 ( .A1(i_data_bus[862]), .A2(n9693), .B1(
        i_data_bus[798]), .B2(n9673), .ZN(n7798) );
  AOI22D1BWP30P140LVT U8397 ( .A1(i_data_bus[574]), .A2(n9695), .B1(
        i_data_bus[606]), .B2(n9697), .ZN(n7797) );
  AOI22D1BWP30P140LVT U8398 ( .A1(i_data_bus[542]), .A2(n9698), .B1(
        i_data_bus[638]), .B2(n9696), .ZN(n7796) );
  ND4D1BWP30P140LVT U8399 ( .A1(n7799), .A2(n7798), .A3(n7797), .A4(n7796), 
        .ZN(n7805) );
  AOI22D1BWP30P140LVT U8400 ( .A1(i_data_bus[382]), .A2(n9691), .B1(
        i_data_bus[894]), .B2(n9710), .ZN(n7803) );
  AOI22D1BWP30P140LVT U8401 ( .A1(i_data_bus[670]), .A2(n9707), .B1(
        i_data_bus[510]), .B2(n9656), .ZN(n7802) );
  AOI22D1BWP30P140LVT U8402 ( .A1(i_data_bus[830]), .A2(n9674), .B1(
        i_data_bus[734]), .B2(n9704), .ZN(n7801) );
  AOI22D1BWP30P140LVT U8403 ( .A1(i_data_bus[286]), .A2(n9694), .B1(
        i_data_bus[478]), .B2(n9703), .ZN(n7800) );
  ND4D1BWP30P140LVT U8404 ( .A1(n7803), .A2(n7802), .A3(n7801), .A4(n7800), 
        .ZN(n7804) );
  INR4D0BWP30P140LVT U8405 ( .A1(n7807), .B1(n7806), .B2(n7805), .B3(n7804), 
        .ZN(n7808) );
  ND4D4BWP30P140LVT U8406 ( .A1(n7811), .A2(n7810), .A3(n7809), .A4(n7808), 
        .ZN(o_data_bus[30]) );
  AOI22D1BWP30P140LVT U8407 ( .A1(i_data_bus[976]), .A2(n9678), .B1(
        i_data_bus[16]), .B2(n9676), .ZN(n7831) );
  AOI22D1BWP30P140LVT U8408 ( .A1(i_data_bus[912]), .A2(n9682), .B1(
        i_data_bus[1008]), .B2(n9677), .ZN(n7830) );
  AOI22D1BWP30P140LVT U8409 ( .A1(i_data_bus[304]), .A2(n9655), .B1(
        i_data_bus[656]), .B2(n9707), .ZN(n7829) );
  AOI22D1BWP30P140LVT U8410 ( .A1(i_data_bus[144]), .A2(n9681), .B1(
        i_data_bus[176]), .B2(n9675), .ZN(n7815) );
  AOI22D1BWP30P140LVT U8411 ( .A1(i_data_bus[48]), .A2(n9670), .B1(
        i_data_bus[240]), .B2(n9671), .ZN(n7814) );
  AOI22D1BWP30P140LVT U8412 ( .A1(i_data_bus[80]), .A2(n9672), .B1(
        i_data_bus[112]), .B2(n9680), .ZN(n7813) );
  AOI22D1BWP30P140LVT U8413 ( .A1(i_data_bus[944]), .A2(n9669), .B1(
        i_data_bus[208]), .B2(n9679), .ZN(n7812) );
  ND4D1BWP30P140LVT U8414 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), 
        .ZN(n7827) );
  INVD1BWP30P140LVT U8415 ( .I(n9708), .ZN(n9626) );
  MOAI22D1BWP30P140LVT U8416 ( .A1(n7899), .A2(n9626), .B1(i_data_bus[880]), 
        .B2(n9710), .ZN(n7826) );
  AOI22D1BWP30P140LVT U8417 ( .A1(i_data_bus[464]), .A2(n9703), .B1(
        i_data_bus[688]), .B2(n9705), .ZN(n7819) );
  AOI22D1BWP30P140LVT U8418 ( .A1(i_data_bus[336]), .A2(n9692), .B1(
        i_data_bus[720]), .B2(n9704), .ZN(n7818) );
  AOI22D1BWP30P140LVT U8419 ( .A1(i_data_bus[560]), .A2(n9695), .B1(
        i_data_bus[624]), .B2(n9696), .ZN(n7817) );
  AOI22D1BWP30P140LVT U8420 ( .A1(i_data_bus[528]), .A2(n9698), .B1(
        i_data_bus[592]), .B2(n9697), .ZN(n7816) );
  ND4D1BWP30P140LVT U8421 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), 
        .ZN(n7825) );
  AOI22D1BWP30P140LVT U8422 ( .A1(i_data_bus[784]), .A2(n9673), .B1(
        i_data_bus[272]), .B2(n9694), .ZN(n7823) );
  AOI22D1BWP30P140LVT U8423 ( .A1(i_data_bus[816]), .A2(n9674), .B1(
        i_data_bus[848]), .B2(n9693), .ZN(n7822) );
  AOI22D1BWP30P140LVT U8424 ( .A1(i_data_bus[496]), .A2(n9656), .B1(
        i_data_bus[368]), .B2(n9691), .ZN(n7821) );
  AOI22D1BWP30P140LVT U8425 ( .A1(i_data_bus[432]), .A2(n9709), .B1(
        i_data_bus[752]), .B2(n9706), .ZN(n7820) );
  ND4D1BWP30P140LVT U8426 ( .A1(n7823), .A2(n7822), .A3(n7821), .A4(n7820), 
        .ZN(n7824) );
  NR4D0BWP30P140LVT U8427 ( .A1(n7827), .A2(n7826), .A3(n7825), .A4(n7824), 
        .ZN(n7828) );
  ND4D4BWP30P140LVT U8428 ( .A1(n7831), .A2(n7830), .A3(n7829), .A4(n7828), 
        .ZN(o_data_bus[16]) );
  AOI22D1BWP30P140LVT U8429 ( .A1(i_data_bus[765]), .A2(n9546), .B1(
        i_data_bus[797]), .B2(n9547), .ZN(n7852) );
  AOI22D1BWP30P140LVT U8430 ( .A1(i_data_bus[669]), .A2(n9558), .B1(
        i_data_bus[829]), .B2(n9552), .ZN(n7851) );
  AOI22D1BWP30P140LVT U8431 ( .A1(i_data_bus[349]), .A2(n9570), .B1(
        i_data_bus[285]), .B2(n9586), .ZN(n7850) );
  AOI22D1BWP30P140LVT U8432 ( .A1(i_data_bus[29]), .A2(n9553), .B1(
        i_data_bus[125]), .B2(n9555), .ZN(n7835) );
  AOI22D1BWP30P140LVT U8433 ( .A1(i_data_bus[61]), .A2(n9548), .B1(
        i_data_bus[893]), .B2(n9556), .ZN(n7834) );
  AOI22D1BWP30P140LVT U8434 ( .A1(i_data_bus[93]), .A2(n9549), .B1(
        i_data_bus[861]), .B2(n9557), .ZN(n7833) );
  AOI22D1BWP30P140LVT U8435 ( .A1(i_data_bus[701]), .A2(n9559), .B1(
        i_data_bus[733]), .B2(n9554), .ZN(n7832) );
  ND4D1BWP30P140LVT U8436 ( .A1(n7835), .A2(n7834), .A3(n7833), .A4(n7832), 
        .ZN(n7848) );
  MOAI22D1BWP30P140LVT U8437 ( .A1(n7836), .A2(n9375), .B1(i_data_bus[157]), 
        .B2(n9533), .ZN(n7847) );
  AOI22D1BWP30P140LVT U8438 ( .A1(i_data_bus[925]), .A2(n9581), .B1(
        i_data_bus[957]), .B2(n9587), .ZN(n7840) );
  AOI22D1BWP30P140LVT U8439 ( .A1(i_data_bus[989]), .A2(n9551), .B1(
        i_data_bus[413]), .B2(n9585), .ZN(n7839) );
  AOI22D1BWP30P140LVT U8440 ( .A1(i_data_bus[573]), .A2(n9575), .B1(
        i_data_bus[541]), .B2(n9573), .ZN(n7838) );
  AOI22D1BWP30P140LVT U8441 ( .A1(i_data_bus[637]), .A2(n9574), .B1(
        i_data_bus[605]), .B2(n9572), .ZN(n7837) );
  ND4D1BWP30P140LVT U8442 ( .A1(n7840), .A2(n7839), .A3(n7838), .A4(n7837), 
        .ZN(n7846) );
  AOI22D1BWP30P140LVT U8443 ( .A1(i_data_bus[1021]), .A2(n9571), .B1(
        i_data_bus[221]), .B2(n9550), .ZN(n7844) );
  AOI22D1BWP30P140LVT U8444 ( .A1(i_data_bus[445]), .A2(n9532), .B1(
        i_data_bus[253]), .B2(n9568), .ZN(n7843) );
  AOI22D1BWP30P140LVT U8445 ( .A1(i_data_bus[317]), .A2(n9584), .B1(
        i_data_bus[509]), .B2(n9580), .ZN(n7842) );
  AOI22D1BWP30P140LVT U8446 ( .A1(i_data_bus[189]), .A2(n9583), .B1(
        i_data_bus[477]), .B2(n9582), .ZN(n7841) );
  ND4D1BWP30P140LVT U8447 ( .A1(n7844), .A2(n7843), .A3(n7842), .A4(n7841), 
        .ZN(n7845) );
  NR4D0BWP30P140LVT U8448 ( .A1(n7848), .A2(n7847), .A3(n7846), .A4(n7845), 
        .ZN(n7849) );
  ND4D4BWP30P140LVT U8449 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), 
        .ZN(o_data_bus[253]) );
  AOI22D1BWP30P140LVT U8450 ( .A1(i_data_bus[120]), .A2(n9555), .B1(
        i_data_bus[696]), .B2(n9559), .ZN(n7873) );
  AOI22D1BWP30P140LVT U8451 ( .A1(i_data_bus[824]), .A2(n9552), .B1(
        i_data_bus[760]), .B2(n9546), .ZN(n7872) );
  AOI22D1BWP30P140LVT U8452 ( .A1(i_data_bus[344]), .A2(n9570), .B1(
        i_data_bus[376]), .B2(n9569), .ZN(n7871) );
  AOI22D1BWP30P140LVT U8453 ( .A1(i_data_bus[56]), .A2(n9548), .B1(
        i_data_bus[664]), .B2(n9558), .ZN(n7856) );
  AOI22D1BWP30P140LVT U8454 ( .A1(i_data_bus[856]), .A2(n9557), .B1(
        i_data_bus[728]), .B2(n9554), .ZN(n7855) );
  AOI22D1BWP30P140LVT U8455 ( .A1(i_data_bus[24]), .A2(n9553), .B1(
        i_data_bus[792]), .B2(n9547), .ZN(n7854) );
  AOI22D1BWP30P140LVT U8456 ( .A1(i_data_bus[88]), .A2(n9549), .B1(
        i_data_bus[888]), .B2(n9556), .ZN(n7853) );
  ND4D1BWP30P140LVT U8457 ( .A1(n7856), .A2(n7855), .A3(n7854), .A4(n7853), 
        .ZN(n7869) );
  INVD1BWP30P140LVT U8458 ( .I(n9586), .ZN(n8390) );
  MOAI22D1BWP30P140LVT U8459 ( .A1(n7857), .A2(n8390), .B1(i_data_bus[152]), 
        .B2(n9533), .ZN(n7868) );
  AOI22D1BWP30P140LVT U8460 ( .A1(i_data_bus[1016]), .A2(n9571), .B1(
        i_data_bus[472]), .B2(n9582), .ZN(n7861) );
  AOI22D1BWP30P140LVT U8461 ( .A1(i_data_bus[248]), .A2(n9568), .B1(
        i_data_bus[312]), .B2(n9584), .ZN(n7860) );
  AOI22D1BWP30P140LVT U8462 ( .A1(i_data_bus[632]), .A2(n9574), .B1(
        i_data_bus[568]), .B2(n9575), .ZN(n7859) );
  AOI22D1BWP30P140LVT U8463 ( .A1(i_data_bus[600]), .A2(n9572), .B1(
        i_data_bus[536]), .B2(n9573), .ZN(n7858) );
  ND4D1BWP30P140LVT U8464 ( .A1(n7861), .A2(n7860), .A3(n7859), .A4(n7858), 
        .ZN(n7867) );
  AOI22D1BWP30P140LVT U8465 ( .A1(i_data_bus[216]), .A2(n9550), .B1(
        i_data_bus[504]), .B2(n9580), .ZN(n7865) );
  AOI22D1BWP30P140LVT U8466 ( .A1(i_data_bus[984]), .A2(n9551), .B1(
        i_data_bus[952]), .B2(n9587), .ZN(n7864) );
  AOI22D1BWP30P140LVT U8467 ( .A1(i_data_bus[920]), .A2(n9581), .B1(
        i_data_bus[184]), .B2(n9583), .ZN(n7863) );
  AOI22D1BWP30P140LVT U8468 ( .A1(i_data_bus[408]), .A2(n9585), .B1(
        i_data_bus[440]), .B2(n9532), .ZN(n7862) );
  ND4D1BWP30P140LVT U8469 ( .A1(n7865), .A2(n7864), .A3(n7863), .A4(n7862), 
        .ZN(n7866) );
  NR4D0BWP30P140LVT U8470 ( .A1(n7869), .A2(n7868), .A3(n7867), .A4(n7866), 
        .ZN(n7870) );
  ND4D4BWP30P140LVT U8471 ( .A1(n7873), .A2(n7872), .A3(n7871), .A4(n7870), 
        .ZN(o_data_bus[248]) );
  AOI22D1BWP30P140LVT U8472 ( .A1(i_data_bus[115]), .A2(n9555), .B1(
        i_data_bus[819]), .B2(n9552), .ZN(n7894) );
  AOI22D1BWP30P140LVT U8473 ( .A1(i_data_bus[691]), .A2(n9559), .B1(
        i_data_bus[723]), .B2(n9554), .ZN(n7893) );
  AOI22D1BWP30P140LVT U8474 ( .A1(i_data_bus[307]), .A2(n9584), .B1(
        i_data_bus[275]), .B2(n9586), .ZN(n7892) );
  AOI22D1BWP30P140LVT U8475 ( .A1(i_data_bus[83]), .A2(n9549), .B1(
        i_data_bus[659]), .B2(n9558), .ZN(n7877) );
  AOI22D1BWP30P140LVT U8476 ( .A1(i_data_bus[19]), .A2(n9553), .B1(
        i_data_bus[851]), .B2(n9557), .ZN(n7876) );
  AOI22D1BWP30P140LVT U8477 ( .A1(i_data_bus[755]), .A2(n9546), .B1(
        i_data_bus[883]), .B2(n9556), .ZN(n7875) );
  AOI22D1BWP30P140LVT U8478 ( .A1(i_data_bus[51]), .A2(n9548), .B1(
        i_data_bus[787]), .B2(n9547), .ZN(n7874) );
  ND4D1BWP30P140LVT U8479 ( .A1(n7877), .A2(n7876), .A3(n7875), .A4(n7874), 
        .ZN(n7890) );
  MOAI22D1BWP30P140LVT U8480 ( .A1(n7878), .A2(n9397), .B1(i_data_bus[947]), 
        .B2(n9587), .ZN(n7889) );
  AOI22D1BWP30P140LVT U8481 ( .A1(i_data_bus[979]), .A2(n9551), .B1(
        i_data_bus[211]), .B2(n9550), .ZN(n7882) );
  AOI22D1BWP30P140LVT U8482 ( .A1(i_data_bus[1011]), .A2(n9571), .B1(
        i_data_bus[403]), .B2(n9585), .ZN(n7881) );
  AOI22D1BWP30P140LVT U8483 ( .A1(i_data_bus[531]), .A2(n9573), .B1(
        i_data_bus[595]), .B2(n9572), .ZN(n7880) );
  AOI22D1BWP30P140LVT U8484 ( .A1(i_data_bus[563]), .A2(n9575), .B1(
        i_data_bus[627]), .B2(n9574), .ZN(n7879) );
  ND4D1BWP30P140LVT U8485 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), 
        .ZN(n7888) );
  AOI22D1BWP30P140LVT U8486 ( .A1(i_data_bus[339]), .A2(n9570), .B1(
        i_data_bus[435]), .B2(n9532), .ZN(n7886) );
  AOI22D1BWP30P140LVT U8487 ( .A1(i_data_bus[915]), .A2(n9581), .B1(
        i_data_bus[467]), .B2(n9582), .ZN(n7885) );
  AOI22D1BWP30P140LVT U8488 ( .A1(i_data_bus[371]), .A2(n9569), .B1(
        i_data_bus[243]), .B2(n9568), .ZN(n7884) );
  AOI22D1BWP30P140LVT U8489 ( .A1(i_data_bus[179]), .A2(n9583), .B1(
        i_data_bus[147]), .B2(n9533), .ZN(n7883) );
  ND4D1BWP30P140LVT U8490 ( .A1(n7886), .A2(n7885), .A3(n7884), .A4(n7883), 
        .ZN(n7887) );
  NR4D0BWP30P140LVT U8491 ( .A1(n7890), .A2(n7889), .A3(n7888), .A4(n7887), 
        .ZN(n7891) );
  ND4D4BWP30P140LVT U8492 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), 
        .ZN(o_data_bus[243]) );
  AOI22D1BWP30P140LVT U8493 ( .A1(i_data_bus[880]), .A2(n9556), .B1(
        i_data_bus[656]), .B2(n9558), .ZN(n7915) );
  AOI22D1BWP30P140LVT U8494 ( .A1(i_data_bus[80]), .A2(n9549), .B1(
        i_data_bus[720]), .B2(n9554), .ZN(n7914) );
  AOI22D1BWP30P140LVT U8495 ( .A1(i_data_bus[304]), .A2(n9584), .B1(
        i_data_bus[272]), .B2(n9586), .ZN(n7913) );
  AOI22D1BWP30P140LVT U8496 ( .A1(i_data_bus[784]), .A2(n9547), .B1(
        i_data_bus[848]), .B2(n9557), .ZN(n7898) );
  AOI22D1BWP30P140LVT U8497 ( .A1(i_data_bus[112]), .A2(n9555), .B1(
        i_data_bus[688]), .B2(n9559), .ZN(n7897) );
  AOI22D1BWP30P140LVT U8498 ( .A1(i_data_bus[48]), .A2(n9548), .B1(
        i_data_bus[752]), .B2(n9546), .ZN(n7896) );
  AOI22D1BWP30P140LVT U8499 ( .A1(i_data_bus[16]), .A2(n9553), .B1(
        i_data_bus[816]), .B2(n9552), .ZN(n7895) );
  ND4D1BWP30P140LVT U8500 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), 
        .ZN(n7911) );
  MOAI22D1BWP30P140LVT U8501 ( .A1(n7899), .A2(n9245), .B1(i_data_bus[208]), 
        .B2(n9550), .ZN(n7910) );
  AOI22D1BWP30P140LVT U8502 ( .A1(i_data_bus[1008]), .A2(n9571), .B1(
        i_data_bus[432]), .B2(n9532), .ZN(n7903) );
  AOI22D1BWP30P140LVT U8503 ( .A1(i_data_bus[944]), .A2(n9587), .B1(
        i_data_bus[144]), .B2(n9533), .ZN(n7902) );
  AOI22D1BWP30P140LVT U8504 ( .A1(i_data_bus[560]), .A2(n9575), .B1(
        i_data_bus[592]), .B2(n9572), .ZN(n7901) );
  AOI22D1BWP30P140LVT U8505 ( .A1(i_data_bus[528]), .A2(n9573), .B1(
        i_data_bus[624]), .B2(n9574), .ZN(n7900) );
  ND4D1BWP30P140LVT U8506 ( .A1(n7903), .A2(n7902), .A3(n7901), .A4(n7900), 
        .ZN(n7909) );
  AOI22D1BWP30P140LVT U8507 ( .A1(i_data_bus[336]), .A2(n9570), .B1(
        i_data_bus[496]), .B2(n9580), .ZN(n7907) );
  AOI22D1BWP30P140LVT U8508 ( .A1(i_data_bus[976]), .A2(n9551), .B1(
        i_data_bus[464]), .B2(n9582), .ZN(n7906) );
  AOI22D1BWP30P140LVT U8509 ( .A1(i_data_bus[912]), .A2(n9581), .B1(
        i_data_bus[240]), .B2(n9568), .ZN(n7905) );
  AOI22D1BWP30P140LVT U8510 ( .A1(i_data_bus[176]), .A2(n9583), .B1(
        i_data_bus[368]), .B2(n9569), .ZN(n7904) );
  ND4D1BWP30P140LVT U8511 ( .A1(n7907), .A2(n7906), .A3(n7905), .A4(n7904), 
        .ZN(n7908) );
  NR4D0BWP30P140LVT U8512 ( .A1(n7911), .A2(n7910), .A3(n7909), .A4(n7908), 
        .ZN(n7912) );
  ND4D4BWP30P140LVT U8513 ( .A1(n7915), .A2(n7914), .A3(n7913), .A4(n7912), 
        .ZN(o_data_bus[240]) );
  AOI22D1BWP30P140LVT U8514 ( .A1(i_data_bus[111]), .A2(n9555), .B1(
        i_data_bus[687]), .B2(n9559), .ZN(n7936) );
  AOI22D1BWP30P140LVT U8515 ( .A1(i_data_bus[47]), .A2(n9548), .B1(
        i_data_bus[783]), .B2(n9547), .ZN(n7935) );
  AOI22D1BWP30P140LVT U8516 ( .A1(i_data_bus[431]), .A2(n9532), .B1(
        i_data_bus[463]), .B2(n9582), .ZN(n7934) );
  AOI22D1BWP30P140LVT U8517 ( .A1(i_data_bus[719]), .A2(n9554), .B1(
        i_data_bus[655]), .B2(n9558), .ZN(n7919) );
  AOI22D1BWP30P140LVT U8518 ( .A1(i_data_bus[15]), .A2(n9553), .B1(
        i_data_bus[751]), .B2(n9546), .ZN(n7918) );
  AOI22D1BWP30P140LVT U8519 ( .A1(i_data_bus[879]), .A2(n9556), .B1(
        i_data_bus[815]), .B2(n9552), .ZN(n7917) );
  AOI22D1BWP30P140LVT U8520 ( .A1(i_data_bus[79]), .A2(n9549), .B1(
        i_data_bus[847]), .B2(n9557), .ZN(n7916) );
  ND4D1BWP30P140LVT U8521 ( .A1(n7919), .A2(n7918), .A3(n7917), .A4(n7916), 
        .ZN(n7932) );
  MOAI22D1BWP30P140LVT U8522 ( .A1(n7920), .A2(n9375), .B1(i_data_bus[335]), 
        .B2(n9570), .ZN(n7931) );
  AOI22D1BWP30P140LVT U8523 ( .A1(i_data_bus[911]), .A2(n9581), .B1(
        i_data_bus[943]), .B2(n9587), .ZN(n7924) );
  AOI22D1BWP30P140LVT U8524 ( .A1(i_data_bus[1007]), .A2(n9571), .B1(
        i_data_bus[239]), .B2(n9568), .ZN(n7923) );
  AOI22D1BWP30P140LVT U8525 ( .A1(i_data_bus[591]), .A2(n9572), .B1(
        i_data_bus[527]), .B2(n9573), .ZN(n7922) );
  AOI22D1BWP30P140LVT U8526 ( .A1(i_data_bus[559]), .A2(n9575), .B1(
        i_data_bus[623]), .B2(n9574), .ZN(n7921) );
  ND4D1BWP30P140LVT U8527 ( .A1(n7924), .A2(n7923), .A3(n7922), .A4(n7921), 
        .ZN(n7930) );
  AOI22D1BWP30P140LVT U8528 ( .A1(i_data_bus[175]), .A2(n9583), .B1(
        i_data_bus[143]), .B2(n9533), .ZN(n7928) );
  AOI22D1BWP30P140LVT U8529 ( .A1(i_data_bus[207]), .A2(n9550), .B1(
        i_data_bus[399]), .B2(n9585), .ZN(n7927) );
  AOI22D1BWP30P140LVT U8530 ( .A1(i_data_bus[975]), .A2(n9551), .B1(
        i_data_bus[271]), .B2(n9586), .ZN(n7926) );
  AOI22D1BWP30P140LVT U8531 ( .A1(i_data_bus[495]), .A2(n9580), .B1(
        i_data_bus[303]), .B2(n9584), .ZN(n7925) );
  ND4D1BWP30P140LVT U8532 ( .A1(n7928), .A2(n7927), .A3(n7926), .A4(n7925), 
        .ZN(n7929) );
  NR4D0BWP30P140LVT U8533 ( .A1(n7932), .A2(n7931), .A3(n7930), .A4(n7929), 
        .ZN(n7933) );
  ND4D4BWP30P140LVT U8534 ( .A1(n7936), .A2(n7935), .A3(n7934), .A4(n7933), 
        .ZN(o_data_bus[239]) );
  AOI22D1BWP30P140LVT U8535 ( .A1(i_data_bus[12]), .A2(n9553), .B1(
        i_data_bus[108]), .B2(n9555), .ZN(n7956) );
  AOI22D1BWP30P140LVT U8536 ( .A1(i_data_bus[44]), .A2(n9548), .B1(
        i_data_bus[684]), .B2(n9559), .ZN(n7955) );
  AOI22D1BWP30P140LVT U8537 ( .A1(i_data_bus[460]), .A2(n9582), .B1(
        i_data_bus[492]), .B2(n9580), .ZN(n7954) );
  AOI22D1BWP30P140LVT U8538 ( .A1(i_data_bus[748]), .A2(n9546), .B1(
        i_data_bus[844]), .B2(n9557), .ZN(n7940) );
  AOI22D1BWP30P140LVT U8539 ( .A1(i_data_bus[780]), .A2(n9547), .B1(
        i_data_bus[876]), .B2(n9556), .ZN(n7939) );
  AOI22D1BWP30P140LVT U8540 ( .A1(i_data_bus[812]), .A2(n9552), .B1(
        i_data_bus[652]), .B2(n9558), .ZN(n7938) );
  AOI22D1BWP30P140LVT U8541 ( .A1(i_data_bus[76]), .A2(n9549), .B1(
        i_data_bus[716]), .B2(n9554), .ZN(n7937) );
  ND4D1BWP30P140LVT U8542 ( .A1(n7940), .A2(n7939), .A3(n7938), .A4(n7937), 
        .ZN(n7952) );
  INVD1BWP30P140LVT U8543 ( .I(i_data_bus[172]), .ZN(n8272) );
  MOAI22D1BWP30P140LVT U8544 ( .A1(n8272), .A2(n9419), .B1(i_data_bus[236]), 
        .B2(n9568), .ZN(n7951) );
  AOI22D1BWP30P140LVT U8545 ( .A1(i_data_bus[1004]), .A2(n9571), .B1(
        i_data_bus[300]), .B2(n9584), .ZN(n7944) );
  AOI22D1BWP30P140LVT U8546 ( .A1(i_data_bus[908]), .A2(n9581), .B1(
        i_data_bus[972]), .B2(n9551), .ZN(n7943) );
  AOI22D1BWP30P140LVT U8547 ( .A1(i_data_bus[524]), .A2(n9573), .B1(
        i_data_bus[588]), .B2(n9572), .ZN(n7942) );
  AOI22D1BWP30P140LVT U8548 ( .A1(i_data_bus[620]), .A2(n9574), .B1(
        i_data_bus[556]), .B2(n9575), .ZN(n7941) );
  ND4D1BWP30P140LVT U8549 ( .A1(n7944), .A2(n7943), .A3(n7942), .A4(n7941), 
        .ZN(n7950) );
  AOI22D1BWP30P140LVT U8550 ( .A1(i_data_bus[940]), .A2(n9587), .B1(
        i_data_bus[140]), .B2(n9533), .ZN(n7948) );
  AOI22D1BWP30P140LVT U8551 ( .A1(i_data_bus[268]), .A2(n9586), .B1(
        i_data_bus[204]), .B2(n9550), .ZN(n7947) );
  AOI22D1BWP30P140LVT U8552 ( .A1(i_data_bus[364]), .A2(n9569), .B1(
        i_data_bus[396]), .B2(n9585), .ZN(n7946) );
  AOI22D1BWP30P140LVT U8553 ( .A1(i_data_bus[428]), .A2(n9532), .B1(
        i_data_bus[332]), .B2(n9570), .ZN(n7945) );
  ND4D1BWP30P140LVT U8554 ( .A1(n7948), .A2(n7947), .A3(n7946), .A4(n7945), 
        .ZN(n7949) );
  NR4D0BWP30P140LVT U8555 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), 
        .ZN(n7953) );
  ND4D4BWP30P140LVT U8556 ( .A1(n7956), .A2(n7955), .A3(n7954), .A4(n7953), 
        .ZN(o_data_bus[236]) );
  AOI22D1BWP30P140LVT U8557 ( .A1(i_data_bus[991]), .A2(n8708), .B1(
        i_data_bus[703]), .B2(n8689), .ZN(n7976) );
  AOI22D1BWP30P140LVT U8558 ( .A1(i_data_bus[671]), .A2(n8693), .B1(
        i_data_bus[767]), .B2(n8696), .ZN(n7975) );
  AOI22D1BWP30P140LVT U8559 ( .A1(i_data_bus[447]), .A2(n8717), .B1(
        i_data_bus[159]), .B2(n8688), .ZN(n7974) );
  AOI22D1BWP30P140LVT U8560 ( .A1(i_data_bus[63]), .A2(n8684), .B1(
        i_data_bus[831]), .B2(n8695), .ZN(n7960) );
  AOI22D1BWP30P140LVT U8561 ( .A1(i_data_bus[799]), .A2(n8707), .B1(
        i_data_bus[351]), .B2(n8685), .ZN(n7959) );
  AOI22D1BWP30P140LVT U8562 ( .A1(i_data_bus[927]), .A2(n8686), .B1(
        i_data_bus[127]), .B2(n8692), .ZN(n7958) );
  AOI22D1BWP30P140LVT U8563 ( .A1(i_data_bus[959]), .A2(n8704), .B1(
        i_data_bus[735]), .B2(n8703), .ZN(n7957) );
  ND4D1BWP30P140LVT U8564 ( .A1(n7960), .A2(n7959), .A3(n7958), .A4(n7957), 
        .ZN(n7972) );
  AOI22D1BWP30P140LVT U8565 ( .A1(i_data_bus[95]), .A2(n8694), .B1(
        i_data_bus[863]), .B2(n8690), .ZN(n7964) );
  AOI22D1BWP30P140LVT U8566 ( .A1(i_data_bus[31]), .A2(n8683), .B1(
        i_data_bus[287]), .B2(n8691), .ZN(n7963) );
  AOI22D1BWP30P140LVT U8567 ( .A1(i_data_bus[1023]), .A2(n8702), .B1(
        i_data_bus[895]), .B2(n8706), .ZN(n7962) );
  AOI22D1BWP30P140LVT U8568 ( .A1(i_data_bus[319]), .A2(n8705), .B1(
        i_data_bus[383]), .B2(n8701), .ZN(n7961) );
  ND4D1BWP30P140LVT U8569 ( .A1(n7964), .A2(n7963), .A3(n7962), .A4(n7961), 
        .ZN(n7971) );
  INVD1BWP30P140LVT U8570 ( .I(i_data_bus[191]), .ZN(n9203) );
  MOAI22D1BWP30P140LVT U8571 ( .A1(n9203), .A2(n8602), .B1(i_data_bus[223]), 
        .B2(n8713), .ZN(n7970) );
  AOI22D1BWP30P140LVT U8572 ( .A1(i_data_bus[511]), .A2(n8718), .B1(
        i_data_bus[255]), .B2(n8687), .ZN(n7968) );
  AOI22D1BWP30P140LVT U8573 ( .A1(i_data_bus[415]), .A2(n8719), .B1(
        i_data_bus[479]), .B2(n8626), .ZN(n7967) );
  AOI22D1BWP30P140LVT U8574 ( .A1(i_data_bus[575]), .A2(n8723), .B1(
        i_data_bus[543]), .B2(n8721), .ZN(n7966) );
  AOI22D1BWP30P140LVT U8575 ( .A1(i_data_bus[607]), .A2(n8722), .B1(
        i_data_bus[639]), .B2(n8720), .ZN(n7965) );
  ND4D1BWP30P140LVT U8576 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), 
        .ZN(n7969) );
  NR4D0BWP30P140LVT U8577 ( .A1(n7972), .A2(n7971), .A3(n7970), .A4(n7969), 
        .ZN(n7973) );
  ND4D4BWP30P140LVT U8578 ( .A1(n7976), .A2(n7975), .A3(n7974), .A4(n7973), 
        .ZN(o_data_bus[191]) );
  AOI22D1BWP30P140LVT U8579 ( .A1(i_data_bus[926]), .A2(n8686), .B1(
        i_data_bus[62]), .B2(n8684), .ZN(n7996) );
  AOI22D1BWP30P140LVT U8580 ( .A1(i_data_bus[30]), .A2(n8683), .B1(
        i_data_bus[734]), .B2(n8703), .ZN(n7995) );
  AOI22D1BWP30P140LVT U8581 ( .A1(i_data_bus[222]), .A2(n8713), .B1(
        i_data_bus[158]), .B2(n8688), .ZN(n7994) );
  AOI22D1BWP30P140LVT U8582 ( .A1(i_data_bus[798]), .A2(n8707), .B1(
        i_data_bus[766]), .B2(n8696), .ZN(n7980) );
  AOI22D1BWP30P140LVT U8583 ( .A1(i_data_bus[990]), .A2(n8708), .B1(
        i_data_bus[702]), .B2(n8689), .ZN(n7979) );
  AOI22D1BWP30P140LVT U8584 ( .A1(i_data_bus[670]), .A2(n8693), .B1(
        i_data_bus[894]), .B2(n8706), .ZN(n7978) );
  AOI22D1BWP30P140LVT U8585 ( .A1(i_data_bus[862]), .A2(n8690), .B1(
        i_data_bus[382]), .B2(n8701), .ZN(n7977) );
  ND4D1BWP30P140LVT U8586 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), 
        .ZN(n7992) );
  AOI22D1BWP30P140LVT U8587 ( .A1(i_data_bus[958]), .A2(n8704), .B1(
        i_data_bus[830]), .B2(n8695), .ZN(n7984) );
  AOI22D1BWP30P140LVT U8588 ( .A1(i_data_bus[126]), .A2(n8692), .B1(
        i_data_bus[318]), .B2(n8705), .ZN(n7983) );
  AOI22D1BWP30P140LVT U8589 ( .A1(i_data_bus[1022]), .A2(n8702), .B1(
        i_data_bus[286]), .B2(n8691), .ZN(n7982) );
  AOI22D1BWP30P140LVT U8590 ( .A1(i_data_bus[94]), .A2(n8694), .B1(
        i_data_bus[350]), .B2(n8685), .ZN(n7981) );
  ND4D1BWP30P140LVT U8591 ( .A1(n7984), .A2(n7983), .A3(n7982), .A4(n7981), 
        .ZN(n7991) );
  MOAI22D1BWP30P140LVT U8592 ( .A1(n9224), .A2(n8647), .B1(i_data_bus[510]), 
        .B2(n8718), .ZN(n7990) );
  AOI22D1BWP30P140LVT U8593 ( .A1(i_data_bus[446]), .A2(n8717), .B1(
        i_data_bus[254]), .B2(n8687), .ZN(n7988) );
  AOI22D1BWP30P140LVT U8594 ( .A1(i_data_bus[190]), .A2(n8716), .B1(
        i_data_bus[478]), .B2(n8626), .ZN(n7987) );
  AOI22D1BWP30P140LVT U8595 ( .A1(i_data_bus[606]), .A2(n8722), .B1(
        i_data_bus[638]), .B2(n8720), .ZN(n7986) );
  AOI22D1BWP30P140LVT U8596 ( .A1(i_data_bus[542]), .A2(n8721), .B1(
        i_data_bus[574]), .B2(n8723), .ZN(n7985) );
  ND4D1BWP30P140LVT U8597 ( .A1(n7988), .A2(n7987), .A3(n7986), .A4(n7985), 
        .ZN(n7989) );
  NR4D0BWP30P140LVT U8598 ( .A1(n7992), .A2(n7991), .A3(n7990), .A4(n7989), 
        .ZN(n7993) );
  ND4D4BWP30P140LVT U8599 ( .A1(n7996), .A2(n7995), .A3(n7994), .A4(n7993), 
        .ZN(o_data_bus[190]) );
  AOI22D1BWP30P140LVT U8600 ( .A1(i_data_bus[60]), .A2(n8684), .B1(
        i_data_bus[860]), .B2(n8690), .ZN(n8017) );
  AOI22D1BWP30P140LVT U8601 ( .A1(i_data_bus[924]), .A2(n8686), .B1(
        i_data_bus[348]), .B2(n8685), .ZN(n8016) );
  AOI22D1BWP30P140LVT U8602 ( .A1(i_data_bus[252]), .A2(n8687), .B1(
        i_data_bus[188]), .B2(n8716), .ZN(n8015) );
  AOI22D1BWP30P140LVT U8603 ( .A1(i_data_bus[92]), .A2(n8694), .B1(
        i_data_bus[700]), .B2(n8689), .ZN(n8000) );
  AOI22D1BWP30P140LVT U8604 ( .A1(i_data_bus[988]), .A2(n8708), .B1(
        i_data_bus[668]), .B2(n8693), .ZN(n7999) );
  AOI22D1BWP30P140LVT U8605 ( .A1(i_data_bus[1020]), .A2(n8702), .B1(
        i_data_bus[892]), .B2(n8706), .ZN(n7998) );
  AOI22D1BWP30P140LVT U8606 ( .A1(i_data_bus[956]), .A2(n8704), .B1(
        i_data_bus[732]), .B2(n8703), .ZN(n7997) );
  ND4D1BWP30P140LVT U8607 ( .A1(n8000), .A2(n7999), .A3(n7998), .A4(n7997), 
        .ZN(n8013) );
  AOI22D1BWP30P140LVT U8608 ( .A1(i_data_bus[28]), .A2(n8683), .B1(
        i_data_bus[828]), .B2(n8695), .ZN(n8004) );
  AOI22D1BWP30P140LVT U8609 ( .A1(i_data_bus[124]), .A2(n8692), .B1(
        i_data_bus[764]), .B2(n8696), .ZN(n8003) );
  AOI22D1BWP30P140LVT U8610 ( .A1(i_data_bus[284]), .A2(n8691), .B1(
        i_data_bus[316]), .B2(n8705), .ZN(n8002) );
  AOI22D1BWP30P140LVT U8611 ( .A1(i_data_bus[380]), .A2(n8701), .B1(
        i_data_bus[796]), .B2(n8707), .ZN(n8001) );
  ND4D1BWP30P140LVT U8612 ( .A1(n8004), .A2(n8003), .A3(n8002), .A4(n8001), 
        .ZN(n8012) );
  MOAI22D1BWP30P140LVT U8613 ( .A1(n8005), .A2(n8714), .B1(i_data_bus[156]), 
        .B2(n8688), .ZN(n8011) );
  AOI22D1BWP30P140LVT U8614 ( .A1(i_data_bus[508]), .A2(n8718), .B1(
        i_data_bus[412]), .B2(n8719), .ZN(n8009) );
  AOI22D1BWP30P140LVT U8615 ( .A1(i_data_bus[444]), .A2(n8717), .B1(
        i_data_bus[220]), .B2(n8713), .ZN(n8008) );
  AOI22D1BWP30P140LVT U8616 ( .A1(i_data_bus[604]), .A2(n8722), .B1(
        i_data_bus[572]), .B2(n8723), .ZN(n8007) );
  AOI22D1BWP30P140LVT U8617 ( .A1(i_data_bus[540]), .A2(n8721), .B1(
        i_data_bus[636]), .B2(n8720), .ZN(n8006) );
  ND4D1BWP30P140LVT U8618 ( .A1(n8009), .A2(n8008), .A3(n8007), .A4(n8006), 
        .ZN(n8010) );
  NR4D0BWP30P140LVT U8619 ( .A1(n8013), .A2(n8012), .A3(n8011), .A4(n8010), 
        .ZN(n8014) );
  ND4D4BWP30P140LVT U8620 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), 
        .ZN(o_data_bus[188]) );
  AOI22D1BWP30P140LVT U8621 ( .A1(i_data_bus[922]), .A2(n8686), .B1(
        i_data_bus[378]), .B2(n8701), .ZN(n8037) );
  AOI22D1BWP30P140LVT U8622 ( .A1(i_data_bus[954]), .A2(n8704), .B1(
        i_data_bus[986]), .B2(n8708), .ZN(n8036) );
  AOI22D1BWP30P140LVT U8623 ( .A1(i_data_bus[250]), .A2(n8687), .B1(
        i_data_bus[474]), .B2(n8626), .ZN(n8035) );
  AOI22D1BWP30P140LVT U8624 ( .A1(i_data_bus[858]), .A2(n8690), .B1(
        i_data_bus[346]), .B2(n8685), .ZN(n8021) );
  AOI22D1BWP30P140LVT U8625 ( .A1(i_data_bus[58]), .A2(n8684), .B1(
        i_data_bus[826]), .B2(n8695), .ZN(n8020) );
  AOI22D1BWP30P140LVT U8626 ( .A1(i_data_bus[90]), .A2(n8694), .B1(
        i_data_bus[762]), .B2(n8696), .ZN(n8019) );
  AOI22D1BWP30P140LVT U8627 ( .A1(i_data_bus[1018]), .A2(n8702), .B1(
        i_data_bus[666]), .B2(n8693), .ZN(n8018) );
  ND4D1BWP30P140LVT U8628 ( .A1(n8021), .A2(n8020), .A3(n8019), .A4(n8018), 
        .ZN(n8033) );
  AOI22D1BWP30P140LVT U8629 ( .A1(i_data_bus[122]), .A2(n8692), .B1(
        i_data_bus[314]), .B2(n8705), .ZN(n8025) );
  AOI22D1BWP30P140LVT U8630 ( .A1(i_data_bus[890]), .A2(n8706), .B1(
        i_data_bus[730]), .B2(n8703), .ZN(n8024) );
  AOI22D1BWP30P140LVT U8631 ( .A1(i_data_bus[282]), .A2(n8691), .B1(
        i_data_bus[794]), .B2(n8707), .ZN(n8023) );
  AOI22D1BWP30P140LVT U8632 ( .A1(i_data_bus[26]), .A2(n8683), .B1(
        i_data_bus[698]), .B2(n8689), .ZN(n8022) );
  ND4D1BWP30P140LVT U8633 ( .A1(n8025), .A2(n8024), .A3(n8023), .A4(n8022), 
        .ZN(n8032) );
  MOAI22D1BWP30P140LVT U8634 ( .A1(n9627), .A2(n8647), .B1(i_data_bus[186]), 
        .B2(n8716), .ZN(n8031) );
  AOI22D1BWP30P140LVT U8635 ( .A1(i_data_bus[442]), .A2(n8717), .B1(
        i_data_bus[154]), .B2(n8688), .ZN(n8029) );
  AOI22D1BWP30P140LVT U8636 ( .A1(i_data_bus[218]), .A2(n8713), .B1(
        i_data_bus[506]), .B2(n8718), .ZN(n8028) );
  AOI22D1BWP30P140LVT U8637 ( .A1(i_data_bus[634]), .A2(n8720), .B1(
        i_data_bus[570]), .B2(n8723), .ZN(n8027) );
  AOI22D1BWP30P140LVT U8638 ( .A1(i_data_bus[602]), .A2(n8722), .B1(
        i_data_bus[538]), .B2(n8721), .ZN(n8026) );
  ND4D1BWP30P140LVT U8639 ( .A1(n8029), .A2(n8028), .A3(n8027), .A4(n8026), 
        .ZN(n8030) );
  NR4D0BWP30P140LVT U8640 ( .A1(n8033), .A2(n8032), .A3(n8031), .A4(n8030), 
        .ZN(n8034) );
  ND4D4BWP30P140LVT U8641 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), 
        .ZN(o_data_bus[186]) );
  AOI22D1BWP30P140LVT U8642 ( .A1(i_data_bus[984]), .A2(n8708), .B1(
        i_data_bus[120]), .B2(n8692), .ZN(n8058) );
  AOI22D1BWP30P140LVT U8643 ( .A1(i_data_bus[280]), .A2(n8691), .B1(
        i_data_bus[792]), .B2(n8707), .ZN(n8057) );
  AOI22D1BWP30P140LVT U8644 ( .A1(i_data_bus[248]), .A2(n8687), .B1(
        i_data_bus[472]), .B2(n8626), .ZN(n8056) );
  AOI22D1BWP30P140LVT U8645 ( .A1(i_data_bus[696]), .A2(n8689), .B1(
        i_data_bus[824]), .B2(n8695), .ZN(n8041) );
  AOI22D1BWP30P140LVT U8646 ( .A1(i_data_bus[24]), .A2(n8683), .B1(
        i_data_bus[760]), .B2(n8696), .ZN(n8040) );
  AOI22D1BWP30P140LVT U8647 ( .A1(i_data_bus[344]), .A2(n8685), .B1(
        i_data_bus[312]), .B2(n8705), .ZN(n8039) );
  AOI22D1BWP30P140LVT U8648 ( .A1(i_data_bus[1016]), .A2(n8702), .B1(
        i_data_bus[856]), .B2(n8690), .ZN(n8038) );
  ND4D1BWP30P140LVT U8649 ( .A1(n8041), .A2(n8040), .A3(n8039), .A4(n8038), 
        .ZN(n8054) );
  AOI22D1BWP30P140LVT U8650 ( .A1(i_data_bus[376]), .A2(n8701), .B1(
        i_data_bus[888]), .B2(n8706), .ZN(n8045) );
  AOI22D1BWP30P140LVT U8651 ( .A1(i_data_bus[88]), .A2(n8694), .B1(
        i_data_bus[952]), .B2(n8704), .ZN(n8044) );
  AOI22D1BWP30P140LVT U8652 ( .A1(i_data_bus[56]), .A2(n8684), .B1(
        i_data_bus[728]), .B2(n8703), .ZN(n8043) );
  AOI22D1BWP30P140LVT U8653 ( .A1(i_data_bus[920]), .A2(n8686), .B1(
        i_data_bus[664]), .B2(n8693), .ZN(n8042) );
  ND4D1BWP30P140LVT U8654 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), 
        .ZN(n8053) );
  MOAI22D1BWP30P140LVT U8655 ( .A1(n8046), .A2(n8624), .B1(i_data_bus[408]), 
        .B2(n8719), .ZN(n8052) );
  AOI22D1BWP30P140LVT U8656 ( .A1(i_data_bus[152]), .A2(n8688), .B1(
        i_data_bus[216]), .B2(n8713), .ZN(n8050) );
  AOI22D1BWP30P140LVT U8657 ( .A1(i_data_bus[440]), .A2(n8717), .B1(
        i_data_bus[184]), .B2(n8716), .ZN(n8049) );
  AOI22D1BWP30P140LVT U8658 ( .A1(i_data_bus[600]), .A2(n8722), .B1(
        i_data_bus[536]), .B2(n8721), .ZN(n8048) );
  AOI22D1BWP30P140LVT U8659 ( .A1(i_data_bus[632]), .A2(n8720), .B1(
        i_data_bus[568]), .B2(n8723), .ZN(n8047) );
  ND4D1BWP30P140LVT U8660 ( .A1(n8050), .A2(n8049), .A3(n8048), .A4(n8047), 
        .ZN(n8051) );
  NR4D0BWP30P140LVT U8661 ( .A1(n8054), .A2(n8053), .A3(n8052), .A4(n8051), 
        .ZN(n8055) );
  ND4D4BWP30P140LVT U8662 ( .A1(n8058), .A2(n8057), .A3(n8056), .A4(n8055), 
        .ZN(o_data_bus[184]) );
  AOI22D1BWP30P140LVT U8663 ( .A1(i_data_bus[1015]), .A2(n8702), .B1(
        i_data_bus[87]), .B2(n8694), .ZN(n8078) );
  AOI22D1BWP30P140LVT U8664 ( .A1(i_data_bus[919]), .A2(n8686), .B1(
        i_data_bus[279]), .B2(n8691), .ZN(n8077) );
  AOI22D1BWP30P140LVT U8665 ( .A1(i_data_bus[247]), .A2(n8687), .B1(
        i_data_bus[439]), .B2(n8717), .ZN(n8076) );
  AOI22D1BWP30P140LVT U8666 ( .A1(i_data_bus[695]), .A2(n8689), .B1(
        i_data_bus[663]), .B2(n8693), .ZN(n8062) );
  AOI22D1BWP30P140LVT U8667 ( .A1(i_data_bus[311]), .A2(n8705), .B1(
        i_data_bus[375]), .B2(n8701), .ZN(n8061) );
  AOI22D1BWP30P140LVT U8668 ( .A1(i_data_bus[983]), .A2(n8708), .B1(
        i_data_bus[823]), .B2(n8695), .ZN(n8060) );
  AOI22D1BWP30P140LVT U8669 ( .A1(i_data_bus[55]), .A2(n8684), .B1(
        i_data_bus[887]), .B2(n8706), .ZN(n8059) );
  ND4D1BWP30P140LVT U8670 ( .A1(n8062), .A2(n8061), .A3(n8060), .A4(n8059), 
        .ZN(n8074) );
  AOI22D1BWP30P140LVT U8671 ( .A1(i_data_bus[23]), .A2(n8683), .B1(
        i_data_bus[791]), .B2(n8707), .ZN(n8066) );
  AOI22D1BWP30P140LVT U8672 ( .A1(i_data_bus[119]), .A2(n8692), .B1(
        i_data_bus[727]), .B2(n8703), .ZN(n8065) );
  AOI22D1BWP30P140LVT U8673 ( .A1(i_data_bus[951]), .A2(n8704), .B1(
        i_data_bus[343]), .B2(n8685), .ZN(n8064) );
  AOI22D1BWP30P140LVT U8674 ( .A1(i_data_bus[759]), .A2(n8696), .B1(
        i_data_bus[855]), .B2(n8690), .ZN(n8063) );
  ND4D1BWP30P140LVT U8675 ( .A1(n8066), .A2(n8065), .A3(n8064), .A4(n8063), 
        .ZN(n8073) );
  MOAI22D1BWP30P140LVT U8676 ( .A1(n8950), .A2(n8714), .B1(i_data_bus[183]), 
        .B2(n8716), .ZN(n8072) );
  AOI22D1BWP30P140LVT U8677 ( .A1(i_data_bus[151]), .A2(n8688), .B1(
        i_data_bus[407]), .B2(n8719), .ZN(n8070) );
  AOI22D1BWP30P140LVT U8678 ( .A1(i_data_bus[215]), .A2(n8713), .B1(
        i_data_bus[503]), .B2(n8718), .ZN(n8069) );
  AOI22D1BWP30P140LVT U8679 ( .A1(i_data_bus[631]), .A2(n8720), .B1(
        i_data_bus[567]), .B2(n8723), .ZN(n8068) );
  AOI22D1BWP30P140LVT U8680 ( .A1(i_data_bus[599]), .A2(n8722), .B1(
        i_data_bus[535]), .B2(n8721), .ZN(n8067) );
  ND4D1BWP30P140LVT U8681 ( .A1(n8070), .A2(n8069), .A3(n8068), .A4(n8067), 
        .ZN(n8071) );
  NR4D0BWP30P140LVT U8682 ( .A1(n8074), .A2(n8073), .A3(n8072), .A4(n8071), 
        .ZN(n8075) );
  ND4D4BWP30P140LVT U8683 ( .A1(n8078), .A2(n8077), .A3(n8076), .A4(n8075), 
        .ZN(o_data_bus[183]) );
  AOI22D1BWP30P140LVT U8684 ( .A1(i_data_bus[1014]), .A2(n8702), .B1(
        i_data_bus[918]), .B2(n8686), .ZN(n8098) );
  AOI22D1BWP30P140LVT U8685 ( .A1(i_data_bus[86]), .A2(n8694), .B1(
        i_data_bus[726]), .B2(n8703), .ZN(n8097) );
  AOI22D1BWP30P140LVT U8686 ( .A1(i_data_bus[246]), .A2(n8687), .B1(
        i_data_bus[502]), .B2(n8718), .ZN(n8096) );
  AOI22D1BWP30P140LVT U8687 ( .A1(i_data_bus[982]), .A2(n8708), .B1(
        i_data_bus[662]), .B2(n8693), .ZN(n8082) );
  AOI22D1BWP30P140LVT U8688 ( .A1(i_data_bus[118]), .A2(n8692), .B1(
        i_data_bus[310]), .B2(n8705), .ZN(n8081) );
  AOI22D1BWP30P140LVT U8689 ( .A1(i_data_bus[886]), .A2(n8706), .B1(
        i_data_bus[342]), .B2(n8685), .ZN(n8080) );
  AOI22D1BWP30P140LVT U8690 ( .A1(i_data_bus[22]), .A2(n8683), .B1(
        i_data_bus[822]), .B2(n8695), .ZN(n8079) );
  ND4D1BWP30P140LVT U8691 ( .A1(n8082), .A2(n8081), .A3(n8080), .A4(n8079), 
        .ZN(n8094) );
  AOI22D1BWP30P140LVT U8692 ( .A1(i_data_bus[374]), .A2(n8701), .B1(
        i_data_bus[278]), .B2(n8691), .ZN(n8086) );
  AOI22D1BWP30P140LVT U8693 ( .A1(i_data_bus[694]), .A2(n8689), .B1(
        i_data_bus[854]), .B2(n8690), .ZN(n8085) );
  AOI22D1BWP30P140LVT U8694 ( .A1(i_data_bus[950]), .A2(n8704), .B1(
        i_data_bus[758]), .B2(n8696), .ZN(n8084) );
  AOI22D1BWP30P140LVT U8695 ( .A1(i_data_bus[54]), .A2(n8684), .B1(
        i_data_bus[790]), .B2(n8707), .ZN(n8083) );
  ND4D1BWP30P140LVT U8696 ( .A1(n8086), .A2(n8085), .A3(n8084), .A4(n8083), 
        .ZN(n8093) );
  INVD1BWP30P140LVT U8697 ( .I(i_data_bus[214]), .ZN(n9075) );
  OAI22D1BWP30P140LVT U8698 ( .A1(n8804), .A2(n8714), .B1(n9075), .B2(n8623), 
        .ZN(n8092) );
  AOI22D1BWP30P140LVT U8699 ( .A1(i_data_bus[182]), .A2(n8716), .B1(
        i_data_bus[150]), .B2(n8688), .ZN(n8090) );
  AOI22D1BWP30P140LVT U8700 ( .A1(i_data_bus[438]), .A2(n8717), .B1(
        i_data_bus[406]), .B2(n8719), .ZN(n8089) );
  AOI22D1BWP30P140LVT U8701 ( .A1(i_data_bus[534]), .A2(n8721), .B1(
        i_data_bus[630]), .B2(n8720), .ZN(n8088) );
  AOI22D1BWP30P140LVT U8702 ( .A1(i_data_bus[566]), .A2(n8723), .B1(
        i_data_bus[598]), .B2(n8722), .ZN(n8087) );
  ND4D1BWP30P140LVT U8703 ( .A1(n8090), .A2(n8089), .A3(n8088), .A4(n8087), 
        .ZN(n8091) );
  NR4D0BWP30P140LVT U8704 ( .A1(n8094), .A2(n8093), .A3(n8092), .A4(n8091), 
        .ZN(n8095) );
  ND4D4BWP30P140LVT U8705 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), 
        .ZN(o_data_bus[182]) );
  AOI22D1BWP30P140LVT U8706 ( .A1(i_data_bus[981]), .A2(n8708), .B1(
        i_data_bus[885]), .B2(n8706), .ZN(n8119) );
  AOI22D1BWP30P140LVT U8707 ( .A1(i_data_bus[85]), .A2(n8694), .B1(
        i_data_bus[1013]), .B2(n8702), .ZN(n8118) );
  AOI22D1BWP30P140LVT U8708 ( .A1(i_data_bus[181]), .A2(n8716), .B1(
        i_data_bus[469]), .B2(n8626), .ZN(n8117) );
  AOI22D1BWP30P140LVT U8709 ( .A1(i_data_bus[341]), .A2(n8685), .B1(
        i_data_bus[725]), .B2(n8703), .ZN(n8102) );
  AOI22D1BWP30P140LVT U8710 ( .A1(i_data_bus[21]), .A2(n8683), .B1(
        i_data_bus[661]), .B2(n8693), .ZN(n8101) );
  AOI22D1BWP30P140LVT U8711 ( .A1(i_data_bus[949]), .A2(n8704), .B1(
        i_data_bus[693]), .B2(n8689), .ZN(n8100) );
  AOI22D1BWP30P140LVT U8712 ( .A1(i_data_bus[53]), .A2(n8684), .B1(
        i_data_bus[117]), .B2(n8692), .ZN(n8099) );
  ND4D1BWP30P140LVT U8713 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), 
        .ZN(n8115) );
  AOI22D1BWP30P140LVT U8714 ( .A1(i_data_bus[917]), .A2(n8686), .B1(
        i_data_bus[789]), .B2(n8707), .ZN(n8106) );
  AOI22D1BWP30P140LVT U8715 ( .A1(i_data_bus[277]), .A2(n8691), .B1(
        i_data_bus[373]), .B2(n8701), .ZN(n8105) );
  AOI22D1BWP30P140LVT U8716 ( .A1(i_data_bus[757]), .A2(n8696), .B1(
        i_data_bus[821]), .B2(n8695), .ZN(n8104) );
  AOI22D1BWP30P140LVT U8717 ( .A1(i_data_bus[853]), .A2(n8690), .B1(
        i_data_bus[309]), .B2(n8705), .ZN(n8103) );
  ND4D1BWP30P140LVT U8718 ( .A1(n8106), .A2(n8105), .A3(n8104), .A4(n8103), 
        .ZN(n8114) );
  MOAI22D1BWP30P140LVT U8719 ( .A1(n8107), .A2(n8647), .B1(i_data_bus[149]), 
        .B2(n8688), .ZN(n8113) );
  AOI22D1BWP30P140LVT U8720 ( .A1(i_data_bus[437]), .A2(n8717), .B1(
        i_data_bus[245]), .B2(n8687), .ZN(n8111) );
  AOI22D1BWP30P140LVT U8721 ( .A1(i_data_bus[501]), .A2(n8718), .B1(
        i_data_bus[213]), .B2(n8713), .ZN(n8110) );
  AOI22D1BWP30P140LVT U8722 ( .A1(i_data_bus[597]), .A2(n8722), .B1(
        i_data_bus[533]), .B2(n8721), .ZN(n8109) );
  AOI22D1BWP30P140LVT U8723 ( .A1(i_data_bus[629]), .A2(n8720), .B1(
        i_data_bus[565]), .B2(n8723), .ZN(n8108) );
  ND4D1BWP30P140LVT U8724 ( .A1(n8111), .A2(n8110), .A3(n8109), .A4(n8108), 
        .ZN(n8112) );
  NR4D0BWP30P140LVT U8725 ( .A1(n8115), .A2(n8114), .A3(n8113), .A4(n8112), 
        .ZN(n8116) );
  ND4D4BWP30P140LVT U8726 ( .A1(n8119), .A2(n8118), .A3(n8117), .A4(n8116), 
        .ZN(o_data_bus[181]) );
  AOI22D1BWP30P140LVT U8727 ( .A1(i_data_bus[948]), .A2(n8704), .B1(
        i_data_bus[84]), .B2(n8694), .ZN(n8140) );
  AOI22D1BWP30P140LVT U8728 ( .A1(i_data_bus[1012]), .A2(n8702), .B1(
        i_data_bus[884]), .B2(n8706), .ZN(n8139) );
  AOI22D1BWP30P140LVT U8729 ( .A1(i_data_bus[244]), .A2(n8687), .B1(
        i_data_bus[436]), .B2(n8717), .ZN(n8138) );
  AOI22D1BWP30P140LVT U8730 ( .A1(i_data_bus[276]), .A2(n8691), .B1(
        i_data_bus[660]), .B2(n8693), .ZN(n8123) );
  AOI22D1BWP30P140LVT U8731 ( .A1(i_data_bus[52]), .A2(n8684), .B1(
        i_data_bus[692]), .B2(n8689), .ZN(n8122) );
  AOI22D1BWP30P140LVT U8732 ( .A1(i_data_bus[980]), .A2(n8708), .B1(
        i_data_bus[116]), .B2(n8692), .ZN(n8121) );
  AOI22D1BWP30P140LVT U8733 ( .A1(i_data_bus[916]), .A2(n8686), .B1(
        i_data_bus[724]), .B2(n8703), .ZN(n8120) );
  ND4D1BWP30P140LVT U8734 ( .A1(n8123), .A2(n8122), .A3(n8121), .A4(n8120), 
        .ZN(n8136) );
  AOI22D1BWP30P140LVT U8735 ( .A1(i_data_bus[340]), .A2(n8685), .B1(
        i_data_bus[820]), .B2(n8695), .ZN(n8127) );
  AOI22D1BWP30P140LVT U8736 ( .A1(i_data_bus[20]), .A2(n8683), .B1(
        i_data_bus[756]), .B2(n8696), .ZN(n8126) );
  AOI22D1BWP30P140LVT U8737 ( .A1(i_data_bus[852]), .A2(n8690), .B1(
        i_data_bus[372]), .B2(n8701), .ZN(n8125) );
  AOI22D1BWP30P140LVT U8738 ( .A1(i_data_bus[788]), .A2(n8707), .B1(
        i_data_bus[308]), .B2(n8705), .ZN(n8124) );
  ND4D1BWP30P140LVT U8739 ( .A1(n8127), .A2(n8126), .A3(n8125), .A4(n8124), 
        .ZN(n8135) );
  MOAI22D1BWP30P140LVT U8740 ( .A1(n8128), .A2(n8714), .B1(i_data_bus[212]), 
        .B2(n8713), .ZN(n8134) );
  AOI22D1BWP30P140LVT U8741 ( .A1(i_data_bus[404]), .A2(n8719), .B1(
        i_data_bus[148]), .B2(n8688), .ZN(n8132) );
  AOI22D1BWP30P140LVT U8742 ( .A1(i_data_bus[180]), .A2(n8716), .B1(
        i_data_bus[500]), .B2(n8718), .ZN(n8131) );
  AOI22D1BWP30P140LVT U8743 ( .A1(i_data_bus[532]), .A2(n8721), .B1(
        i_data_bus[628]), .B2(n8720), .ZN(n8130) );
  AOI22D1BWP30P140LVT U8744 ( .A1(i_data_bus[596]), .A2(n8722), .B1(
        i_data_bus[564]), .B2(n8723), .ZN(n8129) );
  ND4D1BWP30P140LVT U8745 ( .A1(n8132), .A2(n8131), .A3(n8130), .A4(n8129), 
        .ZN(n8133) );
  NR4D0BWP30P140LVT U8746 ( .A1(n8136), .A2(n8135), .A3(n8134), .A4(n8133), 
        .ZN(n8137) );
  ND4D4BWP30P140LVT U8747 ( .A1(n8140), .A2(n8139), .A3(n8138), .A4(n8137), 
        .ZN(o_data_bus[180]) );
  AOI22D1BWP30P140LVT U8748 ( .A1(i_data_bus[339]), .A2(n8685), .B1(
        i_data_bus[851]), .B2(n8690), .ZN(n8160) );
  AOI22D1BWP30P140LVT U8749 ( .A1(i_data_bus[83]), .A2(n8694), .B1(
        i_data_bus[659]), .B2(n8693), .ZN(n8159) );
  AOI22D1BWP30P140LVT U8750 ( .A1(i_data_bus[211]), .A2(n8713), .B1(
        i_data_bus[467]), .B2(n8626), .ZN(n8158) );
  AOI22D1BWP30P140LVT U8751 ( .A1(i_data_bus[179]), .A2(n8716), .B1(
        i_data_bus[147]), .B2(n8688), .ZN(n8156) );
  AOI22D1BWP30P140LVT U8752 ( .A1(i_data_bus[115]), .A2(n8692), .B1(
        i_data_bus[275]), .B2(n8691), .ZN(n8144) );
  AOI22D1BWP30P140LVT U8753 ( .A1(i_data_bus[307]), .A2(n8705), .B1(
        i_data_bus[819]), .B2(n8695), .ZN(n8143) );
  AOI22D1BWP30P140LVT U8754 ( .A1(i_data_bus[947]), .A2(n8704), .B1(
        i_data_bus[787]), .B2(n8707), .ZN(n8142) );
  AOI22D1BWP30P140LVT U8755 ( .A1(i_data_bus[979]), .A2(n8708), .B1(
        i_data_bus[883]), .B2(n8706), .ZN(n8141) );
  ND4D1BWP30P140LVT U8756 ( .A1(n8144), .A2(n8143), .A3(n8142), .A4(n8141), 
        .ZN(n8155) );
  AOI22D1BWP30P140LVT U8757 ( .A1(i_data_bus[19]), .A2(n8683), .B1(
        i_data_bus[691]), .B2(n8689), .ZN(n8148) );
  AOI22D1BWP30P140LVT U8758 ( .A1(i_data_bus[915]), .A2(n8686), .B1(
        i_data_bus[755]), .B2(n8696), .ZN(n8147) );
  AOI22D1BWP30P140LVT U8759 ( .A1(i_data_bus[51]), .A2(n8684), .B1(
        i_data_bus[723]), .B2(n8703), .ZN(n8146) );
  AOI22D1BWP30P140LVT U8760 ( .A1(i_data_bus[1011]), .A2(n8702), .B1(
        i_data_bus[371]), .B2(n8701), .ZN(n8145) );
  ND4D1BWP30P140LVT U8761 ( .A1(n8148), .A2(n8147), .A3(n8146), .A4(n8145), 
        .ZN(n8154) );
  AOI22D1BWP30P140LVT U8762 ( .A1(i_data_bus[243]), .A2(n8687), .B1(
        i_data_bus[435]), .B2(n8717), .ZN(n8152) );
  AOI22D1BWP30P140LVT U8763 ( .A1(i_data_bus[403]), .A2(n8719), .B1(
        i_data_bus[499]), .B2(n8718), .ZN(n8151) );
  AOI22D1BWP30P140LVT U8764 ( .A1(i_data_bus[531]), .A2(n8721), .B1(
        i_data_bus[595]), .B2(n8722), .ZN(n8150) );
  AOI22D1BWP30P140LVT U8765 ( .A1(i_data_bus[563]), .A2(n8723), .B1(
        i_data_bus[627]), .B2(n8720), .ZN(n8149) );
  ND4D1BWP30P140LVT U8766 ( .A1(n8152), .A2(n8151), .A3(n8150), .A4(n8149), 
        .ZN(n8153) );
  INR4D0BWP30P140LVT U8767 ( .A1(n8156), .B1(n8155), .B2(n8154), .B3(n8153), 
        .ZN(n8157) );
  ND4D4BWP30P140LVT U8768 ( .A1(n8160), .A2(n8159), .A3(n8158), .A4(n8157), 
        .ZN(o_data_bus[179]) );
  AOI22D1BWP30P140LVT U8769 ( .A1(i_data_bus[1010]), .A2(n8702), .B1(
        i_data_bus[722]), .B2(n8703), .ZN(n8180) );
  AOI22D1BWP30P140LVT U8770 ( .A1(i_data_bus[818]), .A2(n8695), .B1(
        i_data_bus[338]), .B2(n8685), .ZN(n8179) );
  AOI22D1BWP30P140LVT U8771 ( .A1(i_data_bus[210]), .A2(n8713), .B1(
        i_data_bus[498]), .B2(n8718), .ZN(n8178) );
  AOI22D1BWP30P140LVT U8772 ( .A1(i_data_bus[946]), .A2(n8704), .B1(
        i_data_bus[370]), .B2(n8701), .ZN(n8164) );
  AOI22D1BWP30P140LVT U8773 ( .A1(i_data_bus[50]), .A2(n8684), .B1(
        i_data_bus[914]), .B2(n8686), .ZN(n8163) );
  AOI22D1BWP30P140LVT U8774 ( .A1(i_data_bus[882]), .A2(n8706), .B1(
        i_data_bus[658]), .B2(n8693), .ZN(n8162) );
  AOI22D1BWP30P140LVT U8775 ( .A1(i_data_bus[274]), .A2(n8691), .B1(
        i_data_bus[754]), .B2(n8696), .ZN(n8161) );
  ND4D1BWP30P140LVT U8776 ( .A1(n8164), .A2(n8163), .A3(n8162), .A4(n8161), 
        .ZN(n8176) );
  AOI22D1BWP30P140LVT U8777 ( .A1(i_data_bus[306]), .A2(n8705), .B1(
        i_data_bus[786]), .B2(n8707), .ZN(n8168) );
  AOI22D1BWP30P140LVT U8778 ( .A1(i_data_bus[978]), .A2(n8708), .B1(
        i_data_bus[690]), .B2(n8689), .ZN(n8167) );
  AOI22D1BWP30P140LVT U8779 ( .A1(i_data_bus[114]), .A2(n8692), .B1(
        i_data_bus[82]), .B2(n8694), .ZN(n8166) );
  AOI22D1BWP30P140LVT U8780 ( .A1(i_data_bus[18]), .A2(n8683), .B1(
        i_data_bus[850]), .B2(n8690), .ZN(n8165) );
  ND4D1BWP30P140LVT U8781 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), 
        .ZN(n8175) );
  INVD1BWP30P140LVT U8782 ( .I(i_data_bus[146]), .ZN(n9160) );
  INVD1BWP30P140LVT U8783 ( .I(n8688), .ZN(n8670) );
  MOAI22D1BWP30P140LVT U8784 ( .A1(n9160), .A2(n8670), .B1(i_data_bus[178]), 
        .B2(n8716), .ZN(n8174) );
  AOI22D1BWP30P140LVT U8785 ( .A1(i_data_bus[402]), .A2(n8719), .B1(
        i_data_bus[242]), .B2(n8687), .ZN(n8172) );
  AOI22D1BWP30P140LVT U8786 ( .A1(i_data_bus[466]), .A2(n8626), .B1(
        i_data_bus[434]), .B2(n8717), .ZN(n8171) );
  AOI22D1BWP30P140LVT U8787 ( .A1(i_data_bus[594]), .A2(n8722), .B1(
        i_data_bus[530]), .B2(n8721), .ZN(n8170) );
  AOI22D1BWP30P140LVT U8788 ( .A1(i_data_bus[626]), .A2(n8720), .B1(
        i_data_bus[562]), .B2(n8723), .ZN(n8169) );
  ND4D1BWP30P140LVT U8789 ( .A1(n8172), .A2(n8171), .A3(n8170), .A4(n8169), 
        .ZN(n8173) );
  NR4D0BWP30P140LVT U8790 ( .A1(n8176), .A2(n8175), .A3(n8174), .A4(n8173), 
        .ZN(n8177) );
  ND4D4BWP30P140LVT U8791 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n8177), 
        .ZN(o_data_bus[178]) );
  AOI22D1BWP30P140LVT U8792 ( .A1(i_data_bus[337]), .A2(n8685), .B1(
        i_data_bus[273]), .B2(n8691), .ZN(n8200) );
  AOI22D1BWP30P140LVT U8793 ( .A1(i_data_bus[945]), .A2(n8704), .B1(
        i_data_bus[113]), .B2(n8692), .ZN(n8199) );
  AOI22D1BWP30P140LVT U8794 ( .A1(i_data_bus[433]), .A2(n8717), .B1(
        i_data_bus[497]), .B2(n8718), .ZN(n8198) );
  AOI22D1BWP30P140LVT U8795 ( .A1(i_data_bus[209]), .A2(n8713), .B1(
        i_data_bus[177]), .B2(n8716), .ZN(n8196) );
  AOI22D1BWP30P140LVT U8796 ( .A1(i_data_bus[49]), .A2(n8684), .B1(
        i_data_bus[849]), .B2(n8690), .ZN(n8184) );
  AOI22D1BWP30P140LVT U8797 ( .A1(i_data_bus[1009]), .A2(n8702), .B1(
        i_data_bus[817]), .B2(n8695), .ZN(n8183) );
  AOI22D1BWP30P140LVT U8798 ( .A1(i_data_bus[17]), .A2(n8683), .B1(
        i_data_bus[305]), .B2(n8705), .ZN(n8182) );
  AOI22D1BWP30P140LVT U8799 ( .A1(i_data_bus[689]), .A2(n8689), .B1(
        i_data_bus[753]), .B2(n8696), .ZN(n8181) );
  ND4D1BWP30P140LVT U8800 ( .A1(n8184), .A2(n8183), .A3(n8182), .A4(n8181), 
        .ZN(n8195) );
  AOI22D1BWP30P140LVT U8801 ( .A1(i_data_bus[977]), .A2(n8708), .B1(
        i_data_bus[721]), .B2(n8703), .ZN(n8188) );
  AOI22D1BWP30P140LVT U8802 ( .A1(i_data_bus[81]), .A2(n8694), .B1(
        i_data_bus[657]), .B2(n8693), .ZN(n8187) );
  AOI22D1BWP30P140LVT U8803 ( .A1(i_data_bus[913]), .A2(n8686), .B1(
        i_data_bus[881]), .B2(n8706), .ZN(n8186) );
  AOI22D1BWP30P140LVT U8804 ( .A1(i_data_bus[785]), .A2(n8707), .B1(
        i_data_bus[369]), .B2(n8701), .ZN(n8185) );
  ND4D1BWP30P140LVT U8805 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), 
        .ZN(n8194) );
  AOI22D1BWP30P140LVT U8806 ( .A1(i_data_bus[145]), .A2(n8688), .B1(
        i_data_bus[241]), .B2(n8687), .ZN(n8192) );
  AOI22D1BWP30P140LVT U8807 ( .A1(i_data_bus[401]), .A2(n8719), .B1(
        i_data_bus[465]), .B2(n8626), .ZN(n8191) );
  AOI22D1BWP30P140LVT U8808 ( .A1(i_data_bus[593]), .A2(n8722), .B1(
        i_data_bus[561]), .B2(n8723), .ZN(n8190) );
  AOI22D1BWP30P140LVT U8809 ( .A1(i_data_bus[625]), .A2(n8720), .B1(
        i_data_bus[529]), .B2(n8721), .ZN(n8189) );
  ND4D1BWP30P140LVT U8810 ( .A1(n8192), .A2(n8191), .A3(n8190), .A4(n8189), 
        .ZN(n8193) );
  INR4D0BWP30P140LVT U8811 ( .A1(n8196), .B1(n8195), .B2(n8194), .B3(n8193), 
        .ZN(n8197) );
  ND4D4BWP30P140LVT U8812 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), 
        .ZN(o_data_bus[177]) );
  AOI22D1BWP30P140LVT U8813 ( .A1(i_data_bus[112]), .A2(n8692), .B1(
        i_data_bus[752]), .B2(n8696), .ZN(n8221) );
  AOI22D1BWP30P140LVT U8814 ( .A1(i_data_bus[16]), .A2(n8683), .B1(
        i_data_bus[1008]), .B2(n8702), .ZN(n8220) );
  AOI22D1BWP30P140LVT U8815 ( .A1(i_data_bus[432]), .A2(n8717), .B1(
        i_data_bus[240]), .B2(n8687), .ZN(n8219) );
  AOI22D1BWP30P140LVT U8816 ( .A1(i_data_bus[944]), .A2(n8704), .B1(
        i_data_bus[272]), .B2(n8691), .ZN(n8204) );
  AOI22D1BWP30P140LVT U8817 ( .A1(i_data_bus[80]), .A2(n8694), .B1(
        i_data_bus[688]), .B2(n8689), .ZN(n8203) );
  AOI22D1BWP30P140LVT U8818 ( .A1(i_data_bus[656]), .A2(n8693), .B1(
        i_data_bus[816]), .B2(n8695), .ZN(n8202) );
  AOI22D1BWP30P140LVT U8819 ( .A1(i_data_bus[976]), .A2(n8708), .B1(
        i_data_bus[304]), .B2(n8705), .ZN(n8201) );
  ND4D1BWP30P140LVT U8820 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), 
        .ZN(n8217) );
  AOI22D1BWP30P140LVT U8821 ( .A1(i_data_bus[336]), .A2(n8685), .B1(
        i_data_bus[880]), .B2(n8706), .ZN(n8208) );
  AOI22D1BWP30P140LVT U8822 ( .A1(i_data_bus[912]), .A2(n8686), .B1(
        i_data_bus[368]), .B2(n8701), .ZN(n8207) );
  AOI22D1BWP30P140LVT U8823 ( .A1(i_data_bus[784]), .A2(n8707), .B1(
        i_data_bus[848]), .B2(n8690), .ZN(n8206) );
  AOI22D1BWP30P140LVT U8824 ( .A1(i_data_bus[48]), .A2(n8684), .B1(
        i_data_bus[720]), .B2(n8703), .ZN(n8205) );
  ND4D1BWP30P140LVT U8825 ( .A1(n8208), .A2(n8207), .A3(n8206), .A4(n8205), 
        .ZN(n8216) );
  MOAI22D1BWP30P140LVT U8826 ( .A1(n8209), .A2(n8624), .B1(i_data_bus[176]), 
        .B2(n8716), .ZN(n8215) );
  AOI22D1BWP30P140LVT U8827 ( .A1(i_data_bus[144]), .A2(n8688), .B1(
        i_data_bus[400]), .B2(n8719), .ZN(n8213) );
  AOI22D1BWP30P140LVT U8828 ( .A1(i_data_bus[208]), .A2(n8713), .B1(
        i_data_bus[464]), .B2(n8626), .ZN(n8212) );
  AOI22D1BWP30P140LVT U8829 ( .A1(i_data_bus[560]), .A2(n8723), .B1(
        i_data_bus[528]), .B2(n8721), .ZN(n8211) );
  AOI22D1BWP30P140LVT U8830 ( .A1(i_data_bus[624]), .A2(n8720), .B1(
        i_data_bus[592]), .B2(n8722), .ZN(n8210) );
  ND4D1BWP30P140LVT U8831 ( .A1(n8213), .A2(n8212), .A3(n8211), .A4(n8210), 
        .ZN(n8214) );
  NR4D0BWP30P140LVT U8832 ( .A1(n8217), .A2(n8216), .A3(n8215), .A4(n8214), 
        .ZN(n8218) );
  ND4D4BWP30P140LVT U8833 ( .A1(n8221), .A2(n8220), .A3(n8219), .A4(n8218), 
        .ZN(o_data_bus[176]) );
  AOI22D1BWP30P140LVT U8834 ( .A1(i_data_bus[847]), .A2(n8690), .B1(
        i_data_bus[303]), .B2(n8705), .ZN(n8242) );
  AOI22D1BWP30P140LVT U8835 ( .A1(i_data_bus[111]), .A2(n8692), .B1(
        i_data_bus[335]), .B2(n8685), .ZN(n8241) );
  AOI22D1BWP30P140LVT U8836 ( .A1(i_data_bus[239]), .A2(n8687), .B1(
        i_data_bus[495]), .B2(n8718), .ZN(n8240) );
  AOI22D1BWP30P140LVT U8837 ( .A1(i_data_bus[271]), .A2(n8691), .B1(
        i_data_bus[815]), .B2(n8695), .ZN(n8225) );
  AOI22D1BWP30P140LVT U8838 ( .A1(i_data_bus[15]), .A2(n8683), .B1(
        i_data_bus[783]), .B2(n8707), .ZN(n8224) );
  AOI22D1BWP30P140LVT U8839 ( .A1(i_data_bus[911]), .A2(n8686), .B1(
        i_data_bus[879]), .B2(n8706), .ZN(n8223) );
  AOI22D1BWP30P140LVT U8840 ( .A1(i_data_bus[719]), .A2(n8703), .B1(
        i_data_bus[655]), .B2(n8693), .ZN(n8222) );
  ND4D1BWP30P140LVT U8841 ( .A1(n8225), .A2(n8224), .A3(n8223), .A4(n8222), 
        .ZN(n8238) );
  AOI22D1BWP30P140LVT U8842 ( .A1(i_data_bus[975]), .A2(n8708), .B1(
        i_data_bus[367]), .B2(n8701), .ZN(n8229) );
  AOI22D1BWP30P140LVT U8843 ( .A1(i_data_bus[943]), .A2(n8704), .B1(
        i_data_bus[687]), .B2(n8689), .ZN(n8228) );
  AOI22D1BWP30P140LVT U8844 ( .A1(i_data_bus[1007]), .A2(n8702), .B1(
        i_data_bus[751]), .B2(n8696), .ZN(n8227) );
  AOI22D1BWP30P140LVT U8845 ( .A1(i_data_bus[79]), .A2(n8694), .B1(
        i_data_bus[47]), .B2(n8684), .ZN(n8226) );
  ND4D1BWP30P140LVT U8846 ( .A1(n8229), .A2(n8228), .A3(n8227), .A4(n8226), 
        .ZN(n8237) );
  MOAI22D1BWP30P140LVT U8847 ( .A1(n8230), .A2(n8714), .B1(i_data_bus[143]), 
        .B2(n8688), .ZN(n8236) );
  AOI22D1BWP30P140LVT U8848 ( .A1(i_data_bus[431]), .A2(n8717), .B1(
        i_data_bus[399]), .B2(n8719), .ZN(n8234) );
  AOI22D1BWP30P140LVT U8849 ( .A1(i_data_bus[207]), .A2(n8713), .B1(
        i_data_bus[175]), .B2(n8716), .ZN(n8233) );
  AOI22D1BWP30P140LVT U8850 ( .A1(i_data_bus[559]), .A2(n8723), .B1(
        i_data_bus[527]), .B2(n8721), .ZN(n8232) );
  AOI22D1BWP30P140LVT U8851 ( .A1(i_data_bus[591]), .A2(n8722), .B1(
        i_data_bus[623]), .B2(n8720), .ZN(n8231) );
  ND4D1BWP30P140LVT U8852 ( .A1(n8234), .A2(n8233), .A3(n8232), .A4(n8231), 
        .ZN(n8235) );
  NR4D0BWP30P140LVT U8853 ( .A1(n8238), .A2(n8237), .A3(n8236), .A4(n8235), 
        .ZN(n8239) );
  ND4D4BWP30P140LVT U8854 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n8239), 
        .ZN(o_data_bus[175]) );
  AOI22D1BWP30P140LVT U8855 ( .A1(i_data_bus[110]), .A2(n8692), .B1(
        i_data_bus[686]), .B2(n8689), .ZN(n8263) );
  AOI22D1BWP30P140LVT U8856 ( .A1(i_data_bus[302]), .A2(n8705), .B1(
        i_data_bus[718]), .B2(n8703), .ZN(n8262) );
  AOI22D1BWP30P140LVT U8857 ( .A1(i_data_bus[430]), .A2(n8717), .B1(
        i_data_bus[494]), .B2(n8718), .ZN(n8261) );
  AOI22D1BWP30P140LVT U8858 ( .A1(i_data_bus[942]), .A2(n8704), .B1(
        i_data_bus[782]), .B2(n8707), .ZN(n8246) );
  AOI22D1BWP30P140LVT U8859 ( .A1(i_data_bus[910]), .A2(n8686), .B1(
        i_data_bus[878]), .B2(n8706), .ZN(n8245) );
  AOI22D1BWP30P140LVT U8860 ( .A1(i_data_bus[814]), .A2(n8695), .B1(
        i_data_bus[846]), .B2(n8690), .ZN(n8244) );
  AOI22D1BWP30P140LVT U8861 ( .A1(i_data_bus[1006]), .A2(n8702), .B1(
        i_data_bus[46]), .B2(n8684), .ZN(n8243) );
  ND4D1BWP30P140LVT U8862 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), 
        .ZN(n8259) );
  AOI22D1BWP30P140LVT U8863 ( .A1(i_data_bus[974]), .A2(n8708), .B1(
        i_data_bus[270]), .B2(n8691), .ZN(n8250) );
  AOI22D1BWP30P140LVT U8864 ( .A1(i_data_bus[14]), .A2(n8683), .B1(
        i_data_bus[750]), .B2(n8696), .ZN(n8249) );
  AOI22D1BWP30P140LVT U8865 ( .A1(i_data_bus[78]), .A2(n8694), .B1(
        i_data_bus[366]), .B2(n8701), .ZN(n8248) );
  AOI22D1BWP30P140LVT U8866 ( .A1(i_data_bus[334]), .A2(n8685), .B1(
        i_data_bus[654]), .B2(n8693), .ZN(n8247) );
  ND4D1BWP30P140LVT U8867 ( .A1(n8250), .A2(n8249), .A3(n8248), .A4(n8247), 
        .ZN(n8258) );
  MOAI22D1BWP30P140LVT U8868 ( .A1(n8251), .A2(n8647), .B1(i_data_bus[462]), 
        .B2(n8626), .ZN(n8257) );
  AOI22D1BWP30P140LVT U8869 ( .A1(i_data_bus[174]), .A2(n8716), .B1(
        i_data_bus[238]), .B2(n8687), .ZN(n8255) );
  AOI22D1BWP30P140LVT U8870 ( .A1(i_data_bus[206]), .A2(n8713), .B1(
        i_data_bus[142]), .B2(n8688), .ZN(n8254) );
  AOI22D1BWP30P140LVT U8871 ( .A1(i_data_bus[590]), .A2(n8722), .B1(
        i_data_bus[526]), .B2(n8721), .ZN(n8253) );
  AOI22D1BWP30P140LVT U8872 ( .A1(i_data_bus[558]), .A2(n8723), .B1(
        i_data_bus[622]), .B2(n8720), .ZN(n8252) );
  ND4D1BWP30P140LVT U8873 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), 
        .ZN(n8256) );
  NR4D0BWP30P140LVT U8874 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), 
        .ZN(n8260) );
  ND4D4BWP30P140LVT U8875 ( .A1(n8263), .A2(n8262), .A3(n8261), .A4(n8260), 
        .ZN(o_data_bus[174]) );
  AOI22D1BWP30P140LVT U8876 ( .A1(i_data_bus[876]), .A2(n8706), .B1(
        i_data_bus[332]), .B2(n8685), .ZN(n8284) );
  AOI22D1BWP30P140LVT U8877 ( .A1(i_data_bus[12]), .A2(n8683), .B1(
        i_data_bus[972]), .B2(n8708), .ZN(n8283) );
  AOI22D1BWP30P140LVT U8878 ( .A1(i_data_bus[460]), .A2(n8626), .B1(
        i_data_bus[396]), .B2(n8719), .ZN(n8282) );
  AOI22D1BWP30P140LVT U8879 ( .A1(i_data_bus[908]), .A2(n8686), .B1(
        i_data_bus[108]), .B2(n8692), .ZN(n8267) );
  AOI22D1BWP30P140LVT U8880 ( .A1(i_data_bus[76]), .A2(n8694), .B1(
        i_data_bus[844]), .B2(n8690), .ZN(n8266) );
  AOI22D1BWP30P140LVT U8881 ( .A1(i_data_bus[364]), .A2(n8701), .B1(
        i_data_bus[652]), .B2(n8693), .ZN(n8265) );
  AOI22D1BWP30P140LVT U8882 ( .A1(i_data_bus[780]), .A2(n8707), .B1(
        i_data_bus[812]), .B2(n8695), .ZN(n8264) );
  ND4D1BWP30P140LVT U8883 ( .A1(n8267), .A2(n8266), .A3(n8265), .A4(n8264), 
        .ZN(n8280) );
  AOI22D1BWP30P140LVT U8884 ( .A1(i_data_bus[44]), .A2(n8684), .B1(
        i_data_bus[1004]), .B2(n8702), .ZN(n8271) );
  AOI22D1BWP30P140LVT U8885 ( .A1(i_data_bus[940]), .A2(n8704), .B1(
        i_data_bus[300]), .B2(n8705), .ZN(n8270) );
  AOI22D1BWP30P140LVT U8886 ( .A1(i_data_bus[716]), .A2(n8703), .B1(
        i_data_bus[748]), .B2(n8696), .ZN(n8269) );
  AOI22D1BWP30P140LVT U8887 ( .A1(i_data_bus[684]), .A2(n8689), .B1(
        i_data_bus[268]), .B2(n8691), .ZN(n8268) );
  ND4D1BWP30P140LVT U8888 ( .A1(n8271), .A2(n8270), .A3(n8269), .A4(n8268), 
        .ZN(n8279) );
  OAI22D1BWP30P140LVT U8889 ( .A1(n8971), .A2(n8624), .B1(n8272), .B2(n8602), 
        .ZN(n8278) );
  AOI22D1BWP30P140LVT U8890 ( .A1(i_data_bus[204]), .A2(n8713), .B1(
        i_data_bus[236]), .B2(n8687), .ZN(n8276) );
  AOI22D1BWP30P140LVT U8891 ( .A1(i_data_bus[428]), .A2(n8717), .B1(
        i_data_bus[140]), .B2(n8688), .ZN(n8275) );
  AOI22D1BWP30P140LVT U8892 ( .A1(i_data_bus[620]), .A2(n8720), .B1(
        i_data_bus[524]), .B2(n8721), .ZN(n8274) );
  AOI22D1BWP30P140LVT U8893 ( .A1(i_data_bus[556]), .A2(n8723), .B1(
        i_data_bus[588]), .B2(n8722), .ZN(n8273) );
  ND4D1BWP30P140LVT U8894 ( .A1(n8276), .A2(n8275), .A3(n8274), .A4(n8273), 
        .ZN(n8277) );
  NR4D0BWP30P140LVT U8895 ( .A1(n8280), .A2(n8279), .A3(n8278), .A4(n8277), 
        .ZN(n8281) );
  ND4D4BWP30P140LVT U8896 ( .A1(n8284), .A2(n8283), .A3(n8282), .A4(n8281), 
        .ZN(o_data_bus[172]) );
  AOI22D1BWP30P140LVT U8897 ( .A1(i_data_bus[75]), .A2(n8694), .B1(
        i_data_bus[651]), .B2(n8693), .ZN(n8304) );
  AOI22D1BWP30P140LVT U8898 ( .A1(i_data_bus[747]), .A2(n8696), .B1(
        i_data_bus[299]), .B2(n8705), .ZN(n8303) );
  AOI22D1BWP30P140LVT U8899 ( .A1(i_data_bus[203]), .A2(n8713), .B1(
        i_data_bus[139]), .B2(n8688), .ZN(n8302) );
  AOI22D1BWP30P140LVT U8900 ( .A1(i_data_bus[43]), .A2(n8684), .B1(
        i_data_bus[779]), .B2(n8707), .ZN(n8288) );
  AOI22D1BWP30P140LVT U8901 ( .A1(i_data_bus[907]), .A2(n8686), .B1(
        i_data_bus[363]), .B2(n8701), .ZN(n8287) );
  AOI22D1BWP30P140LVT U8902 ( .A1(i_data_bus[107]), .A2(n8692), .B1(
        i_data_bus[683]), .B2(n8689), .ZN(n8286) );
  AOI22D1BWP30P140LVT U8903 ( .A1(i_data_bus[939]), .A2(n8704), .B1(
        i_data_bus[11]), .B2(n8683), .ZN(n8285) );
  ND4D1BWP30P140LVT U8904 ( .A1(n8288), .A2(n8287), .A3(n8286), .A4(n8285), 
        .ZN(n8300) );
  AOI22D1BWP30P140LVT U8905 ( .A1(i_data_bus[875]), .A2(n8706), .B1(
        i_data_bus[715]), .B2(n8703), .ZN(n8292) );
  AOI22D1BWP30P140LVT U8906 ( .A1(i_data_bus[971]), .A2(n8708), .B1(
        i_data_bus[843]), .B2(n8690), .ZN(n8291) );
  AOI22D1BWP30P140LVT U8907 ( .A1(i_data_bus[811]), .A2(n8695), .B1(
        i_data_bus[331]), .B2(n8685), .ZN(n8290) );
  AOI22D1BWP30P140LVT U8908 ( .A1(i_data_bus[1003]), .A2(n8702), .B1(
        i_data_bus[267]), .B2(n8691), .ZN(n8289) );
  ND4D1BWP30P140LVT U8909 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), 
        .ZN(n8299) );
  MOAI22D1BWP30P140LVT U8910 ( .A1(n9650), .A2(n8714), .B1(i_data_bus[171]), 
        .B2(n8716), .ZN(n8298) );
  AOI22D1BWP30P140LVT U8911 ( .A1(i_data_bus[395]), .A2(n8719), .B1(
        i_data_bus[235]), .B2(n8687), .ZN(n8296) );
  AOI22D1BWP30P140LVT U8912 ( .A1(i_data_bus[491]), .A2(n8718), .B1(
        i_data_bus[427]), .B2(n8717), .ZN(n8295) );
  AOI22D1BWP30P140LVT U8913 ( .A1(i_data_bus[619]), .A2(n8720), .B1(
        i_data_bus[587]), .B2(n8722), .ZN(n8294) );
  AOI22D1BWP30P140LVT U8914 ( .A1(i_data_bus[523]), .A2(n8721), .B1(
        i_data_bus[555]), .B2(n8723), .ZN(n8293) );
  ND4D1BWP30P140LVT U8915 ( .A1(n8296), .A2(n8295), .A3(n8294), .A4(n8293), 
        .ZN(n8297) );
  NR4D0BWP30P140LVT U8916 ( .A1(n8300), .A2(n8299), .A3(n8298), .A4(n8297), 
        .ZN(n8301) );
  ND4D4BWP30P140LVT U8917 ( .A1(n8304), .A2(n8303), .A3(n8302), .A4(n8301), 
        .ZN(o_data_bus[171]) );
  AOI22D1BWP30P140LVT U8918 ( .A1(i_data_bus[105]), .A2(n8692), .B1(
        i_data_bus[41]), .B2(n8684), .ZN(n8325) );
  AOI22D1BWP30P140LVT U8919 ( .A1(i_data_bus[969]), .A2(n8708), .B1(
        i_data_bus[713]), .B2(n8703), .ZN(n8324) );
  AOI22D1BWP30P140LVT U8920 ( .A1(i_data_bus[233]), .A2(n8687), .B1(
        i_data_bus[457]), .B2(n8626), .ZN(n8323) );
  AOI22D1BWP30P140LVT U8921 ( .A1(i_data_bus[873]), .A2(n8706), .B1(
        i_data_bus[649]), .B2(n8693), .ZN(n8308) );
  AOI22D1BWP30P140LVT U8922 ( .A1(i_data_bus[1001]), .A2(n8702), .B1(
        i_data_bus[361]), .B2(n8701), .ZN(n8307) );
  AOI22D1BWP30P140LVT U8923 ( .A1(i_data_bus[745]), .A2(n8696), .B1(
        i_data_bus[297]), .B2(n8705), .ZN(n8306) );
  AOI22D1BWP30P140LVT U8924 ( .A1(i_data_bus[681]), .A2(n8689), .B1(
        i_data_bus[809]), .B2(n8695), .ZN(n8305) );
  ND4D1BWP30P140LVT U8925 ( .A1(n8308), .A2(n8307), .A3(n8306), .A4(n8305), 
        .ZN(n8321) );
  AOI22D1BWP30P140LVT U8926 ( .A1(i_data_bus[9]), .A2(n8683), .B1(
        i_data_bus[329]), .B2(n8685), .ZN(n8312) );
  AOI22D1BWP30P140LVT U8927 ( .A1(i_data_bus[905]), .A2(n8686), .B1(
        i_data_bus[73]), .B2(n8694), .ZN(n8311) );
  AOI22D1BWP30P140LVT U8928 ( .A1(i_data_bus[937]), .A2(n8704), .B1(
        i_data_bus[265]), .B2(n8691), .ZN(n8310) );
  AOI22D1BWP30P140LVT U8929 ( .A1(i_data_bus[777]), .A2(n8707), .B1(
        i_data_bus[841]), .B2(n8690), .ZN(n8309) );
  ND4D1BWP30P140LVT U8930 ( .A1(n8312), .A2(n8311), .A3(n8310), .A4(n8309), 
        .ZN(n8320) );
  INVD1BWP30P140LVT U8931 ( .I(i_data_bus[489]), .ZN(n9690) );
  OAI22D1BWP30P140LVT U8932 ( .A1(n9690), .A2(n8624), .B1(n8313), .B2(n8647), 
        .ZN(n8319) );
  AOI22D1BWP30P140LVT U8933 ( .A1(i_data_bus[201]), .A2(n8713), .B1(
        i_data_bus[425]), .B2(n8717), .ZN(n8317) );
  AOI22D1BWP30P140LVT U8934 ( .A1(i_data_bus[169]), .A2(n8716), .B1(
        i_data_bus[137]), .B2(n8688), .ZN(n8316) );
  AOI22D1BWP30P140LVT U8935 ( .A1(i_data_bus[521]), .A2(n8721), .B1(
        i_data_bus[617]), .B2(n8720), .ZN(n8315) );
  AOI22D1BWP30P140LVT U8936 ( .A1(i_data_bus[585]), .A2(n8722), .B1(
        i_data_bus[553]), .B2(n8723), .ZN(n8314) );
  ND4D1BWP30P140LVT U8937 ( .A1(n8317), .A2(n8316), .A3(n8315), .A4(n8314), 
        .ZN(n8318) );
  NR4D0BWP30P140LVT U8938 ( .A1(n8321), .A2(n8320), .A3(n8319), .A4(n8318), 
        .ZN(n8322) );
  ND4D4BWP30P140LVT U8939 ( .A1(n8325), .A2(n8324), .A3(n8323), .A4(n8322), 
        .ZN(o_data_bus[169]) );
  AOI22D1BWP30P140LVT U8940 ( .A1(i_data_bus[6]), .A2(n8683), .B1(
        i_data_bus[838]), .B2(n8690), .ZN(n8345) );
  AOI22D1BWP30P140LVT U8941 ( .A1(i_data_bus[998]), .A2(n8702), .B1(
        i_data_bus[678]), .B2(n8689), .ZN(n8344) );
  AOI22D1BWP30P140LVT U8942 ( .A1(i_data_bus[230]), .A2(n8687), .B1(
        i_data_bus[422]), .B2(n8717), .ZN(n8343) );
  AOI22D1BWP30P140LVT U8943 ( .A1(i_data_bus[742]), .A2(n8696), .B1(
        i_data_bus[774]), .B2(n8707), .ZN(n8329) );
  AOI22D1BWP30P140LVT U8944 ( .A1(i_data_bus[966]), .A2(n8708), .B1(
        i_data_bus[262]), .B2(n8691), .ZN(n8328) );
  AOI22D1BWP30P140LVT U8945 ( .A1(i_data_bus[102]), .A2(n8692), .B1(
        i_data_bus[806]), .B2(n8695), .ZN(n8327) );
  AOI22D1BWP30P140LVT U8946 ( .A1(i_data_bus[710]), .A2(n8703), .B1(
        i_data_bus[294]), .B2(n8705), .ZN(n8326) );
  ND4D1BWP30P140LVT U8947 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), 
        .ZN(n8341) );
  AOI22D1BWP30P140LVT U8948 ( .A1(i_data_bus[902]), .A2(n8686), .B1(
        i_data_bus[358]), .B2(n8701), .ZN(n8333) );
  AOI22D1BWP30P140LVT U8949 ( .A1(i_data_bus[934]), .A2(n8704), .B1(
        i_data_bus[870]), .B2(n8706), .ZN(n8332) );
  AOI22D1BWP30P140LVT U8950 ( .A1(i_data_bus[38]), .A2(n8684), .B1(
        i_data_bus[70]), .B2(n8694), .ZN(n8331) );
  AOI22D1BWP30P140LVT U8951 ( .A1(i_data_bus[646]), .A2(n8693), .B1(
        i_data_bus[326]), .B2(n8685), .ZN(n8330) );
  ND4D1BWP30P140LVT U8952 ( .A1(n8333), .A2(n8332), .A3(n8331), .A4(n8330), 
        .ZN(n8340) );
  MOAI22D1BWP30P140LVT U8953 ( .A1(n9505), .A2(n8714), .B1(i_data_bus[198]), 
        .B2(n8713), .ZN(n8339) );
  AOI22D1BWP30P140LVT U8954 ( .A1(i_data_bus[486]), .A2(n8718), .B1(
        i_data_bus[390]), .B2(n8719), .ZN(n8337) );
  AOI22D1BWP30P140LVT U8955 ( .A1(i_data_bus[166]), .A2(n8716), .B1(
        i_data_bus[134]), .B2(n8688), .ZN(n8336) );
  AOI22D1BWP30P140LVT U8956 ( .A1(i_data_bus[582]), .A2(n8722), .B1(
        i_data_bus[518]), .B2(n8721), .ZN(n8335) );
  AOI22D1BWP30P140LVT U8957 ( .A1(i_data_bus[614]), .A2(n8720), .B1(
        i_data_bus[550]), .B2(n8723), .ZN(n8334) );
  ND4D1BWP30P140LVT U8958 ( .A1(n8337), .A2(n8336), .A3(n8335), .A4(n8334), 
        .ZN(n8338) );
  NR4D0BWP30P140LVT U8959 ( .A1(n8341), .A2(n8340), .A3(n8339), .A4(n8338), 
        .ZN(n8342) );
  ND4D4BWP30P140LVT U8960 ( .A1(n8345), .A2(n8344), .A3(n8343), .A4(n8342), 
        .ZN(o_data_bus[166]) );
  AOI22D1BWP30P140LVT U8961 ( .A1(i_data_bus[901]), .A2(n8686), .B1(
        i_data_bus[869]), .B2(n8706), .ZN(n8365) );
  AOI22D1BWP30P140LVT U8962 ( .A1(i_data_bus[997]), .A2(n8702), .B1(
        i_data_bus[805]), .B2(n8695), .ZN(n8364) );
  AOI22D1BWP30P140LVT U8963 ( .A1(i_data_bus[165]), .A2(n8716), .B1(
        i_data_bus[485]), .B2(n8718), .ZN(n8363) );
  AOI22D1BWP30P140LVT U8964 ( .A1(i_data_bus[197]), .A2(n8713), .B1(
        i_data_bus[133]), .B2(n8688), .ZN(n8361) );
  AOI22D1BWP30P140LVT U8965 ( .A1(i_data_bus[677]), .A2(n8689), .B1(
        i_data_bus[837]), .B2(n8690), .ZN(n8349) );
  AOI22D1BWP30P140LVT U8966 ( .A1(i_data_bus[933]), .A2(n8704), .B1(
        i_data_bus[69]), .B2(n8694), .ZN(n8348) );
  AOI22D1BWP30P140LVT U8967 ( .A1(i_data_bus[773]), .A2(n8707), .B1(
        i_data_bus[709]), .B2(n8703), .ZN(n8347) );
  AOI22D1BWP30P140LVT U8968 ( .A1(i_data_bus[965]), .A2(n8708), .B1(
        i_data_bus[293]), .B2(n8705), .ZN(n8346) );
  ND4D1BWP30P140LVT U8969 ( .A1(n8349), .A2(n8348), .A3(n8347), .A4(n8346), 
        .ZN(n8360) );
  AOI22D1BWP30P140LVT U8970 ( .A1(i_data_bus[5]), .A2(n8683), .B1(
        i_data_bus[261]), .B2(n8691), .ZN(n8353) );
  AOI22D1BWP30P140LVT U8971 ( .A1(i_data_bus[645]), .A2(n8693), .B1(
        i_data_bus[741]), .B2(n8696), .ZN(n8352) );
  AOI22D1BWP30P140LVT U8972 ( .A1(i_data_bus[101]), .A2(n8692), .B1(
        i_data_bus[357]), .B2(n8701), .ZN(n8351) );
  AOI22D1BWP30P140LVT U8973 ( .A1(i_data_bus[37]), .A2(n8684), .B1(
        i_data_bus[325]), .B2(n8685), .ZN(n8350) );
  ND4D1BWP30P140LVT U8974 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), 
        .ZN(n8359) );
  AOI22D1BWP30P140LVT U8975 ( .A1(i_data_bus[421]), .A2(n8717), .B1(
        i_data_bus[389]), .B2(n8719), .ZN(n8357) );
  AOI22D1BWP30P140LVT U8976 ( .A1(i_data_bus[453]), .A2(n8626), .B1(
        i_data_bus[229]), .B2(n8687), .ZN(n8356) );
  AOI22D1BWP30P140LVT U8977 ( .A1(i_data_bus[517]), .A2(n8721), .B1(
        i_data_bus[549]), .B2(n8723), .ZN(n8355) );
  AOI22D1BWP30P140LVT U8978 ( .A1(i_data_bus[581]), .A2(n8722), .B1(
        i_data_bus[613]), .B2(n8720), .ZN(n8354) );
  ND4D1BWP30P140LVT U8979 ( .A1(n8357), .A2(n8356), .A3(n8355), .A4(n8354), 
        .ZN(n8358) );
  INR4D0BWP30P140LVT U8980 ( .A1(n8361), .B1(n8360), .B2(n8359), .B3(n8358), 
        .ZN(n8362) );
  ND4D4BWP30P140LVT U8981 ( .A1(n8365), .A2(n8364), .A3(n8363), .A4(n8362), 
        .ZN(o_data_bus[165]) );
  AOI22D1BWP30P140LVT U8982 ( .A1(i_data_bus[673]), .A2(n8689), .B1(
        i_data_bus[865]), .B2(n8706), .ZN(n8385) );
  AOI22D1BWP30P140LVT U8983 ( .A1(i_data_bus[289]), .A2(n8705), .B1(
        i_data_bus[321]), .B2(n8685), .ZN(n8384) );
  AOI22D1BWP30P140LVT U8984 ( .A1(i_data_bus[161]), .A2(n8716), .B1(
        i_data_bus[193]), .B2(n8713), .ZN(n8383) );
  AOI22D1BWP30P140LVT U8985 ( .A1(i_data_bus[97]), .A2(n8692), .B1(
        i_data_bus[1]), .B2(n8683), .ZN(n8369) );
  AOI22D1BWP30P140LVT U8986 ( .A1(i_data_bus[897]), .A2(n8686), .B1(
        i_data_bus[641]), .B2(n8693), .ZN(n8368) );
  AOI22D1BWP30P140LVT U8987 ( .A1(i_data_bus[33]), .A2(n8684), .B1(
        i_data_bus[65]), .B2(n8694), .ZN(n8367) );
  AOI22D1BWP30P140LVT U8988 ( .A1(i_data_bus[961]), .A2(n8708), .B1(
        i_data_bus[833]), .B2(n8690), .ZN(n8366) );
  ND4D1BWP30P140LVT U8989 ( .A1(n8369), .A2(n8368), .A3(n8367), .A4(n8366), 
        .ZN(n8381) );
  AOI22D1BWP30P140LVT U8990 ( .A1(i_data_bus[929]), .A2(n8704), .B1(
        i_data_bus[769]), .B2(n8707), .ZN(n8373) );
  AOI22D1BWP30P140LVT U8991 ( .A1(i_data_bus[993]), .A2(n8702), .B1(
        i_data_bus[737]), .B2(n8696), .ZN(n8372) );
  AOI22D1BWP30P140LVT U8992 ( .A1(i_data_bus[705]), .A2(n8703), .B1(
        i_data_bus[353]), .B2(n8701), .ZN(n8371) );
  AOI22D1BWP30P140LVT U8993 ( .A1(i_data_bus[801]), .A2(n8695), .B1(
        i_data_bus[257]), .B2(n8691), .ZN(n8370) );
  ND4D1BWP30P140LVT U8994 ( .A1(n8373), .A2(n8372), .A3(n8371), .A4(n8370), 
        .ZN(n8380) );
  MOAI22D1BWP30P140LVT U8995 ( .A1(n8556), .A2(n8624), .B1(i_data_bus[449]), 
        .B2(n8626), .ZN(n8379) );
  AOI22D1BWP30P140LVT U8996 ( .A1(i_data_bus[417]), .A2(n8717), .B1(
        i_data_bus[129]), .B2(n8688), .ZN(n8377) );
  AOI22D1BWP30P140LVT U8997 ( .A1(i_data_bus[385]), .A2(n8719), .B1(
        i_data_bus[225]), .B2(n8687), .ZN(n8376) );
  AOI22D1BWP30P140LVT U8998 ( .A1(i_data_bus[577]), .A2(n8722), .B1(
        i_data_bus[609]), .B2(n8720), .ZN(n8375) );
  AOI22D1BWP30P140LVT U8999 ( .A1(i_data_bus[545]), .A2(n8723), .B1(
        i_data_bus[513]), .B2(n8721), .ZN(n8374) );
  ND4D1BWP30P140LVT U9000 ( .A1(n8377), .A2(n8376), .A3(n8375), .A4(n8374), 
        .ZN(n8378) );
  NR4D0BWP30P140LVT U9001 ( .A1(n8381), .A2(n8380), .A3(n8379), .A4(n8378), 
        .ZN(n8382) );
  ND4D4BWP30P140LVT U9002 ( .A1(n8385), .A2(n8384), .A3(n8383), .A4(n8382), 
        .ZN(o_data_bus[161]) );
  AOI22D1BWP30P140LVT U9003 ( .A1(i_data_bus[66]), .A2(n9549), .B1(
        i_data_bus[34]), .B2(n9548), .ZN(n8407) );
  AOI22D1BWP30P140LVT U9004 ( .A1(i_data_bus[770]), .A2(n9547), .B1(
        i_data_bus[706]), .B2(n9554), .ZN(n8406) );
  AOI22D1BWP30P140LVT U9005 ( .A1(i_data_bus[386]), .A2(n9585), .B1(
        i_data_bus[130]), .B2(n9533), .ZN(n8405) );
  AOI22D1BWP30P140LVT U9006 ( .A1(i_data_bus[802]), .A2(n9552), .B1(
        i_data_bus[738]), .B2(n9546), .ZN(n8389) );
  AOI22D1BWP30P140LVT U9007 ( .A1(i_data_bus[98]), .A2(n9555), .B1(
        i_data_bus[642]), .B2(n9558), .ZN(n8388) );
  AOI22D1BWP30P140LVT U9008 ( .A1(i_data_bus[2]), .A2(n9553), .B1(
        i_data_bus[834]), .B2(n9557), .ZN(n8387) );
  AOI22D1BWP30P140LVT U9009 ( .A1(i_data_bus[866]), .A2(n9556), .B1(
        i_data_bus[674]), .B2(n9559), .ZN(n8386) );
  ND4D1BWP30P140LVT U9010 ( .A1(n8389), .A2(n8388), .A3(n8387), .A4(n8386), 
        .ZN(n8403) );
  INVD1BWP30P140LVT U9011 ( .I(n9550), .ZN(n9483) );
  OAI22D1BWP30P140LVT U9012 ( .A1(n8391), .A2(n9483), .B1(n9139), .B2(n8390), 
        .ZN(n8402) );
  AOI22D1BWP30P140LVT U9013 ( .A1(i_data_bus[962]), .A2(n9551), .B1(
        i_data_bus[322]), .B2(n9570), .ZN(n8395) );
  AOI22D1BWP30P140LVT U9014 ( .A1(i_data_bus[290]), .A2(n9584), .B1(
        i_data_bus[482]), .B2(n9580), .ZN(n8394) );
  AOI22D1BWP30P140LVT U9015 ( .A1(i_data_bus[578]), .A2(n9572), .B1(
        i_data_bus[610]), .B2(n9574), .ZN(n8393) );
  AOI22D1BWP30P140LVT U9016 ( .A1(i_data_bus[546]), .A2(n9575), .B1(
        i_data_bus[514]), .B2(n9573), .ZN(n8392) );
  ND4D1BWP30P140LVT U9017 ( .A1(n8395), .A2(n8394), .A3(n8393), .A4(n8392), 
        .ZN(n8401) );
  AOI22D1BWP30P140LVT U9018 ( .A1(i_data_bus[930]), .A2(n9587), .B1(
        i_data_bus[418]), .B2(n9532), .ZN(n8399) );
  AOI22D1BWP30P140LVT U9019 ( .A1(i_data_bus[898]), .A2(n9581), .B1(
        i_data_bus[450]), .B2(n9582), .ZN(n8398) );
  AOI22D1BWP30P140LVT U9020 ( .A1(i_data_bus[994]), .A2(n9571), .B1(
        i_data_bus[354]), .B2(n9569), .ZN(n8397) );
  AOI22D1BWP30P140LVT U9021 ( .A1(i_data_bus[162]), .A2(n9583), .B1(
        i_data_bus[226]), .B2(n9568), .ZN(n8396) );
  ND4D1BWP30P140LVT U9022 ( .A1(n8399), .A2(n8398), .A3(n8397), .A4(n8396), 
        .ZN(n8400) );
  NR4D0BWP30P140LVT U9023 ( .A1(n8403), .A2(n8402), .A3(n8401), .A4(n8400), 
        .ZN(n8404) );
  ND4D4BWP30P140LVT U9024 ( .A1(n8407), .A2(n8406), .A3(n8405), .A4(n8404), 
        .ZN(o_data_bus[226]) );
  AOI22D1BWP30P140LVT U9025 ( .A1(i_data_bus[53]), .A2(n9670), .B1(
        i_data_bus[181]), .B2(n9675), .ZN(n8428) );
  AOI22D1BWP30P140LVT U9026 ( .A1(i_data_bus[117]), .A2(n9680), .B1(
        i_data_bus[21]), .B2(n9676), .ZN(n8427) );
  AOI22D1BWP30P140LVT U9027 ( .A1(i_data_bus[757]), .A2(n9706), .B1(
        i_data_bus[501]), .B2(n9656), .ZN(n8426) );
  AOI22D1BWP30P140LVT U9028 ( .A1(i_data_bus[85]), .A2(n9672), .B1(
        i_data_bus[149]), .B2(n9681), .ZN(n8411) );
  AOI22D1BWP30P140LVT U9029 ( .A1(i_data_bus[213]), .A2(n9679), .B1(
        i_data_bus[245]), .B2(n9671), .ZN(n8410) );
  AOI22D1BWP30P140LVT U9030 ( .A1(i_data_bus[917]), .A2(n9682), .B1(
        i_data_bus[1013]), .B2(n9677), .ZN(n8409) );
  AOI22D1BWP30P140LVT U9031 ( .A1(i_data_bus[949]), .A2(n9669), .B1(
        i_data_bus[981]), .B2(n9678), .ZN(n8408) );
  ND4D1BWP30P140LVT U9032 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), 
        .ZN(n8424) );
  MOAI22D1BWP30P140LVT U9033 ( .A1(n8412), .A2(n9687), .B1(i_data_bus[725]), 
        .B2(n9704), .ZN(n8423) );
  AOI22D1BWP30P140LVT U9034 ( .A1(i_data_bus[341]), .A2(n9692), .B1(
        i_data_bus[277]), .B2(n9694), .ZN(n8416) );
  AOI22D1BWP30P140LVT U9035 ( .A1(i_data_bus[853]), .A2(n9693), .B1(
        i_data_bus[405]), .B2(n9708), .ZN(n8415) );
  AOI22D1BWP30P140LVT U9036 ( .A1(i_data_bus[597]), .A2(n9697), .B1(
        i_data_bus[565]), .B2(n9695), .ZN(n8414) );
  AOI22D1BWP30P140LVT U9037 ( .A1(i_data_bus[629]), .A2(n9696), .B1(
        i_data_bus[533]), .B2(n9698), .ZN(n8413) );
  ND4D1BWP30P140LVT U9038 ( .A1(n8416), .A2(n8415), .A3(n8414), .A4(n8413), 
        .ZN(n8422) );
  AOI22D1BWP30P140LVT U9039 ( .A1(i_data_bus[789]), .A2(n9673), .B1(
        i_data_bus[373]), .B2(n9691), .ZN(n8420) );
  AOI22D1BWP30P140LVT U9040 ( .A1(i_data_bus[821]), .A2(n9674), .B1(
        i_data_bus[437]), .B2(n9709), .ZN(n8419) );
  AOI22D1BWP30P140LVT U9041 ( .A1(i_data_bus[661]), .A2(n9707), .B1(
        i_data_bus[885]), .B2(n9710), .ZN(n8418) );
  AOI22D1BWP30P140LVT U9042 ( .A1(i_data_bus[693]), .A2(n9705), .B1(
        i_data_bus[469]), .B2(n9703), .ZN(n8417) );
  ND4D1BWP30P140LVT U9043 ( .A1(n8420), .A2(n8419), .A3(n8418), .A4(n8417), 
        .ZN(n8421) );
  NR4D0BWP30P140LVT U9044 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), 
        .ZN(n8425) );
  ND4D4BWP30P140LVT U9045 ( .A1(n8428), .A2(n8427), .A3(n8426), .A4(n8425), 
        .ZN(o_data_bus[21]) );
  AOI22D1BWP30P140LVT U9046 ( .A1(i_data_bus[947]), .A2(n9669), .B1(
        i_data_bus[915]), .B2(n9682), .ZN(n8449) );
  AOI22D1BWP30P140LVT U9047 ( .A1(i_data_bus[51]), .A2(n9670), .B1(
        i_data_bus[243]), .B2(n9671), .ZN(n8448) );
  AOI22D1BWP30P140LVT U9048 ( .A1(i_data_bus[275]), .A2(n9694), .B1(
        i_data_bus[467]), .B2(n9703), .ZN(n8447) );
  AOI22D1BWP30P140LVT U9049 ( .A1(i_data_bus[115]), .A2(n9680), .B1(
        i_data_bus[83]), .B2(n9672), .ZN(n8432) );
  AOI22D1BWP30P140LVT U9050 ( .A1(i_data_bus[1011]), .A2(n9677), .B1(
        i_data_bus[19]), .B2(n9676), .ZN(n8431) );
  AOI22D1BWP30P140LVT U9051 ( .A1(i_data_bus[979]), .A2(n9678), .B1(
        i_data_bus[211]), .B2(n9679), .ZN(n8430) );
  AOI22D1BWP30P140LVT U9052 ( .A1(i_data_bus[179]), .A2(n9675), .B1(
        i_data_bus[147]), .B2(n9681), .ZN(n8429) );
  ND4D1BWP30P140LVT U9053 ( .A1(n8432), .A2(n8431), .A3(n8430), .A4(n8429), 
        .ZN(n8445) );
  MOAI22D1BWP30P140LVT U9054 ( .A1(n8433), .A2(n9687), .B1(i_data_bus[371]), 
        .B2(n9691), .ZN(n8444) );
  AOI22D1BWP30P140LVT U9055 ( .A1(i_data_bus[403]), .A2(n9708), .B1(
        i_data_bus[691]), .B2(n9705), .ZN(n8437) );
  AOI22D1BWP30P140LVT U9056 ( .A1(i_data_bus[819]), .A2(n9674), .B1(
        i_data_bus[723]), .B2(n9704), .ZN(n8436) );
  AOI22D1BWP30P140LVT U9057 ( .A1(i_data_bus[563]), .A2(n9695), .B1(
        i_data_bus[627]), .B2(n9696), .ZN(n8435) );
  AOI22D1BWP30P140LVT U9058 ( .A1(i_data_bus[531]), .A2(n9698), .B1(
        i_data_bus[595]), .B2(n9697), .ZN(n8434) );
  ND4D1BWP30P140LVT U9059 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), 
        .ZN(n8443) );
  AOI22D1BWP30P140LVT U9060 ( .A1(i_data_bus[787]), .A2(n9673), .B1(
        i_data_bus[883]), .B2(n9710), .ZN(n8441) );
  AOI22D1BWP30P140LVT U9061 ( .A1(i_data_bus[755]), .A2(n9706), .B1(
        i_data_bus[659]), .B2(n9707), .ZN(n8440) );
  AOI22D1BWP30P140LVT U9062 ( .A1(i_data_bus[851]), .A2(n9693), .B1(
        i_data_bus[435]), .B2(n9709), .ZN(n8439) );
  AOI22D1BWP30P140LVT U9063 ( .A1(i_data_bus[339]), .A2(n9692), .B1(
        i_data_bus[499]), .B2(n9656), .ZN(n8438) );
  ND4D1BWP30P140LVT U9064 ( .A1(n8441), .A2(n8440), .A3(n8439), .A4(n8438), 
        .ZN(n8442) );
  NR4D0BWP30P140LVT U9065 ( .A1(n8445), .A2(n8444), .A3(n8443), .A4(n8442), 
        .ZN(n8446) );
  ND4D4BWP30P140LVT U9066 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8446), 
        .ZN(o_data_bus[19]) );
  AOI22D1BWP30P140LVT U9067 ( .A1(i_data_bus[82]), .A2(n9672), .B1(
        i_data_bus[914]), .B2(n9682), .ZN(n8469) );
  AOI22D1BWP30P140LVT U9068 ( .A1(i_data_bus[946]), .A2(n9669), .B1(
        i_data_bus[210]), .B2(n9679), .ZN(n8468) );
  AOI22D1BWP30P140LVT U9069 ( .A1(i_data_bus[370]), .A2(n9691), .B1(
        i_data_bus[306]), .B2(n9655), .ZN(n8467) );
  AOI22D1BWP30P140LVT U9070 ( .A1(i_data_bus[882]), .A2(n9710), .B1(
        i_data_bus[722]), .B2(n9704), .ZN(n8465) );
  AOI22D1BWP30P140LVT U9071 ( .A1(i_data_bus[978]), .A2(n9678), .B1(
        i_data_bus[114]), .B2(n9680), .ZN(n8453) );
  AOI22D1BWP30P140LVT U9072 ( .A1(i_data_bus[1010]), .A2(n9677), .B1(
        i_data_bus[146]), .B2(n9681), .ZN(n8452) );
  AOI22D1BWP30P140LVT U9073 ( .A1(i_data_bus[50]), .A2(n9670), .B1(
        i_data_bus[18]), .B2(n9676), .ZN(n8451) );
  AOI22D1BWP30P140LVT U9074 ( .A1(i_data_bus[242]), .A2(n9671), .B1(
        i_data_bus[178]), .B2(n9675), .ZN(n8450) );
  ND4D1BWP30P140LVT U9075 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), 
        .ZN(n8464) );
  AOI22D1BWP30P140LVT U9076 ( .A1(i_data_bus[818]), .A2(n9674), .B1(
        i_data_bus[498]), .B2(n9656), .ZN(n8457) );
  AOI22D1BWP30P140LVT U9077 ( .A1(i_data_bus[690]), .A2(n9705), .B1(
        i_data_bus[274]), .B2(n9694), .ZN(n8456) );
  AOI22D1BWP30P140LVT U9078 ( .A1(i_data_bus[530]), .A2(n9698), .B1(
        i_data_bus[562]), .B2(n9695), .ZN(n8455) );
  AOI22D1BWP30P140LVT U9079 ( .A1(i_data_bus[626]), .A2(n9696), .B1(
        i_data_bus[594]), .B2(n9697), .ZN(n8454) );
  ND4D1BWP30P140LVT U9080 ( .A1(n8457), .A2(n8456), .A3(n8455), .A4(n8454), 
        .ZN(n8463) );
  AOI22D1BWP30P140LVT U9081 ( .A1(i_data_bus[466]), .A2(n9703), .B1(
        i_data_bus[754]), .B2(n9706), .ZN(n8461) );
  AOI22D1BWP30P140LVT U9082 ( .A1(i_data_bus[402]), .A2(n9708), .B1(
        i_data_bus[850]), .B2(n9693), .ZN(n8460) );
  AOI22D1BWP30P140LVT U9083 ( .A1(i_data_bus[658]), .A2(n9707), .B1(
        i_data_bus[786]), .B2(n9673), .ZN(n8459) );
  AOI22D1BWP30P140LVT U9084 ( .A1(i_data_bus[434]), .A2(n9709), .B1(
        i_data_bus[338]), .B2(n9692), .ZN(n8458) );
  ND4D1BWP30P140LVT U9085 ( .A1(n8461), .A2(n8460), .A3(n8459), .A4(n8458), 
        .ZN(n8462) );
  INR4D0BWP30P140LVT U9086 ( .A1(n8465), .B1(n8464), .B2(n8463), .B3(n8462), 
        .ZN(n8466) );
  ND4D4BWP30P140LVT U9087 ( .A1(n8469), .A2(n8468), .A3(n8467), .A4(n8466), 
        .ZN(o_data_bus[18]) );
  AOI22D1BWP30P140LVT U9088 ( .A1(i_data_bus[913]), .A2(n9682), .B1(
        i_data_bus[145]), .B2(n9681), .ZN(n8489) );
  AOI22D1BWP30P140LVT U9089 ( .A1(i_data_bus[1009]), .A2(n9677), .B1(
        i_data_bus[209]), .B2(n9679), .ZN(n8488) );
  AOI22D1BWP30P140LVT U9090 ( .A1(i_data_bus[721]), .A2(n9704), .B1(
        i_data_bus[273]), .B2(n9694), .ZN(n8487) );
  AOI22D1BWP30P140LVT U9091 ( .A1(i_data_bus[689]), .A2(n9705), .B1(
        i_data_bus[465]), .B2(n9703), .ZN(n8485) );
  AOI22D1BWP30P140LVT U9092 ( .A1(i_data_bus[17]), .A2(n9676), .B1(
        i_data_bus[177]), .B2(n9675), .ZN(n8473) );
  AOI22D1BWP30P140LVT U9093 ( .A1(i_data_bus[49]), .A2(n9670), .B1(
        i_data_bus[945]), .B2(n9669), .ZN(n8472) );
  AOI22D1BWP30P140LVT U9094 ( .A1(i_data_bus[977]), .A2(n9678), .B1(
        i_data_bus[241]), .B2(n9671), .ZN(n8471) );
  AOI22D1BWP30P140LVT U9095 ( .A1(i_data_bus[81]), .A2(n9672), .B1(
        i_data_bus[113]), .B2(n9680), .ZN(n8470) );
  ND4D1BWP30P140LVT U9096 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), 
        .ZN(n8484) );
  AOI22D1BWP30P140LVT U9097 ( .A1(i_data_bus[753]), .A2(n9706), .B1(
        i_data_bus[497]), .B2(n9656), .ZN(n8477) );
  AOI22D1BWP30P140LVT U9098 ( .A1(i_data_bus[433]), .A2(n9709), .B1(
        i_data_bus[401]), .B2(n9708), .ZN(n8476) );
  AOI22D1BWP30P140LVT U9099 ( .A1(i_data_bus[625]), .A2(n9696), .B1(
        i_data_bus[561]), .B2(n9695), .ZN(n8475) );
  AOI22D1BWP30P140LVT U9100 ( .A1(i_data_bus[593]), .A2(n9697), .B1(
        i_data_bus[529]), .B2(n9698), .ZN(n8474) );
  ND4D1BWP30P140LVT U9101 ( .A1(n8477), .A2(n8476), .A3(n8475), .A4(n8474), 
        .ZN(n8483) );
  AOI22D1BWP30P140LVT U9102 ( .A1(i_data_bus[305]), .A2(n9655), .B1(
        i_data_bus[369]), .B2(n9691), .ZN(n8481) );
  AOI22D1BWP30P140LVT U9103 ( .A1(i_data_bus[337]), .A2(n9692), .B1(
        i_data_bus[785]), .B2(n9673), .ZN(n8480) );
  AOI22D1BWP30P140LVT U9104 ( .A1(i_data_bus[849]), .A2(n9693), .B1(
        i_data_bus[817]), .B2(n9674), .ZN(n8479) );
  AOI22D1BWP30P140LVT U9105 ( .A1(i_data_bus[881]), .A2(n9710), .B1(
        i_data_bus[657]), .B2(n9707), .ZN(n8478) );
  ND4D1BWP30P140LVT U9106 ( .A1(n8481), .A2(n8480), .A3(n8479), .A4(n8478), 
        .ZN(n8482) );
  INR4D0BWP30P140LVT U9107 ( .A1(n8485), .B1(n8484), .B2(n8483), .B3(n8482), 
        .ZN(n8486) );
  ND4D4BWP30P140LVT U9108 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), 
        .ZN(o_data_bus[17]) );
  AOI22D1BWP30P140LVT U9109 ( .A1(i_data_bus[904]), .A2(n9682), .B1(
        i_data_bus[232]), .B2(n9671), .ZN(n8509) );
  AOI22D1BWP30P140LVT U9110 ( .A1(i_data_bus[936]), .A2(n9669), .B1(
        i_data_bus[40]), .B2(n9670), .ZN(n8508) );
  AOI22D1BWP30P140LVT U9111 ( .A1(i_data_bus[680]), .A2(n9705), .B1(
        i_data_bus[488]), .B2(n9656), .ZN(n8507) );
  AOI22D1BWP30P140LVT U9112 ( .A1(i_data_bus[72]), .A2(n9672), .B1(
        i_data_bus[200]), .B2(n9679), .ZN(n8493) );
  AOI22D1BWP30P140LVT U9113 ( .A1(i_data_bus[168]), .A2(n9675), .B1(
        i_data_bus[136]), .B2(n9681), .ZN(n8492) );
  AOI22D1BWP30P140LVT U9114 ( .A1(i_data_bus[8]), .A2(n9676), .B1(
        i_data_bus[1000]), .B2(n9677), .ZN(n8491) );
  AOI22D1BWP30P140LVT U9115 ( .A1(i_data_bus[968]), .A2(n9678), .B1(
        i_data_bus[104]), .B2(n9680), .ZN(n8490) );
  ND4D1BWP30P140LVT U9116 ( .A1(n8493), .A2(n8492), .A3(n8491), .A4(n8490), 
        .ZN(n8505) );
  MOAI22D1BWP30P140LVT U9117 ( .A1(n9462), .A2(n9687), .B1(i_data_bus[712]), 
        .B2(n9704), .ZN(n8504) );
  AOI22D1BWP30P140LVT U9118 ( .A1(i_data_bus[456]), .A2(n9703), .B1(
        i_data_bus[360]), .B2(n9691), .ZN(n8497) );
  AOI22D1BWP30P140LVT U9119 ( .A1(i_data_bus[424]), .A2(n9709), .B1(
        i_data_bus[648]), .B2(n9707), .ZN(n8496) );
  AOI22D1BWP30P140LVT U9120 ( .A1(i_data_bus[552]), .A2(n9695), .B1(
        i_data_bus[520]), .B2(n9698), .ZN(n8495) );
  AOI22D1BWP30P140LVT U9121 ( .A1(i_data_bus[616]), .A2(n9696), .B1(
        i_data_bus[584]), .B2(n9697), .ZN(n8494) );
  ND4D1BWP30P140LVT U9122 ( .A1(n8497), .A2(n8496), .A3(n8495), .A4(n8494), 
        .ZN(n8503) );
  AOI22D1BWP30P140LVT U9123 ( .A1(i_data_bus[328]), .A2(n9692), .B1(
        i_data_bus[776]), .B2(n9673), .ZN(n8501) );
  AOI22D1BWP30P140LVT U9124 ( .A1(i_data_bus[264]), .A2(n9694), .B1(
        i_data_bus[808]), .B2(n9674), .ZN(n8500) );
  AOI22D1BWP30P140LVT U9125 ( .A1(i_data_bus[840]), .A2(n9693), .B1(
        i_data_bus[872]), .B2(n9710), .ZN(n8499) );
  AOI22D1BWP30P140LVT U9126 ( .A1(i_data_bus[744]), .A2(n9706), .B1(
        i_data_bus[392]), .B2(n9708), .ZN(n8498) );
  ND4D1BWP30P140LVT U9127 ( .A1(n8501), .A2(n8500), .A3(n8499), .A4(n8498), 
        .ZN(n8502) );
  NR4D0BWP30P140LVT U9128 ( .A1(n8505), .A2(n8504), .A3(n8503), .A4(n8502), 
        .ZN(n8506) );
  ND4D4BWP30P140LVT U9129 ( .A1(n8509), .A2(n8508), .A3(n8507), .A4(n8506), 
        .ZN(o_data_bus[8]) );
  AOI22D1BWP30P140LVT U9130 ( .A1(i_data_bus[651]), .A2(n9558), .B1(
        i_data_bus[715]), .B2(n9554), .ZN(n8530) );
  AOI22D1BWP30P140LVT U9131 ( .A1(i_data_bus[107]), .A2(n9555), .B1(
        i_data_bus[683]), .B2(n9559), .ZN(n8529) );
  AOI22D1BWP30P140LVT U9132 ( .A1(i_data_bus[907]), .A2(n9581), .B1(
        i_data_bus[203]), .B2(n9550), .ZN(n8528) );
  AOI22D1BWP30P140LVT U9133 ( .A1(i_data_bus[843]), .A2(n9557), .B1(
        i_data_bus[811]), .B2(n9552), .ZN(n8513) );
  AOI22D1BWP30P140LVT U9134 ( .A1(i_data_bus[43]), .A2(n9548), .B1(
        i_data_bus[779]), .B2(n9547), .ZN(n8512) );
  AOI22D1BWP30P140LVT U9135 ( .A1(i_data_bus[11]), .A2(n9553), .B1(
        i_data_bus[875]), .B2(n9556), .ZN(n8511) );
  AOI22D1BWP30P140LVT U9136 ( .A1(i_data_bus[75]), .A2(n9549), .B1(
        i_data_bus[747]), .B2(n9546), .ZN(n8510) );
  ND4D1BWP30P140LVT U9137 ( .A1(n8513), .A2(n8512), .A3(n8511), .A4(n8510), 
        .ZN(n8526) );
  OAI22D1BWP30P140LVT U9138 ( .A1(n9650), .A2(n9526), .B1(n8514), .B2(n9247), 
        .ZN(n8525) );
  AOI22D1BWP30P140LVT U9139 ( .A1(i_data_bus[1003]), .A2(n9571), .B1(
        i_data_bus[139]), .B2(n9533), .ZN(n8518) );
  AOI22D1BWP30P140LVT U9140 ( .A1(i_data_bus[491]), .A2(n9580), .B1(
        i_data_bus[235]), .B2(n9568), .ZN(n8517) );
  AOI22D1BWP30P140LVT U9141 ( .A1(i_data_bus[619]), .A2(n9574), .B1(
        i_data_bus[555]), .B2(n9575), .ZN(n8516) );
  AOI22D1BWP30P140LVT U9142 ( .A1(i_data_bus[523]), .A2(n9573), .B1(
        i_data_bus[587]), .B2(n9572), .ZN(n8515) );
  ND4D1BWP30P140LVT U9143 ( .A1(n8518), .A2(n8517), .A3(n8516), .A4(n8515), 
        .ZN(n8524) );
  AOI22D1BWP30P140LVT U9144 ( .A1(i_data_bus[939]), .A2(n9587), .B1(
        i_data_bus[395]), .B2(n9585), .ZN(n8522) );
  AOI22D1BWP30P140LVT U9145 ( .A1(i_data_bus[971]), .A2(n9551), .B1(
        i_data_bus[363]), .B2(n9569), .ZN(n8521) );
  AOI22D1BWP30P140LVT U9146 ( .A1(i_data_bus[427]), .A2(n9532), .B1(
        i_data_bus[299]), .B2(n9584), .ZN(n8520) );
  AOI22D1BWP30P140LVT U9147 ( .A1(i_data_bus[171]), .A2(n9583), .B1(
        i_data_bus[267]), .B2(n9586), .ZN(n8519) );
  ND4D1BWP30P140LVT U9148 ( .A1(n8522), .A2(n8521), .A3(n8520), .A4(n8519), 
        .ZN(n8523) );
  NR4D0BWP30P140LVT U9149 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), 
        .ZN(n8527) );
  ND4D4BWP30P140LVT U9150 ( .A1(n8530), .A2(n8529), .A3(n8528), .A4(n8527), 
        .ZN(o_data_bus[235]) );
  AOI22D1BWP30P140LVT U9151 ( .A1(i_data_bus[810]), .A2(n9552), .B1(
        i_data_bus[682]), .B2(n9559), .ZN(n8551) );
  AOI22D1BWP30P140LVT U9152 ( .A1(i_data_bus[10]), .A2(n9553), .B1(
        i_data_bus[874]), .B2(n9556), .ZN(n8550) );
  AOI22D1BWP30P140LVT U9153 ( .A1(i_data_bus[266]), .A2(n9586), .B1(
        i_data_bus[138]), .B2(n9533), .ZN(n8549) );
  AOI22D1BWP30P140LVT U9154 ( .A1(i_data_bus[106]), .A2(n9555), .B1(
        i_data_bus[842]), .B2(n9557), .ZN(n8534) );
  AOI22D1BWP30P140LVT U9155 ( .A1(i_data_bus[650]), .A2(n9558), .B1(
        i_data_bus[746]), .B2(n9546), .ZN(n8533) );
  AOI22D1BWP30P140LVT U9156 ( .A1(i_data_bus[778]), .A2(n9547), .B1(
        i_data_bus[714]), .B2(n9554), .ZN(n8532) );
  AOI22D1BWP30P140LVT U9157 ( .A1(i_data_bus[42]), .A2(n9548), .B1(
        i_data_bus[74]), .B2(n9549), .ZN(n8531) );
  ND4D1BWP30P140LVT U9158 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), 
        .ZN(n8547) );
  OAI22D1BWP30P140LVT U9159 ( .A1(n8887), .A2(n9397), .B1(n8535), .B2(n9245), 
        .ZN(n8546) );
  AOI22D1BWP30P140LVT U9160 ( .A1(i_data_bus[234]), .A2(n9568), .B1(
        i_data_bus[458]), .B2(n9582), .ZN(n8539) );
  AOI22D1BWP30P140LVT U9161 ( .A1(i_data_bus[1002]), .A2(n9571), .B1(
        i_data_bus[330]), .B2(n9570), .ZN(n8538) );
  AOI22D1BWP30P140LVT U9162 ( .A1(i_data_bus[618]), .A2(n9574), .B1(
        i_data_bus[586]), .B2(n9572), .ZN(n8537) );
  AOI22D1BWP30P140LVT U9163 ( .A1(i_data_bus[554]), .A2(n9575), .B1(
        i_data_bus[522]), .B2(n9573), .ZN(n8536) );
  ND4D1BWP30P140LVT U9164 ( .A1(n8539), .A2(n8538), .A3(n8537), .A4(n8536), 
        .ZN(n8545) );
  AOI22D1BWP30P140LVT U9165 ( .A1(i_data_bus[938]), .A2(n9587), .B1(
        i_data_bus[298]), .B2(n9584), .ZN(n8543) );
  AOI22D1BWP30P140LVT U9166 ( .A1(i_data_bus[906]), .A2(n9581), .B1(
        i_data_bus[202]), .B2(n9550), .ZN(n8542) );
  AOI22D1BWP30P140LVT U9167 ( .A1(i_data_bus[170]), .A2(n9583), .B1(
        i_data_bus[426]), .B2(n9532), .ZN(n8541) );
  AOI22D1BWP30P140LVT U9168 ( .A1(i_data_bus[970]), .A2(n9551), .B1(
        i_data_bus[362]), .B2(n9569), .ZN(n8540) );
  ND4D1BWP30P140LVT U9169 ( .A1(n8543), .A2(n8542), .A3(n8541), .A4(n8540), 
        .ZN(n8544) );
  NR4D0BWP30P140LVT U9170 ( .A1(n8547), .A2(n8546), .A3(n8545), .A4(n8544), 
        .ZN(n8548) );
  ND4D4BWP30P140LVT U9171 ( .A1(n8551), .A2(n8550), .A3(n8549), .A4(n8548), 
        .ZN(o_data_bus[234]) );
  AOI22D1BWP30P140LVT U9172 ( .A1(i_data_bus[865]), .A2(n9556), .B1(
        i_data_bus[833]), .B2(n9557), .ZN(n8572) );
  AOI22D1BWP30P140LVT U9173 ( .A1(i_data_bus[1]), .A2(n9553), .B1(
        i_data_bus[641]), .B2(n9558), .ZN(n8571) );
  AOI22D1BWP30P140LVT U9174 ( .A1(i_data_bus[897]), .A2(n9581), .B1(
        i_data_bus[321]), .B2(n9570), .ZN(n8570) );
  AOI22D1BWP30P140LVT U9175 ( .A1(i_data_bus[33]), .A2(n9548), .B1(
        i_data_bus[705]), .B2(n9554), .ZN(n8555) );
  AOI22D1BWP30P140LVT U9176 ( .A1(i_data_bus[97]), .A2(n9555), .B1(
        i_data_bus[673]), .B2(n9559), .ZN(n8554) );
  AOI22D1BWP30P140LVT U9177 ( .A1(i_data_bus[65]), .A2(n9549), .B1(
        i_data_bus[769]), .B2(n9547), .ZN(n8553) );
  AOI22D1BWP30P140LVT U9178 ( .A1(i_data_bus[801]), .A2(n9552), .B1(
        i_data_bus[737]), .B2(n9546), .ZN(n8552) );
  ND4D1BWP30P140LVT U9179 ( .A1(n8555), .A2(n8554), .A3(n8553), .A4(n8552), 
        .ZN(n8568) );
  MOAI22D1BWP30P140LVT U9180 ( .A1(n8556), .A2(n9397), .B1(i_data_bus[193]), 
        .B2(n9550), .ZN(n8567) );
  AOI22D1BWP30P140LVT U9181 ( .A1(i_data_bus[961]), .A2(n9551), .B1(
        i_data_bus[385]), .B2(n9585), .ZN(n8560) );
  AOI22D1BWP30P140LVT U9182 ( .A1(i_data_bus[353]), .A2(n9569), .B1(
        i_data_bus[289]), .B2(n9584), .ZN(n8559) );
  AOI22D1BWP30P140LVT U9183 ( .A1(i_data_bus[545]), .A2(n9575), .B1(
        i_data_bus[513]), .B2(n9573), .ZN(n8558) );
  AOI22D1BWP30P140LVT U9184 ( .A1(i_data_bus[577]), .A2(n9572), .B1(
        i_data_bus[609]), .B2(n9574), .ZN(n8557) );
  ND4D1BWP30P140LVT U9185 ( .A1(n8560), .A2(n8559), .A3(n8558), .A4(n8557), 
        .ZN(n8566) );
  AOI22D1BWP30P140LVT U9186 ( .A1(i_data_bus[993]), .A2(n9571), .B1(
        i_data_bus[225]), .B2(n9568), .ZN(n8564) );
  AOI22D1BWP30P140LVT U9187 ( .A1(i_data_bus[161]), .A2(n9583), .B1(
        i_data_bus[417]), .B2(n9532), .ZN(n8563) );
  AOI22D1BWP30P140LVT U9188 ( .A1(i_data_bus[929]), .A2(n9587), .B1(
        i_data_bus[449]), .B2(n9582), .ZN(n8562) );
  AOI22D1BWP30P140LVT U9189 ( .A1(i_data_bus[257]), .A2(n9586), .B1(
        i_data_bus[129]), .B2(n9533), .ZN(n8561) );
  ND4D1BWP30P140LVT U9190 ( .A1(n8564), .A2(n8563), .A3(n8562), .A4(n8561), 
        .ZN(n8565) );
  NR4D0BWP30P140LVT U9191 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), 
        .ZN(n8569) );
  ND4D4BWP30P140LVT U9192 ( .A1(n8572), .A2(n8571), .A3(n8570), .A4(n8569), 
        .ZN(o_data_bus[225]) );
  AOI22D1BWP30P140LVT U9193 ( .A1(i_data_bus[953]), .A2(n8704), .B1(
        i_data_bus[729]), .B2(n8703), .ZN(n8593) );
  AOI22D1BWP30P140LVT U9194 ( .A1(i_data_bus[121]), .A2(n8692), .B1(
        i_data_bus[889]), .B2(n8706), .ZN(n8592) );
  AOI22D1BWP30P140LVT U9195 ( .A1(i_data_bus[153]), .A2(n8688), .B1(
        i_data_bus[217]), .B2(n8713), .ZN(n8591) );
  AOI22D1BWP30P140LVT U9196 ( .A1(i_data_bus[665]), .A2(n8693), .B1(
        i_data_bus[377]), .B2(n8701), .ZN(n8576) );
  AOI22D1BWP30P140LVT U9197 ( .A1(i_data_bus[825]), .A2(n8695), .B1(
        i_data_bus[697]), .B2(n8689), .ZN(n8575) );
  AOI22D1BWP30P140LVT U9198 ( .A1(i_data_bus[313]), .A2(n8705), .B1(
        i_data_bus[857]), .B2(n8690), .ZN(n8574) );
  AOI22D1BWP30P140LVT U9199 ( .A1(i_data_bus[921]), .A2(n8686), .B1(
        i_data_bus[793]), .B2(n8707), .ZN(n8573) );
  ND4D1BWP30P140LVT U9200 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), 
        .ZN(n8589) );
  AOI22D1BWP30P140LVT U9201 ( .A1(i_data_bus[1017]), .A2(n8702), .B1(
        i_data_bus[985]), .B2(n8708), .ZN(n8580) );
  AOI22D1BWP30P140LVT U9202 ( .A1(i_data_bus[89]), .A2(n8694), .B1(
        i_data_bus[281]), .B2(n8691), .ZN(n8579) );
  AOI22D1BWP30P140LVT U9203 ( .A1(i_data_bus[25]), .A2(n8683), .B1(
        i_data_bus[345]), .B2(n8685), .ZN(n8578) );
  AOI22D1BWP30P140LVT U9204 ( .A1(i_data_bus[57]), .A2(n8684), .B1(
        i_data_bus[761]), .B2(n8696), .ZN(n8577) );
  ND4D1BWP30P140LVT U9205 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n8577), 
        .ZN(n8588) );
  OAI22D1BWP30P140LVT U9206 ( .A1(n8581), .A2(n8647), .B1(n8761), .B2(n8624), 
        .ZN(n8587) );
  AOI22D1BWP30P140LVT U9207 ( .A1(i_data_bus[473]), .A2(n8626), .B1(
        i_data_bus[249]), .B2(n8687), .ZN(n8585) );
  AOI22D1BWP30P140LVT U9208 ( .A1(i_data_bus[185]), .A2(n8716), .B1(
        i_data_bus[441]), .B2(n8717), .ZN(n8584) );
  AOI22D1BWP30P140LVT U9209 ( .A1(i_data_bus[569]), .A2(n8723), .B1(
        i_data_bus[633]), .B2(n8720), .ZN(n8583) );
  AOI22D1BWP30P140LVT U9210 ( .A1(i_data_bus[601]), .A2(n8722), .B1(
        i_data_bus[537]), .B2(n8721), .ZN(n8582) );
  ND4D1BWP30P140LVT U9211 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), 
        .ZN(n8586) );
  NR4D0BWP30P140LVT U9212 ( .A1(n8589), .A2(n8588), .A3(n8587), .A4(n8586), 
        .ZN(n8590) );
  ND4D4BWP30P140LVT U9213 ( .A1(n8593), .A2(n8592), .A3(n8591), .A4(n8590), 
        .ZN(o_data_bus[185]) );
  AOI22D1BWP30P140LVT U9214 ( .A1(i_data_bus[77]), .A2(n8694), .B1(
        i_data_bus[813]), .B2(n8695), .ZN(n8614) );
  AOI22D1BWP30P140LVT U9215 ( .A1(i_data_bus[365]), .A2(n8701), .B1(
        i_data_bus[877]), .B2(n8706), .ZN(n8613) );
  AOI22D1BWP30P140LVT U9216 ( .A1(i_data_bus[141]), .A2(n8688), .B1(
        i_data_bus[461]), .B2(n8626), .ZN(n8612) );
  AOI22D1BWP30P140LVT U9217 ( .A1(i_data_bus[749]), .A2(n8696), .B1(
        i_data_bus[717]), .B2(n8703), .ZN(n8597) );
  AOI22D1BWP30P140LVT U9218 ( .A1(i_data_bus[1005]), .A2(n8702), .B1(
        i_data_bus[653]), .B2(n8693), .ZN(n8596) );
  AOI22D1BWP30P140LVT U9219 ( .A1(i_data_bus[909]), .A2(n8686), .B1(
        i_data_bus[301]), .B2(n8705), .ZN(n8595) );
  AOI22D1BWP30P140LVT U9220 ( .A1(i_data_bus[973]), .A2(n8708), .B1(
        i_data_bus[109]), .B2(n8692), .ZN(n8594) );
  ND4D1BWP30P140LVT U9221 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), 
        .ZN(n8610) );
  AOI22D1BWP30P140LVT U9222 ( .A1(i_data_bus[269]), .A2(n8691), .B1(
        i_data_bus[845]), .B2(n8690), .ZN(n8601) );
  AOI22D1BWP30P140LVT U9223 ( .A1(i_data_bus[45]), .A2(n8684), .B1(
        i_data_bus[685]), .B2(n8689), .ZN(n8600) );
  AOI22D1BWP30P140LVT U9224 ( .A1(i_data_bus[941]), .A2(n8704), .B1(
        i_data_bus[781]), .B2(n8707), .ZN(n8599) );
  AOI22D1BWP30P140LVT U9225 ( .A1(i_data_bus[13]), .A2(n8683), .B1(
        i_data_bus[333]), .B2(n8685), .ZN(n8598) );
  ND4D1BWP30P140LVT U9226 ( .A1(n8601), .A2(n8600), .A3(n8599), .A4(n8598), 
        .ZN(n8609) );
  INVD1BWP30P140LVT U9227 ( .I(i_data_bus[173]), .ZN(n9420) );
  OAI22D1BWP30P140LVT U9228 ( .A1(n8866), .A2(n8624), .B1(n9420), .B2(n8602), 
        .ZN(n8608) );
  AOI22D1BWP30P140LVT U9229 ( .A1(i_data_bus[237]), .A2(n8687), .B1(
        i_data_bus[397]), .B2(n8719), .ZN(n8606) );
  AOI22D1BWP30P140LVT U9230 ( .A1(i_data_bus[429]), .A2(n8717), .B1(
        i_data_bus[205]), .B2(n8713), .ZN(n8605) );
  AOI22D1BWP30P140LVT U9231 ( .A1(i_data_bus[525]), .A2(n8721), .B1(
        i_data_bus[557]), .B2(n8723), .ZN(n8604) );
  AOI22D1BWP30P140LVT U9232 ( .A1(i_data_bus[621]), .A2(n8720), .B1(
        i_data_bus[589]), .B2(n8722), .ZN(n8603) );
  ND4D1BWP30P140LVT U9233 ( .A1(n8606), .A2(n8605), .A3(n8604), .A4(n8603), 
        .ZN(n8607) );
  NR4D0BWP30P140LVT U9234 ( .A1(n8610), .A2(n8609), .A3(n8608), .A4(n8607), 
        .ZN(n8611) );
  ND4D4BWP30P140LVT U9235 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), 
        .ZN(o_data_bus[173]) );
  AOI22D1BWP30P140LVT U9236 ( .A1(i_data_bus[775]), .A2(n8707), .B1(
        i_data_bus[295]), .B2(n8705), .ZN(n8638) );
  AOI22D1BWP30P140LVT U9237 ( .A1(i_data_bus[967]), .A2(n8708), .B1(
        i_data_bus[935]), .B2(n8704), .ZN(n8637) );
  AOI22D1BWP30P140LVT U9238 ( .A1(i_data_bus[391]), .A2(n8719), .B1(
        i_data_bus[135]), .B2(n8688), .ZN(n8636) );
  AOI22D1BWP30P140LVT U9239 ( .A1(i_data_bus[871]), .A2(n8706), .B1(
        i_data_bus[679]), .B2(n8689), .ZN(n8618) );
  AOI22D1BWP30P140LVT U9240 ( .A1(i_data_bus[359]), .A2(n8701), .B1(
        i_data_bus[327]), .B2(n8685), .ZN(n8617) );
  AOI22D1BWP30P140LVT U9241 ( .A1(i_data_bus[263]), .A2(n8691), .B1(
        i_data_bus[807]), .B2(n8695), .ZN(n8616) );
  AOI22D1BWP30P140LVT U9242 ( .A1(i_data_bus[7]), .A2(n8683), .B1(
        i_data_bus[71]), .B2(n8694), .ZN(n8615) );
  ND4D1BWP30P140LVT U9243 ( .A1(n8618), .A2(n8617), .A3(n8616), .A4(n8615), 
        .ZN(n8634) );
  AOI22D1BWP30P140LVT U9244 ( .A1(i_data_bus[839]), .A2(n8690), .B1(
        i_data_bus[647]), .B2(n8693), .ZN(n8622) );
  AOI22D1BWP30P140LVT U9245 ( .A1(i_data_bus[903]), .A2(n8686), .B1(
        i_data_bus[743]), .B2(n8696), .ZN(n8621) );
  AOI22D1BWP30P140LVT U9246 ( .A1(i_data_bus[103]), .A2(n8692), .B1(
        i_data_bus[999]), .B2(n8702), .ZN(n8620) );
  AOI22D1BWP30P140LVT U9247 ( .A1(i_data_bus[39]), .A2(n8684), .B1(
        i_data_bus[711]), .B2(n8703), .ZN(n8619) );
  ND4D1BWP30P140LVT U9248 ( .A1(n8622), .A2(n8621), .A3(n8620), .A4(n8619), 
        .ZN(n8633) );
  INVD1BWP30P140LVT U9249 ( .I(i_data_bus[199]), .ZN(n9484) );
  OAI22D1BWP30P140LVT U9250 ( .A1(n8625), .A2(n8624), .B1(n9484), .B2(n8623), 
        .ZN(n8632) );
  AOI22D1BWP30P140LVT U9251 ( .A1(i_data_bus[167]), .A2(n8716), .B1(
        i_data_bus[231]), .B2(n8687), .ZN(n8630) );
  AOI22D1BWP30P140LVT U9252 ( .A1(i_data_bus[455]), .A2(n8626), .B1(
        i_data_bus[423]), .B2(n8717), .ZN(n8629) );
  AOI22D1BWP30P140LVT U9253 ( .A1(i_data_bus[615]), .A2(n8720), .B1(
        i_data_bus[551]), .B2(n8723), .ZN(n8628) );
  AOI22D1BWP30P140LVT U9254 ( .A1(i_data_bus[519]), .A2(n8721), .B1(
        i_data_bus[583]), .B2(n8722), .ZN(n8627) );
  ND4D1BWP30P140LVT U9255 ( .A1(n8630), .A2(n8629), .A3(n8628), .A4(n8627), 
        .ZN(n8631) );
  NR4D0BWP30P140LVT U9256 ( .A1(n8634), .A2(n8633), .A3(n8632), .A4(n8631), 
        .ZN(n8635) );
  ND4D4BWP30P140LVT U9257 ( .A1(n8638), .A2(n8637), .A3(n8636), .A4(n8635), 
        .ZN(o_data_bus[167]) );
  AOI22D1BWP30P140LVT U9258 ( .A1(i_data_bus[4]), .A2(n8683), .B1(
        i_data_bus[740]), .B2(n8696), .ZN(n8660) );
  AOI22D1BWP30P140LVT U9259 ( .A1(i_data_bus[964]), .A2(n8708), .B1(
        i_data_bus[932]), .B2(n8704), .ZN(n8659) );
  AOI22D1BWP30P140LVT U9260 ( .A1(i_data_bus[132]), .A2(n8688), .B1(
        i_data_bus[420]), .B2(n8717), .ZN(n8658) );
  AOI22D1BWP30P140LVT U9261 ( .A1(i_data_bus[996]), .A2(n8702), .B1(
        i_data_bus[324]), .B2(n8685), .ZN(n8642) );
  AOI22D1BWP30P140LVT U9262 ( .A1(i_data_bus[68]), .A2(n8694), .B1(
        i_data_bus[644]), .B2(n8693), .ZN(n8641) );
  AOI22D1BWP30P140LVT U9263 ( .A1(i_data_bus[676]), .A2(n8689), .B1(
        i_data_bus[836]), .B2(n8690), .ZN(n8640) );
  AOI22D1BWP30P140LVT U9264 ( .A1(i_data_bus[356]), .A2(n8701), .B1(
        i_data_bus[260]), .B2(n8691), .ZN(n8639) );
  ND4D1BWP30P140LVT U9265 ( .A1(n8642), .A2(n8641), .A3(n8640), .A4(n8639), 
        .ZN(n8656) );
  AOI22D1BWP30P140LVT U9266 ( .A1(i_data_bus[772]), .A2(n8707), .B1(
        i_data_bus[804]), .B2(n8695), .ZN(n8646) );
  AOI22D1BWP30P140LVT U9267 ( .A1(i_data_bus[900]), .A2(n8686), .B1(
        i_data_bus[36]), .B2(n8684), .ZN(n8645) );
  AOI22D1BWP30P140LVT U9268 ( .A1(i_data_bus[100]), .A2(n8692), .B1(
        i_data_bus[868]), .B2(n8706), .ZN(n8644) );
  AOI22D1BWP30P140LVT U9269 ( .A1(i_data_bus[708]), .A2(n8703), .B1(
        i_data_bus[292]), .B2(n8705), .ZN(n8643) );
  ND4D1BWP30P140LVT U9270 ( .A1(n8646), .A2(n8645), .A3(n8644), .A4(n8643), 
        .ZN(n8655) );
  OAI22D1BWP30P140LVT U9271 ( .A1(n9527), .A2(n8714), .B1(n8648), .B2(n8647), 
        .ZN(n8654) );
  AOI22D1BWP30P140LVT U9272 ( .A1(i_data_bus[228]), .A2(n8687), .B1(
        i_data_bus[164]), .B2(n8716), .ZN(n8652) );
  AOI22D1BWP30P140LVT U9273 ( .A1(i_data_bus[196]), .A2(n8713), .B1(
        i_data_bus[484]), .B2(n8718), .ZN(n8651) );
  AOI22D1BWP30P140LVT U9274 ( .A1(i_data_bus[548]), .A2(n8723), .B1(
        i_data_bus[612]), .B2(n8720), .ZN(n8650) );
  AOI22D1BWP30P140LVT U9275 ( .A1(i_data_bus[516]), .A2(n8721), .B1(
        i_data_bus[580]), .B2(n8722), .ZN(n8649) );
  ND4D1BWP30P140LVT U9276 ( .A1(n8652), .A2(n8651), .A3(n8650), .A4(n8649), 
        .ZN(n8653) );
  NR4D0BWP30P140LVT U9277 ( .A1(n8656), .A2(n8655), .A3(n8654), .A4(n8653), 
        .ZN(n8657) );
  ND4D4BWP30P140LVT U9278 ( .A1(n8660), .A2(n8659), .A3(n8658), .A4(n8657), 
        .ZN(o_data_bus[164]) );
  AOI22D1BWP30P140LVT U9279 ( .A1(i_data_bus[771]), .A2(n8707), .B1(
        i_data_bus[803]), .B2(n8695), .ZN(n8682) );
  AOI22D1BWP30P140LVT U9280 ( .A1(i_data_bus[867]), .A2(n8706), .B1(
        i_data_bus[707]), .B2(n8703), .ZN(n8681) );
  AOI22D1BWP30P140LVT U9281 ( .A1(i_data_bus[387]), .A2(n8719), .B1(
        i_data_bus[483]), .B2(n8718), .ZN(n8680) );
  AOI22D1BWP30P140LVT U9282 ( .A1(i_data_bus[355]), .A2(n8701), .B1(
        i_data_bus[291]), .B2(n8705), .ZN(n8664) );
  AOI22D1BWP30P140LVT U9283 ( .A1(i_data_bus[259]), .A2(n8691), .B1(
        i_data_bus[323]), .B2(n8685), .ZN(n8663) );
  AOI22D1BWP30P140LVT U9284 ( .A1(i_data_bus[995]), .A2(n8702), .B1(
        i_data_bus[643]), .B2(n8693), .ZN(n8662) );
  AOI22D1BWP30P140LVT U9285 ( .A1(i_data_bus[99]), .A2(n8692), .B1(
        i_data_bus[835]), .B2(n8690), .ZN(n8661) );
  ND4D1BWP30P140LVT U9286 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), 
        .ZN(n8678) );
  AOI22D1BWP30P140LVT U9287 ( .A1(i_data_bus[67]), .A2(n8694), .B1(
        i_data_bus[675]), .B2(n8689), .ZN(n8668) );
  AOI22D1BWP30P140LVT U9288 ( .A1(i_data_bus[899]), .A2(n8686), .B1(
        i_data_bus[3]), .B2(n8683), .ZN(n8667) );
  AOI22D1BWP30P140LVT U9289 ( .A1(i_data_bus[931]), .A2(n8704), .B1(
        i_data_bus[739]), .B2(n8696), .ZN(n8666) );
  AOI22D1BWP30P140LVT U9290 ( .A1(i_data_bus[35]), .A2(n8684), .B1(
        i_data_bus[963]), .B2(n8708), .ZN(n8665) );
  ND4D1BWP30P140LVT U9291 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), 
        .ZN(n8677) );
  INVD1BWP30P140LVT U9292 ( .I(i_data_bus[131]), .ZN(n9565) );
  OAI22D1BWP30P140LVT U9293 ( .A1(n9565), .A2(n8670), .B1(n8669), .B2(n8714), 
        .ZN(n8676) );
  AOI22D1BWP30P140LVT U9294 ( .A1(i_data_bus[163]), .A2(n8716), .B1(
        i_data_bus[195]), .B2(n8713), .ZN(n8674) );
  AOI22D1BWP30P140LVT U9295 ( .A1(i_data_bus[419]), .A2(n8717), .B1(
        i_data_bus[227]), .B2(n8687), .ZN(n8673) );
  AOI22D1BWP30P140LVT U9296 ( .A1(i_data_bus[515]), .A2(n8721), .B1(
        i_data_bus[547]), .B2(n8723), .ZN(n8672) );
  AOI22D1BWP30P140LVT U9297 ( .A1(i_data_bus[579]), .A2(n8722), .B1(
        i_data_bus[611]), .B2(n8720), .ZN(n8671) );
  ND4D1BWP30P140LVT U9298 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), 
        .ZN(n8675) );
  NR4D0BWP30P140LVT U9299 ( .A1(n8678), .A2(n8677), .A3(n8676), .A4(n8675), 
        .ZN(n8679) );
  ND4D4BWP30P140LVT U9300 ( .A1(n8682), .A2(n8681), .A3(n8680), .A4(n8679), 
        .ZN(o_data_bus[163]) );
  AOI22D1BWP30P140LVT U9301 ( .A1(i_data_bus[32]), .A2(n8684), .B1(
        i_data_bus[0]), .B2(n8683), .ZN(n8735) );
  AOI22D1BWP30P140LVT U9302 ( .A1(i_data_bus[896]), .A2(n8686), .B1(
        i_data_bus[320]), .B2(n8685), .ZN(n8734) );
  AOI22D1BWP30P140LVT U9303 ( .A1(i_data_bus[128]), .A2(n8688), .B1(
        i_data_bus[224]), .B2(n8687), .ZN(n8733) );
  AOI22D1BWP30P140LVT U9304 ( .A1(i_data_bus[832]), .A2(n8690), .B1(
        i_data_bus[672]), .B2(n8689), .ZN(n8700) );
  AOI22D1BWP30P140LVT U9305 ( .A1(i_data_bus[96]), .A2(n8692), .B1(
        i_data_bus[256]), .B2(n8691), .ZN(n8699) );
  AOI22D1BWP30P140LVT U9306 ( .A1(i_data_bus[64]), .A2(n8694), .B1(
        i_data_bus[640]), .B2(n8693), .ZN(n8698) );
  AOI22D1BWP30P140LVT U9307 ( .A1(i_data_bus[736]), .A2(n8696), .B1(
        i_data_bus[800]), .B2(n8695), .ZN(n8697) );
  ND4D1BWP30P140LVT U9308 ( .A1(n8700), .A2(n8699), .A3(n8698), .A4(n8697), 
        .ZN(n8731) );
  AOI22D1BWP30P140LVT U9309 ( .A1(i_data_bus[992]), .A2(n8702), .B1(
        i_data_bus[352]), .B2(n8701), .ZN(n8712) );
  AOI22D1BWP30P140LVT U9310 ( .A1(i_data_bus[928]), .A2(n8704), .B1(
        i_data_bus[704]), .B2(n8703), .ZN(n8711) );
  AOI22D1BWP30P140LVT U9311 ( .A1(i_data_bus[864]), .A2(n8706), .B1(
        i_data_bus[288]), .B2(n8705), .ZN(n8710) );
  AOI22D1BWP30P140LVT U9312 ( .A1(i_data_bus[960]), .A2(n8708), .B1(
        i_data_bus[768]), .B2(n8707), .ZN(n8709) );
  ND4D1BWP30P140LVT U9313 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), 
        .ZN(n8730) );
  MOAI22D1BWP30P140LVT U9314 ( .A1(n8715), .A2(n8714), .B1(i_data_bus[192]), 
        .B2(n8713), .ZN(n8729) );
  AOI22D1BWP30P140LVT U9315 ( .A1(i_data_bus[416]), .A2(n8717), .B1(
        i_data_bus[160]), .B2(n8716), .ZN(n8727) );
  AOI22D1BWP30P140LVT U9316 ( .A1(i_data_bus[384]), .A2(n8719), .B1(
        i_data_bus[480]), .B2(n8718), .ZN(n8726) );
  AOI22D1BWP30P140LVT U9317 ( .A1(i_data_bus[512]), .A2(n8721), .B1(
        i_data_bus[608]), .B2(n8720), .ZN(n8725) );
  AOI22D1BWP30P140LVT U9318 ( .A1(i_data_bus[544]), .A2(n8723), .B1(
        i_data_bus[576]), .B2(n8722), .ZN(n8724) );
  ND4D1BWP30P140LVT U9319 ( .A1(n8727), .A2(n8726), .A3(n8725), .A4(n8724), 
        .ZN(n8728) );
  NR4D0BWP30P140LVT U9320 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), 
        .ZN(n8732) );
  ND4D4BWP30P140LVT U9321 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), 
        .ZN(o_data_bus[160]) );
  AOI22D1BWP30P140LVT U9322 ( .A1(i_data_bus[29]), .A2(n9676), .B1(
        i_data_bus[93]), .B2(n9672), .ZN(n8756) );
  AOI22D1BWP30P140LVT U9323 ( .A1(i_data_bus[957]), .A2(n9669), .B1(
        i_data_bus[1021]), .B2(n9677), .ZN(n8755) );
  AOI22D1BWP30P140LVT U9324 ( .A1(i_data_bus[765]), .A2(n9706), .B1(
        i_data_bus[829]), .B2(n9674), .ZN(n8754) );
  AOI22D1BWP30P140LVT U9325 ( .A1(i_data_bus[61]), .A2(n9670), .B1(
        i_data_bus[157]), .B2(n9681), .ZN(n8739) );
  AOI22D1BWP30P140LVT U9326 ( .A1(i_data_bus[925]), .A2(n9682), .B1(
        i_data_bus[189]), .B2(n9675), .ZN(n8738) );
  AOI22D1BWP30P140LVT U9327 ( .A1(i_data_bus[989]), .A2(n9678), .B1(
        i_data_bus[253]), .B2(n9671), .ZN(n8737) );
  AOI22D1BWP30P140LVT U9328 ( .A1(i_data_bus[125]), .A2(n9680), .B1(
        i_data_bus[221]), .B2(n9679), .ZN(n8736) );
  ND4D1BWP30P140LVT U9329 ( .A1(n8739), .A2(n8738), .A3(n8737), .A4(n8736), 
        .ZN(n8752) );
  MOAI22D1BWP30P140LVT U9330 ( .A1(n8740), .A2(n9181), .B1(i_data_bus[733]), 
        .B2(n9704), .ZN(n8751) );
  AOI22D1BWP30P140LVT U9331 ( .A1(i_data_bus[349]), .A2(n9692), .B1(
        i_data_bus[477]), .B2(n9703), .ZN(n8744) );
  AOI22D1BWP30P140LVT U9332 ( .A1(i_data_bus[509]), .A2(n9656), .B1(
        i_data_bus[797]), .B2(n9673), .ZN(n8743) );
  AOI22D1BWP30P140LVT U9333 ( .A1(i_data_bus[637]), .A2(n9696), .B1(
        i_data_bus[541]), .B2(n9698), .ZN(n8742) );
  AOI22D1BWP30P140LVT U9334 ( .A1(i_data_bus[573]), .A2(n9695), .B1(
        i_data_bus[605]), .B2(n9697), .ZN(n8741) );
  ND4D1BWP30P140LVT U9335 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), 
        .ZN(n8750) );
  AOI22D1BWP30P140LVT U9336 ( .A1(i_data_bus[445]), .A2(n9709), .B1(
        i_data_bus[381]), .B2(n9691), .ZN(n8748) );
  AOI22D1BWP30P140LVT U9337 ( .A1(i_data_bus[669]), .A2(n9707), .B1(
        i_data_bus[317]), .B2(n9655), .ZN(n8747) );
  AOI22D1BWP30P140LVT U9338 ( .A1(i_data_bus[701]), .A2(n9705), .B1(
        i_data_bus[413]), .B2(n9708), .ZN(n8746) );
  AOI22D1BWP30P140LVT U9339 ( .A1(i_data_bus[861]), .A2(n9693), .B1(
        i_data_bus[893]), .B2(n9710), .ZN(n8745) );
  ND4D1BWP30P140LVT U9340 ( .A1(n8748), .A2(n8747), .A3(n8746), .A4(n8745), 
        .ZN(n8749) );
  NR4D0BWP30P140LVT U9341 ( .A1(n8752), .A2(n8751), .A3(n8750), .A4(n8749), 
        .ZN(n8753) );
  ND4D4BWP30P140LVT U9342 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), 
        .ZN(o_data_bus[29]) );
  AOI22D1BWP30P140LVT U9343 ( .A1(i_data_bus[121]), .A2(n9680), .B1(
        i_data_bus[249]), .B2(n9671), .ZN(n8777) );
  AOI22D1BWP30P140LVT U9344 ( .A1(i_data_bus[1017]), .A2(n9677), .B1(
        i_data_bus[89]), .B2(n9672), .ZN(n8776) );
  AOI22D1BWP30P140LVT U9345 ( .A1(i_data_bus[665]), .A2(n9707), .B1(
        i_data_bus[857]), .B2(n9693), .ZN(n8775) );
  AOI22D1BWP30P140LVT U9346 ( .A1(i_data_bus[25]), .A2(n9676), .B1(
        i_data_bus[153]), .B2(n9681), .ZN(n8760) );
  AOI22D1BWP30P140LVT U9347 ( .A1(i_data_bus[57]), .A2(n9670), .B1(
        i_data_bus[921]), .B2(n9682), .ZN(n8759) );
  AOI22D1BWP30P140LVT U9348 ( .A1(i_data_bus[953]), .A2(n9669), .B1(
        i_data_bus[185]), .B2(n9675), .ZN(n8758) );
  AOI22D1BWP30P140LVT U9349 ( .A1(i_data_bus[985]), .A2(n9678), .B1(
        i_data_bus[217]), .B2(n9679), .ZN(n8757) );
  ND4D1BWP30P140LVT U9350 ( .A1(n8760), .A2(n8759), .A3(n8758), .A4(n8757), 
        .ZN(n8773) );
  INVD1BWP30P140LVT U9351 ( .I(n9656), .ZN(n9689) );
  MOAI22D1BWP30P140LVT U9352 ( .A1(n8761), .A2(n9689), .B1(i_data_bus[729]), 
        .B2(n9704), .ZN(n8772) );
  AOI22D1BWP30P140LVT U9353 ( .A1(i_data_bus[345]), .A2(n9692), .B1(
        i_data_bus[761]), .B2(n9706), .ZN(n8765) );
  AOI22D1BWP30P140LVT U9354 ( .A1(i_data_bus[793]), .A2(n9673), .B1(
        i_data_bus[281]), .B2(n9694), .ZN(n8764) );
  AOI22D1BWP30P140LVT U9355 ( .A1(i_data_bus[569]), .A2(n9695), .B1(
        i_data_bus[601]), .B2(n9697), .ZN(n8763) );
  AOI22D1BWP30P140LVT U9356 ( .A1(i_data_bus[633]), .A2(n9696), .B1(
        i_data_bus[537]), .B2(n9698), .ZN(n8762) );
  ND4D1BWP30P140LVT U9357 ( .A1(n8765), .A2(n8764), .A3(n8763), .A4(n8762), 
        .ZN(n8771) );
  AOI22D1BWP30P140LVT U9358 ( .A1(i_data_bus[825]), .A2(n9674), .B1(
        i_data_bus[409]), .B2(n9708), .ZN(n8769) );
  AOI22D1BWP30P140LVT U9359 ( .A1(i_data_bus[377]), .A2(n9691), .B1(
        i_data_bus[473]), .B2(n9703), .ZN(n8768) );
  AOI22D1BWP30P140LVT U9360 ( .A1(i_data_bus[313]), .A2(n9655), .B1(
        i_data_bus[441]), .B2(n9709), .ZN(n8767) );
  AOI22D1BWP30P140LVT U9361 ( .A1(i_data_bus[697]), .A2(n9705), .B1(
        i_data_bus[889]), .B2(n9710), .ZN(n8766) );
  ND4D1BWP30P140LVT U9362 ( .A1(n8769), .A2(n8768), .A3(n8767), .A4(n8766), 
        .ZN(n8770) );
  NR4D0BWP30P140LVT U9363 ( .A1(n8773), .A2(n8772), .A3(n8771), .A4(n8770), 
        .ZN(n8774) );
  ND4D4BWP30P140LVT U9364 ( .A1(n8777), .A2(n8776), .A3(n8775), .A4(n8774), 
        .ZN(o_data_bus[25]) );
  AOI22D1BWP30P140LVT U9365 ( .A1(i_data_bus[152]), .A2(n9681), .B1(
        i_data_bus[184]), .B2(n9675), .ZN(n8798) );
  AOI22D1BWP30P140LVT U9366 ( .A1(i_data_bus[120]), .A2(n9680), .B1(
        i_data_bus[248]), .B2(n9671), .ZN(n8797) );
  AOI22D1BWP30P140LVT U9367 ( .A1(i_data_bus[408]), .A2(n9708), .B1(
        i_data_bus[664]), .B2(n9707), .ZN(n8796) );
  AOI22D1BWP30P140LVT U9368 ( .A1(i_data_bus[1016]), .A2(n9677), .B1(
        i_data_bus[24]), .B2(n9676), .ZN(n8781) );
  AOI22D1BWP30P140LVT U9369 ( .A1(i_data_bus[56]), .A2(n9670), .B1(
        i_data_bus[920]), .B2(n9682), .ZN(n8780) );
  AOI22D1BWP30P140LVT U9370 ( .A1(i_data_bus[984]), .A2(n9678), .B1(
        i_data_bus[88]), .B2(n9672), .ZN(n8779) );
  AOI22D1BWP30P140LVT U9371 ( .A1(i_data_bus[952]), .A2(n9669), .B1(
        i_data_bus[216]), .B2(n9679), .ZN(n8778) );
  ND4D1BWP30P140LVT U9372 ( .A1(n8781), .A2(n8780), .A3(n8779), .A4(n8778), 
        .ZN(n8794) );
  MOAI22D1BWP30P140LVT U9373 ( .A1(n8782), .A2(n9687), .B1(i_data_bus[728]), 
        .B2(n9704), .ZN(n8793) );
  AOI22D1BWP30P140LVT U9374 ( .A1(i_data_bus[792]), .A2(n9673), .B1(
        i_data_bus[824]), .B2(n9674), .ZN(n8786) );
  AOI22D1BWP30P140LVT U9375 ( .A1(i_data_bus[344]), .A2(n9692), .B1(
        i_data_bus[376]), .B2(n9691), .ZN(n8785) );
  AOI22D1BWP30P140LVT U9376 ( .A1(i_data_bus[632]), .A2(n9696), .B1(
        i_data_bus[536]), .B2(n9698), .ZN(n8784) );
  AOI22D1BWP30P140LVT U9377 ( .A1(i_data_bus[600]), .A2(n9697), .B1(
        i_data_bus[568]), .B2(n9695), .ZN(n8783) );
  ND4D1BWP30P140LVT U9378 ( .A1(n8786), .A2(n8785), .A3(n8784), .A4(n8783), 
        .ZN(n8792) );
  AOI22D1BWP30P140LVT U9379 ( .A1(i_data_bus[280]), .A2(n9694), .B1(
        i_data_bus[472]), .B2(n9703), .ZN(n8790) );
  AOI22D1BWP30P140LVT U9380 ( .A1(i_data_bus[856]), .A2(n9693), .B1(
        i_data_bus[504]), .B2(n9656), .ZN(n8789) );
  AOI22D1BWP30P140LVT U9381 ( .A1(i_data_bus[696]), .A2(n9705), .B1(
        i_data_bus[888]), .B2(n9710), .ZN(n8788) );
  AOI22D1BWP30P140LVT U9382 ( .A1(i_data_bus[440]), .A2(n9709), .B1(
        i_data_bus[760]), .B2(n9706), .ZN(n8787) );
  ND4D1BWP30P140LVT U9383 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), 
        .ZN(n8791) );
  NR4D0BWP30P140LVT U9384 ( .A1(n8794), .A2(n8793), .A3(n8792), .A4(n8791), 
        .ZN(n8795) );
  ND4D4BWP30P140LVT U9385 ( .A1(n8798), .A2(n8797), .A3(n8796), .A4(n8795), 
        .ZN(o_data_bus[24]) );
  AOI22D1BWP30P140LVT U9386 ( .A1(i_data_bus[182]), .A2(n9675), .B1(
        i_data_bus[214]), .B2(n9679), .ZN(n8820) );
  AOI22D1BWP30P140LVT U9387 ( .A1(i_data_bus[54]), .A2(n9670), .B1(
        i_data_bus[22]), .B2(n9676), .ZN(n8819) );
  AOI22D1BWP30P140LVT U9388 ( .A1(i_data_bus[310]), .A2(n9655), .B1(
        i_data_bus[854]), .B2(n9693), .ZN(n8818) );
  AOI22D1BWP30P140LVT U9389 ( .A1(i_data_bus[918]), .A2(n9682), .B1(
        i_data_bus[950]), .B2(n9669), .ZN(n8802) );
  AOI22D1BWP30P140LVT U9390 ( .A1(i_data_bus[246]), .A2(n9671), .B1(
        i_data_bus[150]), .B2(n9681), .ZN(n8801) );
  AOI22D1BWP30P140LVT U9391 ( .A1(i_data_bus[118]), .A2(n9680), .B1(
        i_data_bus[86]), .B2(n9672), .ZN(n8800) );
  AOI22D1BWP30P140LVT U9392 ( .A1(i_data_bus[1014]), .A2(n9677), .B1(
        i_data_bus[982]), .B2(n9678), .ZN(n8799) );
  ND4D1BWP30P140LVT U9393 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), 
        .ZN(n8816) );
  OAI22D1BWP30P140LVT U9394 ( .A1(n8804), .A2(n9649), .B1(n8803), .B2(n9137), 
        .ZN(n8815) );
  AOI22D1BWP30P140LVT U9395 ( .A1(i_data_bus[438]), .A2(n9709), .B1(
        i_data_bus[374]), .B2(n9691), .ZN(n8808) );
  AOI22D1BWP30P140LVT U9396 ( .A1(i_data_bus[822]), .A2(n9674), .B1(
        i_data_bus[758]), .B2(n9706), .ZN(n8807) );
  AOI22D1BWP30P140LVT U9397 ( .A1(i_data_bus[534]), .A2(n9698), .B1(
        i_data_bus[598]), .B2(n9697), .ZN(n8806) );
  AOI22D1BWP30P140LVT U9398 ( .A1(i_data_bus[566]), .A2(n9695), .B1(
        i_data_bus[630]), .B2(n9696), .ZN(n8805) );
  ND4D1BWP30P140LVT U9399 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), 
        .ZN(n8814) );
  AOI22D1BWP30P140LVT U9400 ( .A1(i_data_bus[406]), .A2(n9708), .B1(
        i_data_bus[278]), .B2(n9694), .ZN(n8812) );
  AOI22D1BWP30P140LVT U9401 ( .A1(i_data_bus[790]), .A2(n9673), .B1(
        i_data_bus[502]), .B2(n9656), .ZN(n8811) );
  AOI22D1BWP30P140LVT U9402 ( .A1(i_data_bus[726]), .A2(n9704), .B1(
        i_data_bus[886]), .B2(n9710), .ZN(n8810) );
  AOI22D1BWP30P140LVT U9403 ( .A1(i_data_bus[694]), .A2(n9705), .B1(
        i_data_bus[662]), .B2(n9707), .ZN(n8809) );
  ND4D1BWP30P140LVT U9404 ( .A1(n8812), .A2(n8811), .A3(n8810), .A4(n8809), 
        .ZN(n8813) );
  NR4D0BWP30P140LVT U9405 ( .A1(n8816), .A2(n8815), .A3(n8814), .A4(n8813), 
        .ZN(n8817) );
  ND4D4BWP30P140LVT U9406 ( .A1(n8820), .A2(n8819), .A3(n8818), .A4(n8817), 
        .ZN(o_data_bus[22]) );
  AOI22D1BWP30P140LVT U9407 ( .A1(i_data_bus[84]), .A2(n9672), .B1(
        i_data_bus[180]), .B2(n9675), .ZN(n8840) );
  AOI22D1BWP30P140LVT U9408 ( .A1(i_data_bus[948]), .A2(n9669), .B1(
        i_data_bus[244]), .B2(n9671), .ZN(n8839) );
  AOI22D1BWP30P140LVT U9409 ( .A1(i_data_bus[724]), .A2(n9704), .B1(
        i_data_bus[436]), .B2(n9709), .ZN(n8838) );
  AOI22D1BWP30P140LVT U9410 ( .A1(i_data_bus[660]), .A2(n9707), .B1(
        i_data_bus[404]), .B2(n9708), .ZN(n8836) );
  AOI22D1BWP30P140LVT U9411 ( .A1(i_data_bus[20]), .A2(n9676), .B1(
        i_data_bus[212]), .B2(n9679), .ZN(n8824) );
  AOI22D1BWP30P140LVT U9412 ( .A1(i_data_bus[116]), .A2(n9680), .B1(
        i_data_bus[148]), .B2(n9681), .ZN(n8823) );
  AOI22D1BWP30P140LVT U9413 ( .A1(i_data_bus[980]), .A2(n9678), .B1(
        i_data_bus[1012]), .B2(n9677), .ZN(n8822) );
  AOI22D1BWP30P140LVT U9414 ( .A1(i_data_bus[52]), .A2(n9670), .B1(
        i_data_bus[916]), .B2(n9682), .ZN(n8821) );
  ND4D1BWP30P140LVT U9415 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), 
        .ZN(n8835) );
  AOI22D1BWP30P140LVT U9416 ( .A1(i_data_bus[852]), .A2(n9693), .B1(
        i_data_bus[276]), .B2(n9694), .ZN(n8828) );
  AOI22D1BWP30P140LVT U9417 ( .A1(i_data_bus[756]), .A2(n9706), .B1(
        i_data_bus[500]), .B2(n9656), .ZN(n8827) );
  AOI22D1BWP30P140LVT U9418 ( .A1(i_data_bus[596]), .A2(n9697), .B1(
        i_data_bus[532]), .B2(n9698), .ZN(n8826) );
  AOI22D1BWP30P140LVT U9419 ( .A1(i_data_bus[564]), .A2(n9695), .B1(
        i_data_bus[628]), .B2(n9696), .ZN(n8825) );
  ND4D1BWP30P140LVT U9420 ( .A1(n8828), .A2(n8827), .A3(n8826), .A4(n8825), 
        .ZN(n8834) );
  AOI22D1BWP30P140LVT U9421 ( .A1(i_data_bus[692]), .A2(n9705), .B1(
        i_data_bus[468]), .B2(n9703), .ZN(n8832) );
  AOI22D1BWP30P140LVT U9422 ( .A1(i_data_bus[340]), .A2(n9692), .B1(
        i_data_bus[788]), .B2(n9673), .ZN(n8831) );
  AOI22D1BWP30P140LVT U9423 ( .A1(i_data_bus[820]), .A2(n9674), .B1(
        i_data_bus[308]), .B2(n9655), .ZN(n8830) );
  AOI22D1BWP30P140LVT U9424 ( .A1(i_data_bus[884]), .A2(n9710), .B1(
        i_data_bus[372]), .B2(n9691), .ZN(n8829) );
  ND4D1BWP30P140LVT U9425 ( .A1(n8832), .A2(n8831), .A3(n8830), .A4(n8829), 
        .ZN(n8833) );
  INR4D0BWP30P140LVT U9426 ( .A1(n8836), .B1(n8835), .B2(n8834), .B3(n8833), 
        .ZN(n8837) );
  ND4D4BWP30P140LVT U9427 ( .A1(n8840), .A2(n8839), .A3(n8838), .A4(n8837), 
        .ZN(o_data_bus[20]) );
  AOI22D1BWP30P140LVT U9428 ( .A1(i_data_bus[943]), .A2(n9669), .B1(
        i_data_bus[207]), .B2(n9679), .ZN(n8861) );
  AOI22D1BWP30P140LVT U9429 ( .A1(i_data_bus[975]), .A2(n9678), .B1(
        i_data_bus[175]), .B2(n9675), .ZN(n8860) );
  AOI22D1BWP30P140LVT U9430 ( .A1(i_data_bus[783]), .A2(n9673), .B1(
        i_data_bus[335]), .B2(n9692), .ZN(n8859) );
  AOI22D1BWP30P140LVT U9431 ( .A1(i_data_bus[111]), .A2(n9680), .B1(
        i_data_bus[1007]), .B2(n9677), .ZN(n8844) );
  AOI22D1BWP30P140LVT U9432 ( .A1(i_data_bus[911]), .A2(n9682), .B1(
        i_data_bus[15]), .B2(n9676), .ZN(n8843) );
  AOI22D1BWP30P140LVT U9433 ( .A1(i_data_bus[239]), .A2(n9671), .B1(
        i_data_bus[143]), .B2(n9681), .ZN(n8842) );
  AOI22D1BWP30P140LVT U9434 ( .A1(i_data_bus[79]), .A2(n9672), .B1(
        i_data_bus[47]), .B2(n9670), .ZN(n8841) );
  ND4D1BWP30P140LVT U9435 ( .A1(n8844), .A2(n8843), .A3(n8842), .A4(n8841), 
        .ZN(n8857) );
  MOAI22D1BWP30P140LVT U9436 ( .A1(n8845), .A2(n9626), .B1(i_data_bus[655]), 
        .B2(n9707), .ZN(n8856) );
  AOI22D1BWP30P140LVT U9437 ( .A1(i_data_bus[719]), .A2(n9704), .B1(
        i_data_bus[687]), .B2(n9705), .ZN(n8849) );
  AOI22D1BWP30P140LVT U9438 ( .A1(i_data_bus[847]), .A2(n9693), .B1(
        i_data_bus[303]), .B2(n9655), .ZN(n8848) );
  AOI22D1BWP30P140LVT U9439 ( .A1(i_data_bus[527]), .A2(n9698), .B1(
        i_data_bus[623]), .B2(n9696), .ZN(n8847) );
  AOI22D1BWP30P140LVT U9440 ( .A1(i_data_bus[591]), .A2(n9697), .B1(
        i_data_bus[559]), .B2(n9695), .ZN(n8846) );
  ND4D1BWP30P140LVT U9441 ( .A1(n8849), .A2(n8848), .A3(n8847), .A4(n8846), 
        .ZN(n8855) );
  AOI22D1BWP30P140LVT U9442 ( .A1(i_data_bus[495]), .A2(n9656), .B1(
        i_data_bus[879]), .B2(n9710), .ZN(n8853) );
  AOI22D1BWP30P140LVT U9443 ( .A1(i_data_bus[815]), .A2(n9674), .B1(
        i_data_bus[367]), .B2(n9691), .ZN(n8852) );
  AOI22D1BWP30P140LVT U9444 ( .A1(i_data_bus[271]), .A2(n9694), .B1(
        i_data_bus[463]), .B2(n9703), .ZN(n8851) );
  AOI22D1BWP30P140LVT U9445 ( .A1(i_data_bus[751]), .A2(n9706), .B1(
        i_data_bus[431]), .B2(n9709), .ZN(n8850) );
  ND4D1BWP30P140LVT U9446 ( .A1(n8853), .A2(n8852), .A3(n8851), .A4(n8850), 
        .ZN(n8854) );
  NR4D0BWP30P140LVT U9447 ( .A1(n8857), .A2(n8856), .A3(n8855), .A4(n8854), 
        .ZN(n8858) );
  ND4D4BWP30P140LVT U9448 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), 
        .ZN(o_data_bus[15]) );
  AOI22D1BWP30P140LVT U9449 ( .A1(i_data_bus[109]), .A2(n9680), .B1(
        i_data_bus[173]), .B2(n9675), .ZN(n8882) );
  AOI22D1BWP30P140LVT U9450 ( .A1(i_data_bus[237]), .A2(n9671), .B1(
        i_data_bus[141]), .B2(n9681), .ZN(n8881) );
  AOI22D1BWP30P140LVT U9451 ( .A1(i_data_bus[333]), .A2(n9692), .B1(
        i_data_bus[813]), .B2(n9674), .ZN(n8880) );
  AOI22D1BWP30P140LVT U9452 ( .A1(i_data_bus[45]), .A2(n9670), .B1(
        i_data_bus[77]), .B2(n9672), .ZN(n8865) );
  AOI22D1BWP30P140LVT U9453 ( .A1(i_data_bus[909]), .A2(n9682), .B1(
        i_data_bus[941]), .B2(n9669), .ZN(n8864) );
  AOI22D1BWP30P140LVT U9454 ( .A1(i_data_bus[1005]), .A2(n9677), .B1(
        i_data_bus[13]), .B2(n9676), .ZN(n8863) );
  AOI22D1BWP30P140LVT U9455 ( .A1(i_data_bus[973]), .A2(n9678), .B1(
        i_data_bus[205]), .B2(n9679), .ZN(n8862) );
  ND4D1BWP30P140LVT U9456 ( .A1(n8865), .A2(n8864), .A3(n8863), .A4(n8862), 
        .ZN(n8878) );
  MOAI22D1BWP30P140LVT U9457 ( .A1(n8866), .A2(n9689), .B1(i_data_bus[877]), 
        .B2(n9710), .ZN(n8877) );
  AOI22D1BWP30P140LVT U9458 ( .A1(i_data_bus[429]), .A2(n9709), .B1(
        i_data_bus[845]), .B2(n9693), .ZN(n8870) );
  AOI22D1BWP30P140LVT U9459 ( .A1(i_data_bus[653]), .A2(n9707), .B1(
        i_data_bus[461]), .B2(n9703), .ZN(n8869) );
  AOI22D1BWP30P140LVT U9460 ( .A1(i_data_bus[621]), .A2(n9696), .B1(
        i_data_bus[589]), .B2(n9697), .ZN(n8868) );
  AOI22D1BWP30P140LVT U9461 ( .A1(i_data_bus[525]), .A2(n9698), .B1(
        i_data_bus[557]), .B2(n9695), .ZN(n8867) );
  ND4D1BWP30P140LVT U9462 ( .A1(n8870), .A2(n8869), .A3(n8868), .A4(n8867), 
        .ZN(n8876) );
  AOI22D1BWP30P140LVT U9463 ( .A1(i_data_bus[397]), .A2(n9708), .B1(
        i_data_bus[717]), .B2(n9704), .ZN(n8874) );
  AOI22D1BWP30P140LVT U9464 ( .A1(i_data_bus[269]), .A2(n9694), .B1(
        i_data_bus[781]), .B2(n9673), .ZN(n8873) );
  AOI22D1BWP30P140LVT U9465 ( .A1(i_data_bus[365]), .A2(n9691), .B1(
        i_data_bus[301]), .B2(n9655), .ZN(n8872) );
  AOI22D1BWP30P140LVT U9466 ( .A1(i_data_bus[749]), .A2(n9706), .B1(
        i_data_bus[685]), .B2(n9705), .ZN(n8871) );
  ND4D1BWP30P140LVT U9467 ( .A1(n8874), .A2(n8873), .A3(n8872), .A4(n8871), 
        .ZN(n8875) );
  NR4D0BWP30P140LVT U9468 ( .A1(n8878), .A2(n8877), .A3(n8876), .A4(n8875), 
        .ZN(n8879) );
  ND4D4BWP30P140LVT U9469 ( .A1(n8882), .A2(n8881), .A3(n8880), .A4(n8879), 
        .ZN(o_data_bus[13]) );
  AOI22D1BWP30P140LVT U9470 ( .A1(i_data_bus[74]), .A2(n9672), .B1(
        i_data_bus[170]), .B2(n9675), .ZN(n8903) );
  AOI22D1BWP30P140LVT U9471 ( .A1(i_data_bus[1002]), .A2(n9677), .B1(
        i_data_bus[202]), .B2(n9679), .ZN(n8902) );
  AOI22D1BWP30P140LVT U9472 ( .A1(i_data_bus[298]), .A2(n9655), .B1(
        i_data_bus[426]), .B2(n9709), .ZN(n8901) );
  AOI22D1BWP30P140LVT U9473 ( .A1(i_data_bus[42]), .A2(n9670), .B1(
        i_data_bus[906]), .B2(n9682), .ZN(n8886) );
  AOI22D1BWP30P140LVT U9474 ( .A1(i_data_bus[10]), .A2(n9676), .B1(
        i_data_bus[138]), .B2(n9681), .ZN(n8885) );
  AOI22D1BWP30P140LVT U9475 ( .A1(i_data_bus[106]), .A2(n9680), .B1(
        i_data_bus[938]), .B2(n9669), .ZN(n8884) );
  AOI22D1BWP30P140LVT U9476 ( .A1(i_data_bus[970]), .A2(n9678), .B1(
        i_data_bus[234]), .B2(n9671), .ZN(n8883) );
  ND4D1BWP30P140LVT U9477 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), 
        .ZN(n8899) );
  MOAI22D1BWP30P140LVT U9478 ( .A1(n8887), .A2(n9689), .B1(i_data_bus[458]), 
        .B2(n9703), .ZN(n8898) );
  AOI22D1BWP30P140LVT U9479 ( .A1(i_data_bus[778]), .A2(n9673), .B1(
        i_data_bus[842]), .B2(n9693), .ZN(n8891) );
  AOI22D1BWP30P140LVT U9480 ( .A1(i_data_bus[874]), .A2(n9710), .B1(
        i_data_bus[746]), .B2(n9706), .ZN(n8890) );
  AOI22D1BWP30P140LVT U9481 ( .A1(i_data_bus[618]), .A2(n9696), .B1(
        i_data_bus[586]), .B2(n9697), .ZN(n8889) );
  AOI22D1BWP30P140LVT U9482 ( .A1(i_data_bus[554]), .A2(n9695), .B1(
        i_data_bus[522]), .B2(n9698), .ZN(n8888) );
  ND4D1BWP30P140LVT U9483 ( .A1(n8891), .A2(n8890), .A3(n8889), .A4(n8888), 
        .ZN(n8897) );
  AOI22D1BWP30P140LVT U9484 ( .A1(i_data_bus[362]), .A2(n9691), .B1(
        i_data_bus[266]), .B2(n9694), .ZN(n8895) );
  AOI22D1BWP30P140LVT U9485 ( .A1(i_data_bus[810]), .A2(n9674), .B1(
        i_data_bus[682]), .B2(n9705), .ZN(n8894) );
  AOI22D1BWP30P140LVT U9486 ( .A1(i_data_bus[330]), .A2(n9692), .B1(
        i_data_bus[714]), .B2(n9704), .ZN(n8893) );
  AOI22D1BWP30P140LVT U9487 ( .A1(i_data_bus[650]), .A2(n9707), .B1(
        i_data_bus[394]), .B2(n9708), .ZN(n8892) );
  ND4D1BWP30P140LVT U9488 ( .A1(n8895), .A2(n8894), .A3(n8893), .A4(n8892), 
        .ZN(n8896) );
  NR4D0BWP30P140LVT U9489 ( .A1(n8899), .A2(n8898), .A3(n8897), .A4(n8896), 
        .ZN(n8900) );
  ND4D4BWP30P140LVT U9490 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), 
        .ZN(o_data_bus[10]) );
  AOI22D1BWP30P140LVT U9491 ( .A1(i_data_bus[71]), .A2(n9672), .B1(
        i_data_bus[231]), .B2(n9671), .ZN(n8924) );
  AOI22D1BWP30P140LVT U9492 ( .A1(i_data_bus[967]), .A2(n9678), .B1(
        i_data_bus[999]), .B2(n9677), .ZN(n8923) );
  AOI22D1BWP30P140LVT U9493 ( .A1(i_data_bus[391]), .A2(n9708), .B1(
        i_data_bus[711]), .B2(n9704), .ZN(n8922) );
  AOI22D1BWP30P140LVT U9494 ( .A1(i_data_bus[7]), .A2(n9676), .B1(
        i_data_bus[199]), .B2(n9679), .ZN(n8907) );
  AOI22D1BWP30P140LVT U9495 ( .A1(i_data_bus[39]), .A2(n9670), .B1(
        i_data_bus[135]), .B2(n9681), .ZN(n8906) );
  AOI22D1BWP30P140LVT U9496 ( .A1(i_data_bus[103]), .A2(n9680), .B1(
        i_data_bus[935]), .B2(n9669), .ZN(n8905) );
  AOI22D1BWP30P140LVT U9497 ( .A1(i_data_bus[903]), .A2(n9682), .B1(
        i_data_bus[167]), .B2(n9675), .ZN(n8904) );
  ND4D1BWP30P140LVT U9498 ( .A1(n8907), .A2(n8906), .A3(n8905), .A4(n8904), 
        .ZN(n8920) );
  MOAI22D1BWP30P140LVT U9499 ( .A1(n8908), .A2(n9604), .B1(i_data_bus[423]), 
        .B2(n9709), .ZN(n8919) );
  AOI22D1BWP30P140LVT U9500 ( .A1(i_data_bus[871]), .A2(n9710), .B1(
        i_data_bus[647]), .B2(n9707), .ZN(n8912) );
  AOI22D1BWP30P140LVT U9501 ( .A1(i_data_bus[807]), .A2(n9674), .B1(
        i_data_bus[295]), .B2(n9655), .ZN(n8911) );
  AOI22D1BWP30P140LVT U9502 ( .A1(i_data_bus[519]), .A2(n9698), .B1(
        i_data_bus[583]), .B2(n9697), .ZN(n8910) );
  AOI22D1BWP30P140LVT U9503 ( .A1(i_data_bus[615]), .A2(n9696), .B1(
        i_data_bus[551]), .B2(n9695), .ZN(n8909) );
  ND4D1BWP30P140LVT U9504 ( .A1(n8912), .A2(n8911), .A3(n8910), .A4(n8909), 
        .ZN(n8918) );
  AOI22D1BWP30P140LVT U9505 ( .A1(i_data_bus[455]), .A2(n9703), .B1(
        i_data_bus[775]), .B2(n9673), .ZN(n8916) );
  AOI22D1BWP30P140LVT U9506 ( .A1(i_data_bus[263]), .A2(n9694), .B1(
        i_data_bus[743]), .B2(n9706), .ZN(n8915) );
  AOI22D1BWP30P140LVT U9507 ( .A1(i_data_bus[679]), .A2(n9705), .B1(
        i_data_bus[839]), .B2(n9693), .ZN(n8914) );
  AOI22D1BWP30P140LVT U9508 ( .A1(i_data_bus[487]), .A2(n9656), .B1(
        i_data_bus[327]), .B2(n9692), .ZN(n8913) );
  ND4D1BWP30P140LVT U9509 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), 
        .ZN(n8917) );
  NR4D0BWP30P140LVT U9510 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), 
        .ZN(n8921) );
  ND4D4BWP30P140LVT U9511 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), 
        .ZN(o_data_bus[7]) );
  AOI22D1BWP30P140LVT U9512 ( .A1(i_data_bus[60]), .A2(n9670), .B1(
        i_data_bus[220]), .B2(n9679), .ZN(n8945) );
  AOI22D1BWP30P140LVT U9513 ( .A1(i_data_bus[92]), .A2(n9672), .B1(
        i_data_bus[156]), .B2(n9681), .ZN(n8944) );
  AOI22D1BWP30P140LVT U9514 ( .A1(i_data_bus[508]), .A2(n9656), .B1(
        i_data_bus[700]), .B2(n9705), .ZN(n8943) );
  AOI22D1BWP30P140LVT U9515 ( .A1(i_data_bus[956]), .A2(n9669), .B1(
        i_data_bus[1020]), .B2(n9677), .ZN(n8928) );
  AOI22D1BWP30P140LVT U9516 ( .A1(i_data_bus[988]), .A2(n9678), .B1(
        i_data_bus[252]), .B2(n9671), .ZN(n8927) );
  AOI22D1BWP30P140LVT U9517 ( .A1(i_data_bus[28]), .A2(n9676), .B1(
        i_data_bus[188]), .B2(n9675), .ZN(n8926) );
  AOI22D1BWP30P140LVT U9518 ( .A1(i_data_bus[924]), .A2(n9682), .B1(
        i_data_bus[124]), .B2(n9680), .ZN(n8925) );
  ND4D1BWP30P140LVT U9519 ( .A1(n8928), .A2(n8927), .A3(n8926), .A4(n8925), 
        .ZN(n8941) );
  MOAI22D1BWP30P140LVT U9520 ( .A1(n8929), .A2(n9181), .B1(i_data_bus[316]), 
        .B2(n9655), .ZN(n8940) );
  AOI22D1BWP30P140LVT U9521 ( .A1(i_data_bus[764]), .A2(n9706), .B1(
        i_data_bus[668]), .B2(n9707), .ZN(n8933) );
  AOI22D1BWP30P140LVT U9522 ( .A1(i_data_bus[348]), .A2(n9692), .B1(
        i_data_bus[380]), .B2(n9691), .ZN(n8932) );
  AOI22D1BWP30P140LVT U9523 ( .A1(i_data_bus[636]), .A2(n9696), .B1(
        i_data_bus[572]), .B2(n9695), .ZN(n8931) );
  AOI22D1BWP30P140LVT U9524 ( .A1(i_data_bus[540]), .A2(n9698), .B1(
        i_data_bus[604]), .B2(n9697), .ZN(n8930) );
  ND4D1BWP30P140LVT U9525 ( .A1(n8933), .A2(n8932), .A3(n8931), .A4(n8930), 
        .ZN(n8939) );
  AOI22D1BWP30P140LVT U9526 ( .A1(i_data_bus[828]), .A2(n9674), .B1(
        i_data_bus[860]), .B2(n9693), .ZN(n8937) );
  AOI22D1BWP30P140LVT U9527 ( .A1(i_data_bus[892]), .A2(n9710), .B1(
        i_data_bus[412]), .B2(n9708), .ZN(n8936) );
  AOI22D1BWP30P140LVT U9528 ( .A1(i_data_bus[796]), .A2(n9673), .B1(
        i_data_bus[732]), .B2(n9704), .ZN(n8935) );
  AOI22D1BWP30P140LVT U9529 ( .A1(i_data_bus[444]), .A2(n9709), .B1(
        i_data_bus[476]), .B2(n9703), .ZN(n8934) );
  ND4D1BWP30P140LVT U9530 ( .A1(n8937), .A2(n8936), .A3(n8935), .A4(n8934), 
        .ZN(n8938) );
  NR4D0BWP30P140LVT U9531 ( .A1(n8941), .A2(n8940), .A3(n8939), .A4(n8938), 
        .ZN(n8942) );
  ND4D4BWP30P140LVT U9532 ( .A1(n8945), .A2(n8944), .A3(n8943), .A4(n8942), 
        .ZN(o_data_bus[28]) );
  AOI22D1BWP30P140LVT U9533 ( .A1(i_data_bus[1015]), .A2(n9677), .B1(
        i_data_bus[951]), .B2(n9669), .ZN(n8966) );
  AOI22D1BWP30P140LVT U9534 ( .A1(i_data_bus[119]), .A2(n9680), .B1(
        i_data_bus[215]), .B2(n9679), .ZN(n8965) );
  AOI22D1BWP30P140LVT U9535 ( .A1(i_data_bus[503]), .A2(n9656), .B1(
        i_data_bus[343]), .B2(n9692), .ZN(n8964) );
  AOI22D1BWP30P140LVT U9536 ( .A1(i_data_bus[55]), .A2(n9670), .B1(
        i_data_bus[919]), .B2(n9682), .ZN(n8949) );
  AOI22D1BWP30P140LVT U9537 ( .A1(i_data_bus[983]), .A2(n9678), .B1(
        i_data_bus[151]), .B2(n9681), .ZN(n8948) );
  AOI22D1BWP30P140LVT U9538 ( .A1(i_data_bus[23]), .A2(n9676), .B1(
        i_data_bus[183]), .B2(n9675), .ZN(n8947) );
  AOI22D1BWP30P140LVT U9539 ( .A1(i_data_bus[87]), .A2(n9672), .B1(
        i_data_bus[247]), .B2(n9671), .ZN(n8946) );
  ND4D1BWP30P140LVT U9540 ( .A1(n8949), .A2(n8948), .A3(n8947), .A4(n8946), 
        .ZN(n8962) );
  MOAI22D1BWP30P140LVT U9541 ( .A1(n8950), .A2(n9649), .B1(i_data_bus[823]), 
        .B2(n9674), .ZN(n8961) );
  AOI22D1BWP30P140LVT U9542 ( .A1(i_data_bus[759]), .A2(n9706), .B1(
        i_data_bus[407]), .B2(n9708), .ZN(n8954) );
  AOI22D1BWP30P140LVT U9543 ( .A1(i_data_bus[695]), .A2(n9705), .B1(
        i_data_bus[311]), .B2(n9655), .ZN(n8953) );
  AOI22D1BWP30P140LVT U9544 ( .A1(i_data_bus[631]), .A2(n9696), .B1(
        i_data_bus[599]), .B2(n9697), .ZN(n8952) );
  AOI22D1BWP30P140LVT U9545 ( .A1(i_data_bus[535]), .A2(n9698), .B1(
        i_data_bus[567]), .B2(n9695), .ZN(n8951) );
  ND4D1BWP30P140LVT U9546 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), 
        .ZN(n8960) );
  AOI22D1BWP30P140LVT U9547 ( .A1(i_data_bus[439]), .A2(n9709), .B1(
        i_data_bus[727]), .B2(n9704), .ZN(n8958) );
  AOI22D1BWP30P140LVT U9548 ( .A1(i_data_bus[887]), .A2(n9710), .B1(
        i_data_bus[279]), .B2(n9694), .ZN(n8957) );
  AOI22D1BWP30P140LVT U9549 ( .A1(i_data_bus[663]), .A2(n9707), .B1(
        i_data_bus[375]), .B2(n9691), .ZN(n8956) );
  AOI22D1BWP30P140LVT U9550 ( .A1(i_data_bus[791]), .A2(n9673), .B1(
        i_data_bus[855]), .B2(n9693), .ZN(n8955) );
  ND4D1BWP30P140LVT U9551 ( .A1(n8958), .A2(n8957), .A3(n8956), .A4(n8955), 
        .ZN(n8959) );
  NR4D0BWP30P140LVT U9552 ( .A1(n8962), .A2(n8961), .A3(n8960), .A4(n8959), 
        .ZN(n8963) );
  ND4D4BWP30P140LVT U9553 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), 
        .ZN(o_data_bus[23]) );
  AOI22D1BWP30P140LVT U9554 ( .A1(i_data_bus[12]), .A2(n9676), .B1(
        i_data_bus[140]), .B2(n9681), .ZN(n8988) );
  AOI22D1BWP30P140LVT U9555 ( .A1(i_data_bus[1004]), .A2(n9677), .B1(
        i_data_bus[108]), .B2(n9680), .ZN(n8987) );
  AOI22D1BWP30P140LVT U9556 ( .A1(i_data_bus[780]), .A2(n9673), .B1(
        i_data_bus[332]), .B2(n9692), .ZN(n8986) );
  AOI22D1BWP30P140LVT U9557 ( .A1(i_data_bus[76]), .A2(n9672), .B1(
        i_data_bus[204]), .B2(n9679), .ZN(n8970) );
  AOI22D1BWP30P140LVT U9558 ( .A1(i_data_bus[908]), .A2(n9682), .B1(
        i_data_bus[972]), .B2(n9678), .ZN(n8969) );
  AOI22D1BWP30P140LVT U9559 ( .A1(i_data_bus[940]), .A2(n9669), .B1(
        i_data_bus[172]), .B2(n9675), .ZN(n8968) );
  AOI22D1BWP30P140LVT U9560 ( .A1(i_data_bus[44]), .A2(n9670), .B1(
        i_data_bus[236]), .B2(n9671), .ZN(n8967) );
  ND4D1BWP30P140LVT U9561 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), 
        .ZN(n8984) );
  OAI22D1BWP30P140LVT U9562 ( .A1(n8972), .A2(n9649), .B1(n8971), .B2(n9689), 
        .ZN(n8983) );
  AOI22D1BWP30P140LVT U9563 ( .A1(i_data_bus[652]), .A2(n9707), .B1(
        i_data_bus[876]), .B2(n9710), .ZN(n8976) );
  AOI22D1BWP30P140LVT U9564 ( .A1(i_data_bus[684]), .A2(n9705), .B1(
        i_data_bus[812]), .B2(n9674), .ZN(n8975) );
  AOI22D1BWP30P140LVT U9565 ( .A1(i_data_bus[556]), .A2(n9695), .B1(
        i_data_bus[524]), .B2(n9698), .ZN(n8974) );
  AOI22D1BWP30P140LVT U9566 ( .A1(i_data_bus[620]), .A2(n9696), .B1(
        i_data_bus[588]), .B2(n9697), .ZN(n8973) );
  ND4D1BWP30P140LVT U9567 ( .A1(n8976), .A2(n8975), .A3(n8974), .A4(n8973), 
        .ZN(n8982) );
  AOI22D1BWP30P140LVT U9568 ( .A1(i_data_bus[300]), .A2(n9655), .B1(
        i_data_bus[364]), .B2(n9691), .ZN(n8980) );
  AOI22D1BWP30P140LVT U9569 ( .A1(i_data_bus[428]), .A2(n9709), .B1(
        i_data_bus[268]), .B2(n9694), .ZN(n8979) );
  AOI22D1BWP30P140LVT U9570 ( .A1(i_data_bus[748]), .A2(n9706), .B1(
        i_data_bus[396]), .B2(n9708), .ZN(n8978) );
  AOI22D1BWP30P140LVT U9571 ( .A1(i_data_bus[716]), .A2(n9704), .B1(
        i_data_bus[844]), .B2(n9693), .ZN(n8977) );
  ND4D1BWP30P140LVT U9572 ( .A1(n8980), .A2(n8979), .A3(n8978), .A4(n8977), 
        .ZN(n8981) );
  NR4D0BWP30P140LVT U9573 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), 
        .ZN(n8985) );
  ND4D4BWP30P140LVT U9574 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), 
        .ZN(o_data_bus[12]) );
  AOI22D1BWP30P140LVT U9575 ( .A1(i_data_bus[966]), .A2(n9678), .B1(
        i_data_bus[198]), .B2(n9679), .ZN(n9009) );
  AOI22D1BWP30P140LVT U9576 ( .A1(i_data_bus[934]), .A2(n9669), .B1(
        i_data_bus[166]), .B2(n9675), .ZN(n9008) );
  AOI22D1BWP30P140LVT U9577 ( .A1(i_data_bus[774]), .A2(n9673), .B1(
        i_data_bus[294]), .B2(n9655), .ZN(n9007) );
  AOI22D1BWP30P140LVT U9578 ( .A1(i_data_bus[998]), .A2(n9677), .B1(
        i_data_bus[230]), .B2(n9671), .ZN(n8992) );
  AOI22D1BWP30P140LVT U9579 ( .A1(i_data_bus[102]), .A2(n9680), .B1(
        i_data_bus[134]), .B2(n9681), .ZN(n8991) );
  AOI22D1BWP30P140LVT U9580 ( .A1(i_data_bus[6]), .A2(n9676), .B1(
        i_data_bus[70]), .B2(n9672), .ZN(n8990) );
  AOI22D1BWP30P140LVT U9581 ( .A1(i_data_bus[38]), .A2(n9670), .B1(
        i_data_bus[902]), .B2(n9682), .ZN(n8989) );
  ND4D1BWP30P140LVT U9582 ( .A1(n8992), .A2(n8991), .A3(n8990), .A4(n8989), 
        .ZN(n9005) );
  MOAI22D1BWP30P140LVT U9583 ( .A1(n8993), .A2(n9626), .B1(i_data_bus[422]), 
        .B2(n9709), .ZN(n9004) );
  AOI22D1BWP30P140LVT U9584 ( .A1(i_data_bus[646]), .A2(n9707), .B1(
        i_data_bus[454]), .B2(n9703), .ZN(n8997) );
  AOI22D1BWP30P140LVT U9585 ( .A1(i_data_bus[806]), .A2(n9674), .B1(
        i_data_bus[870]), .B2(n9710), .ZN(n8996) );
  AOI22D1BWP30P140LVT U9586 ( .A1(i_data_bus[550]), .A2(n9695), .B1(
        i_data_bus[518]), .B2(n9698), .ZN(n8995) );
  AOI22D1BWP30P140LVT U9587 ( .A1(i_data_bus[582]), .A2(n9697), .B1(
        i_data_bus[614]), .B2(n9696), .ZN(n8994) );
  ND4D1BWP30P140LVT U9588 ( .A1(n8997), .A2(n8996), .A3(n8995), .A4(n8994), 
        .ZN(n9003) );
  AOI22D1BWP30P140LVT U9589 ( .A1(i_data_bus[838]), .A2(n9693), .B1(
        i_data_bus[710]), .B2(n9704), .ZN(n9001) );
  AOI22D1BWP30P140LVT U9590 ( .A1(i_data_bus[486]), .A2(n9656), .B1(
        i_data_bus[678]), .B2(n9705), .ZN(n9000) );
  AOI22D1BWP30P140LVT U9591 ( .A1(i_data_bus[742]), .A2(n9706), .B1(
        i_data_bus[262]), .B2(n9694), .ZN(n8999) );
  AOI22D1BWP30P140LVT U9592 ( .A1(i_data_bus[358]), .A2(n9691), .B1(
        i_data_bus[326]), .B2(n9692), .ZN(n8998) );
  ND4D1BWP30P140LVT U9593 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), 
        .ZN(n9002) );
  NR4D0BWP30P140LVT U9594 ( .A1(n9005), .A2(n9004), .A3(n9003), .A4(n9002), 
        .ZN(n9006) );
  ND4D4BWP30P140LVT U9595 ( .A1(n9009), .A2(n9008), .A3(n9007), .A4(n9006), 
        .ZN(o_data_bus[6]) );
  AOI22D1BWP30P140LVT U9596 ( .A1(i_data_bus[37]), .A2(n9670), .B1(
        i_data_bus[997]), .B2(n9677), .ZN(n9029) );
  AOI22D1BWP30P140LVT U9597 ( .A1(i_data_bus[901]), .A2(n9682), .B1(
        i_data_bus[229]), .B2(n9671), .ZN(n9028) );
  AOI22D1BWP30P140LVT U9598 ( .A1(i_data_bus[485]), .A2(n9656), .B1(
        i_data_bus[261]), .B2(n9694), .ZN(n9027) );
  AOI22D1BWP30P140LVT U9599 ( .A1(i_data_bus[101]), .A2(n9680), .B1(
        i_data_bus[69]), .B2(n9672), .ZN(n9013) );
  AOI22D1BWP30P140LVT U9600 ( .A1(i_data_bus[5]), .A2(n9676), .B1(
        i_data_bus[133]), .B2(n9681), .ZN(n9012) );
  AOI22D1BWP30P140LVT U9601 ( .A1(i_data_bus[933]), .A2(n9669), .B1(
        i_data_bus[965]), .B2(n9678), .ZN(n9011) );
  AOI22D1BWP30P140LVT U9602 ( .A1(i_data_bus[197]), .A2(n9679), .B1(
        i_data_bus[165]), .B2(n9675), .ZN(n9010) );
  ND4D1BWP30P140LVT U9603 ( .A1(n9013), .A2(n9012), .A3(n9011), .A4(n9010), 
        .ZN(n9025) );
  MOAI22D1BWP30P140LVT U9604 ( .A1(n9333), .A2(n9687), .B1(i_data_bus[741]), 
        .B2(n9706), .ZN(n9024) );
  AOI22D1BWP30P140LVT U9605 ( .A1(i_data_bus[645]), .A2(n9707), .B1(
        i_data_bus[325]), .B2(n9692), .ZN(n9017) );
  AOI22D1BWP30P140LVT U9606 ( .A1(i_data_bus[773]), .A2(n9673), .B1(
        i_data_bus[421]), .B2(n9709), .ZN(n9016) );
  AOI22D1BWP30P140LVT U9607 ( .A1(i_data_bus[549]), .A2(n9695), .B1(
        i_data_bus[581]), .B2(n9697), .ZN(n9015) );
  AOI22D1BWP30P140LVT U9608 ( .A1(i_data_bus[517]), .A2(n9698), .B1(
        i_data_bus[613]), .B2(n9696), .ZN(n9014) );
  ND4D1BWP30P140LVT U9609 ( .A1(n9017), .A2(n9016), .A3(n9015), .A4(n9014), 
        .ZN(n9023) );
  AOI22D1BWP30P140LVT U9610 ( .A1(i_data_bus[453]), .A2(n9703), .B1(
        i_data_bus[357]), .B2(n9691), .ZN(n9021) );
  AOI22D1BWP30P140LVT U9611 ( .A1(i_data_bus[837]), .A2(n9693), .B1(
        i_data_bus[869]), .B2(n9710), .ZN(n9020) );
  AOI22D1BWP30P140LVT U9612 ( .A1(i_data_bus[677]), .A2(n9705), .B1(
        i_data_bus[805]), .B2(n9674), .ZN(n9019) );
  AOI22D1BWP30P140LVT U9613 ( .A1(i_data_bus[709]), .A2(n9704), .B1(
        i_data_bus[389]), .B2(n9708), .ZN(n9018) );
  ND4D1BWP30P140LVT U9614 ( .A1(n9021), .A2(n9020), .A3(n9019), .A4(n9018), 
        .ZN(n9022) );
  NR4D0BWP30P140LVT U9615 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), 
        .ZN(n9026) );
  ND4D4BWP30P140LVT U9616 ( .A1(n9029), .A2(n9028), .A3(n9027), .A4(n9026), 
        .ZN(o_data_bus[5]) );
  AOI22D1BWP30P140LVT U9617 ( .A1(i_data_bus[99]), .A2(n9680), .B1(
        i_data_bus[963]), .B2(n9678), .ZN(n9049) );
  AOI22D1BWP30P140LVT U9618 ( .A1(i_data_bus[899]), .A2(n9682), .B1(
        i_data_bus[35]), .B2(n9670), .ZN(n9048) );
  AOI22D1BWP30P140LVT U9619 ( .A1(i_data_bus[771]), .A2(n9673), .B1(
        i_data_bus[739]), .B2(n9706), .ZN(n9047) );
  AOI22D1BWP30P140LVT U9620 ( .A1(i_data_bus[643]), .A2(n9707), .B1(
        i_data_bus[867]), .B2(n9710), .ZN(n9045) );
  AOI22D1BWP30P140LVT U9621 ( .A1(i_data_bus[931]), .A2(n9669), .B1(
        i_data_bus[227]), .B2(n9671), .ZN(n9033) );
  AOI22D1BWP30P140LVT U9622 ( .A1(i_data_bus[995]), .A2(n9677), .B1(
        i_data_bus[163]), .B2(n9675), .ZN(n9032) );
  AOI22D1BWP30P140LVT U9623 ( .A1(i_data_bus[67]), .A2(n9672), .B1(
        i_data_bus[3]), .B2(n9676), .ZN(n9031) );
  AOI22D1BWP30P140LVT U9624 ( .A1(i_data_bus[131]), .A2(n9681), .B1(
        i_data_bus[195]), .B2(n9679), .ZN(n9030) );
  ND4D1BWP30P140LVT U9625 ( .A1(n9033), .A2(n9032), .A3(n9031), .A4(n9030), 
        .ZN(n9044) );
  AOI22D1BWP30P140LVT U9626 ( .A1(i_data_bus[835]), .A2(n9693), .B1(
        i_data_bus[323]), .B2(n9692), .ZN(n9037) );
  AOI22D1BWP30P140LVT U9627 ( .A1(i_data_bus[387]), .A2(n9708), .B1(
        i_data_bus[675]), .B2(n9705), .ZN(n9036) );
  AOI22D1BWP30P140LVT U9628 ( .A1(i_data_bus[547]), .A2(n9695), .B1(
        i_data_bus[611]), .B2(n9696), .ZN(n9035) );
  AOI22D1BWP30P140LVT U9629 ( .A1(i_data_bus[515]), .A2(n9698), .B1(
        i_data_bus[579]), .B2(n9697), .ZN(n9034) );
  ND4D1BWP30P140LVT U9630 ( .A1(n9037), .A2(n9036), .A3(n9035), .A4(n9034), 
        .ZN(n9043) );
  AOI22D1BWP30P140LVT U9631 ( .A1(i_data_bus[419]), .A2(n9709), .B1(
        i_data_bus[291]), .B2(n9655), .ZN(n9041) );
  AOI22D1BWP30P140LVT U9632 ( .A1(i_data_bus[707]), .A2(n9704), .B1(
        i_data_bus[451]), .B2(n9703), .ZN(n9040) );
  AOI22D1BWP30P140LVT U9633 ( .A1(i_data_bus[355]), .A2(n9691), .B1(
        i_data_bus[259]), .B2(n9694), .ZN(n9039) );
  AOI22D1BWP30P140LVT U9634 ( .A1(i_data_bus[483]), .A2(n9656), .B1(
        i_data_bus[803]), .B2(n9674), .ZN(n9038) );
  ND4D1BWP30P140LVT U9635 ( .A1(n9041), .A2(n9040), .A3(n9039), .A4(n9038), 
        .ZN(n9042) );
  INR4D0BWP30P140LVT U9636 ( .A1(n9045), .B1(n9044), .B2(n9043), .B3(n9042), 
        .ZN(n9046) );
  ND4D4BWP30P140LVT U9637 ( .A1(n9049), .A2(n9048), .A3(n9047), .A4(n9046), 
        .ZN(o_data_bus[3]) );
  AOI22D1BWP30P140LVT U9638 ( .A1(i_data_bus[97]), .A2(n9680), .B1(
        i_data_bus[225]), .B2(n9671), .ZN(n9070) );
  AOI22D1BWP30P140LVT U9639 ( .A1(i_data_bus[65]), .A2(n9672), .B1(
        i_data_bus[193]), .B2(n9679), .ZN(n9069) );
  AOI22D1BWP30P140LVT U9640 ( .A1(i_data_bus[769]), .A2(n9673), .B1(
        i_data_bus[801]), .B2(n9674), .ZN(n9068) );
  AOI22D1BWP30P140LVT U9641 ( .A1(i_data_bus[961]), .A2(n9678), .B1(
        i_data_bus[993]), .B2(n9677), .ZN(n9053) );
  AOI22D1BWP30P140LVT U9642 ( .A1(i_data_bus[33]), .A2(n9670), .B1(
        i_data_bus[1]), .B2(n9676), .ZN(n9052) );
  AOI22D1BWP30P140LVT U9643 ( .A1(i_data_bus[897]), .A2(n9682), .B1(
        i_data_bus[929]), .B2(n9669), .ZN(n9051) );
  AOI22D1BWP30P140LVT U9644 ( .A1(i_data_bus[161]), .A2(n9675), .B1(
        i_data_bus[129]), .B2(n9681), .ZN(n9050) );
  ND4D1BWP30P140LVT U9645 ( .A1(n9053), .A2(n9052), .A3(n9051), .A4(n9050), 
        .ZN(n9066) );
  MOAI22D1BWP30P140LVT U9646 ( .A1(n9054), .A2(n9181), .B1(i_data_bus[865]), 
        .B2(n9710), .ZN(n9065) );
  AOI22D1BWP30P140LVT U9647 ( .A1(i_data_bus[705]), .A2(n9704), .B1(
        i_data_bus[321]), .B2(n9692), .ZN(n9058) );
  AOI22D1BWP30P140LVT U9648 ( .A1(i_data_bus[353]), .A2(n9691), .B1(
        i_data_bus[833]), .B2(n9693), .ZN(n9057) );
  AOI22D1BWP30P140LVT U9649 ( .A1(i_data_bus[577]), .A2(n9697), .B1(
        i_data_bus[545]), .B2(n9695), .ZN(n9056) );
  AOI22D1BWP30P140LVT U9650 ( .A1(i_data_bus[609]), .A2(n9696), .B1(
        i_data_bus[513]), .B2(n9698), .ZN(n9055) );
  ND4D1BWP30P140LVT U9651 ( .A1(n9058), .A2(n9057), .A3(n9056), .A4(n9055), 
        .ZN(n9064) );
  AOI22D1BWP30P140LVT U9652 ( .A1(i_data_bus[673]), .A2(n9705), .B1(
        i_data_bus[417]), .B2(n9709), .ZN(n9062) );
  AOI22D1BWP30P140LVT U9653 ( .A1(i_data_bus[449]), .A2(n9703), .B1(
        i_data_bus[289]), .B2(n9655), .ZN(n9061) );
  AOI22D1BWP30P140LVT U9654 ( .A1(i_data_bus[481]), .A2(n9656), .B1(
        i_data_bus[737]), .B2(n9706), .ZN(n9060) );
  AOI22D1BWP30P140LVT U9655 ( .A1(i_data_bus[385]), .A2(n9708), .B1(
        i_data_bus[641]), .B2(n9707), .ZN(n9059) );
  ND4D1BWP30P140LVT U9656 ( .A1(n9062), .A2(n9061), .A3(n9060), .A4(n9059), 
        .ZN(n9063) );
  NR4D0BWP30P140LVT U9657 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), 
        .ZN(n9067) );
  ND4D4BWP30P140LVT U9658 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), 
        .ZN(o_data_bus[1]) );
  AOI22D1BWP30P140LVT U9659 ( .A1(i_data_bus[822]), .A2(n9552), .B1(
        i_data_bus[662]), .B2(n9558), .ZN(n9091) );
  AOI22D1BWP30P140LVT U9660 ( .A1(i_data_bus[54]), .A2(n9548), .B1(
        i_data_bus[118]), .B2(n9555), .ZN(n9090) );
  AOI22D1BWP30P140LVT U9661 ( .A1(i_data_bus[182]), .A2(n9583), .B1(
        i_data_bus[470]), .B2(n9582), .ZN(n9089) );
  AOI22D1BWP30P140LVT U9662 ( .A1(i_data_bus[86]), .A2(n9549), .B1(
        i_data_bus[726]), .B2(n9554), .ZN(n9074) );
  AOI22D1BWP30P140LVT U9663 ( .A1(i_data_bus[22]), .A2(n9553), .B1(
        i_data_bus[790]), .B2(n9547), .ZN(n9073) );
  AOI22D1BWP30P140LVT U9664 ( .A1(i_data_bus[886]), .A2(n9556), .B1(
        i_data_bus[854]), .B2(n9557), .ZN(n9072) );
  AOI22D1BWP30P140LVT U9665 ( .A1(i_data_bus[694]), .A2(n9559), .B1(
        i_data_bus[758]), .B2(n9546), .ZN(n9071) );
  ND4D1BWP30P140LVT U9666 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), 
        .ZN(n9087) );
  MOAI22D1BWP30P140LVT U9667 ( .A1(n9075), .A2(n9483), .B1(i_data_bus[246]), 
        .B2(n9568), .ZN(n9086) );
  AOI22D1BWP30P140LVT U9668 ( .A1(i_data_bus[502]), .A2(n9580), .B1(
        i_data_bus[310]), .B2(n9584), .ZN(n9079) );
  AOI22D1BWP30P140LVT U9669 ( .A1(i_data_bus[1014]), .A2(n9571), .B1(
        i_data_bus[342]), .B2(n9570), .ZN(n9078) );
  AOI22D1BWP30P140LVT U9670 ( .A1(i_data_bus[534]), .A2(n9573), .B1(
        i_data_bus[630]), .B2(n9574), .ZN(n9077) );
  AOI22D1BWP30P140LVT U9671 ( .A1(i_data_bus[566]), .A2(n9575), .B1(
        i_data_bus[598]), .B2(n9572), .ZN(n9076) );
  ND4D1BWP30P140LVT U9672 ( .A1(n9079), .A2(n9078), .A3(n9077), .A4(n9076), 
        .ZN(n9085) );
  AOI22D1BWP30P140LVT U9673 ( .A1(i_data_bus[950]), .A2(n9587), .B1(
        i_data_bus[374]), .B2(n9569), .ZN(n9083) );
  AOI22D1BWP30P140LVT U9674 ( .A1(i_data_bus[150]), .A2(n9533), .B1(
        i_data_bus[278]), .B2(n9586), .ZN(n9082) );
  AOI22D1BWP30P140LVT U9675 ( .A1(i_data_bus[918]), .A2(n9581), .B1(
        i_data_bus[438]), .B2(n9532), .ZN(n9081) );
  AOI22D1BWP30P140LVT U9676 ( .A1(i_data_bus[982]), .A2(n9551), .B1(
        i_data_bus[406]), .B2(n9585), .ZN(n9080) );
  ND4D1BWP30P140LVT U9677 ( .A1(n9083), .A2(n9082), .A3(n9081), .A4(n9080), 
        .ZN(n9084) );
  NR4D0BWP30P140LVT U9678 ( .A1(n9087), .A2(n9086), .A3(n9085), .A4(n9084), 
        .ZN(n9088) );
  ND4D4BWP30P140LVT U9679 ( .A1(n9091), .A2(n9090), .A3(n9089), .A4(n9088), 
        .ZN(o_data_bus[246]) );
  AOI22D1BWP30P140LVT U9680 ( .A1(i_data_bus[910]), .A2(n9682), .B1(
        i_data_bus[14]), .B2(n9676), .ZN(n9111) );
  AOI22D1BWP30P140LVT U9681 ( .A1(i_data_bus[974]), .A2(n9678), .B1(
        i_data_bus[142]), .B2(n9681), .ZN(n9110) );
  AOI22D1BWP30P140LVT U9682 ( .A1(i_data_bus[462]), .A2(n9703), .B1(
        i_data_bus[398]), .B2(n9708), .ZN(n9109) );
  AOI22D1BWP30P140LVT U9683 ( .A1(i_data_bus[334]), .A2(n9692), .B1(
        i_data_bus[878]), .B2(n9710), .ZN(n9107) );
  AOI22D1BWP30P140LVT U9684 ( .A1(i_data_bus[1006]), .A2(n9677), .B1(
        i_data_bus[942]), .B2(n9669), .ZN(n9095) );
  AOI22D1BWP30P140LVT U9685 ( .A1(i_data_bus[46]), .A2(n9670), .B1(
        i_data_bus[206]), .B2(n9679), .ZN(n9094) );
  AOI22D1BWP30P140LVT U9686 ( .A1(i_data_bus[78]), .A2(n9672), .B1(
        i_data_bus[174]), .B2(n9675), .ZN(n9093) );
  AOI22D1BWP30P140LVT U9687 ( .A1(i_data_bus[110]), .A2(n9680), .B1(
        i_data_bus[238]), .B2(n9671), .ZN(n9092) );
  ND4D1BWP30P140LVT U9688 ( .A1(n9095), .A2(n9094), .A3(n9093), .A4(n9092), 
        .ZN(n9106) );
  AOI22D1BWP30P140LVT U9689 ( .A1(i_data_bus[846]), .A2(n9693), .B1(
        i_data_bus[302]), .B2(n9655), .ZN(n9099) );
  AOI22D1BWP30P140LVT U9690 ( .A1(i_data_bus[270]), .A2(n9694), .B1(
        i_data_bus[814]), .B2(n9674), .ZN(n9098) );
  AOI22D1BWP30P140LVT U9691 ( .A1(i_data_bus[558]), .A2(n9695), .B1(
        i_data_bus[622]), .B2(n9696), .ZN(n9097) );
  AOI22D1BWP30P140LVT U9692 ( .A1(i_data_bus[590]), .A2(n9697), .B1(
        i_data_bus[526]), .B2(n9698), .ZN(n9096) );
  ND4D1BWP30P140LVT U9693 ( .A1(n9099), .A2(n9098), .A3(n9097), .A4(n9096), 
        .ZN(n9105) );
  AOI22D1BWP30P140LVT U9694 ( .A1(i_data_bus[686]), .A2(n9705), .B1(
        i_data_bus[718]), .B2(n9704), .ZN(n9103) );
  AOI22D1BWP30P140LVT U9695 ( .A1(i_data_bus[782]), .A2(n9673), .B1(
        i_data_bus[430]), .B2(n9709), .ZN(n9102) );
  AOI22D1BWP30P140LVT U9696 ( .A1(i_data_bus[366]), .A2(n9691), .B1(
        i_data_bus[494]), .B2(n9656), .ZN(n9101) );
  AOI22D1BWP30P140LVT U9697 ( .A1(i_data_bus[750]), .A2(n9706), .B1(
        i_data_bus[654]), .B2(n9707), .ZN(n9100) );
  ND4D1BWP30P140LVT U9698 ( .A1(n9103), .A2(n9102), .A3(n9101), .A4(n9100), 
        .ZN(n9104) );
  INR4D0BWP30P140LVT U9699 ( .A1(n9107), .B1(n9106), .B2(n9105), .B3(n9104), 
        .ZN(n9108) );
  ND4D4BWP30P140LVT U9700 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), 
        .ZN(o_data_bus[14]) );
  AOI22D1BWP30P140LVT U9701 ( .A1(i_data_bus[932]), .A2(n9669), .B1(
        i_data_bus[132]), .B2(n9681), .ZN(n9132) );
  AOI22D1BWP30P140LVT U9702 ( .A1(i_data_bus[36]), .A2(n9670), .B1(
        i_data_bus[196]), .B2(n9679), .ZN(n9131) );
  AOI22D1BWP30P140LVT U9703 ( .A1(i_data_bus[452]), .A2(n9703), .B1(
        i_data_bus[484]), .B2(n9656), .ZN(n9130) );
  AOI22D1BWP30P140LVT U9704 ( .A1(i_data_bus[964]), .A2(n9678), .B1(
        i_data_bus[996]), .B2(n9677), .ZN(n9115) );
  AOI22D1BWP30P140LVT U9705 ( .A1(i_data_bus[4]), .A2(n9676), .B1(
        i_data_bus[228]), .B2(n9671), .ZN(n9114) );
  AOI22D1BWP30P140LVT U9706 ( .A1(i_data_bus[100]), .A2(n9680), .B1(
        i_data_bus[164]), .B2(n9675), .ZN(n9113) );
  AOI22D1BWP30P140LVT U9707 ( .A1(i_data_bus[900]), .A2(n9682), .B1(
        i_data_bus[68]), .B2(n9672), .ZN(n9112) );
  ND4D1BWP30P140LVT U9708 ( .A1(n9115), .A2(n9114), .A3(n9113), .A4(n9112), 
        .ZN(n9128) );
  MOAI22D1BWP30P140LVT U9709 ( .A1(n9116), .A2(n9137), .B1(i_data_bus[676]), 
        .B2(n9705), .ZN(n9127) );
  AOI22D1BWP30P140LVT U9710 ( .A1(i_data_bus[708]), .A2(n9704), .B1(
        i_data_bus[420]), .B2(n9709), .ZN(n9120) );
  AOI22D1BWP30P140LVT U9711 ( .A1(i_data_bus[740]), .A2(n9706), .B1(
        i_data_bus[772]), .B2(n9673), .ZN(n9119) );
  AOI22D1BWP30P140LVT U9712 ( .A1(i_data_bus[548]), .A2(n9695), .B1(
        i_data_bus[516]), .B2(n9698), .ZN(n9118) );
  AOI22D1BWP30P140LVT U9713 ( .A1(i_data_bus[612]), .A2(n9696), .B1(
        i_data_bus[580]), .B2(n9697), .ZN(n9117) );
  ND4D1BWP30P140LVT U9714 ( .A1(n9120), .A2(n9119), .A3(n9118), .A4(n9117), 
        .ZN(n9126) );
  AOI22D1BWP30P140LVT U9715 ( .A1(i_data_bus[868]), .A2(n9710), .B1(
        i_data_bus[292]), .B2(n9655), .ZN(n9124) );
  AOI22D1BWP30P140LVT U9716 ( .A1(i_data_bus[260]), .A2(n9694), .B1(
        i_data_bus[388]), .B2(n9708), .ZN(n9123) );
  AOI22D1BWP30P140LVT U9717 ( .A1(i_data_bus[836]), .A2(n9693), .B1(
        i_data_bus[804]), .B2(n9674), .ZN(n9122) );
  AOI22D1BWP30P140LVT U9718 ( .A1(i_data_bus[644]), .A2(n9707), .B1(
        i_data_bus[356]), .B2(n9691), .ZN(n9121) );
  ND4D1BWP30P140LVT U9719 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), 
        .ZN(n9125) );
  NR4D0BWP30P140LVT U9720 ( .A1(n9128), .A2(n9127), .A3(n9126), .A4(n9125), 
        .ZN(n9129) );
  ND4D4BWP30P140LVT U9721 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), 
        .ZN(o_data_bus[4]) );
  AOI22D1BWP30P140LVT U9722 ( .A1(i_data_bus[962]), .A2(n9678), .B1(
        i_data_bus[994]), .B2(n9677), .ZN(n9155) );
  AOI22D1BWP30P140LVT U9723 ( .A1(i_data_bus[2]), .A2(n9676), .B1(
        i_data_bus[930]), .B2(n9669), .ZN(n9154) );
  AOI22D1BWP30P140LVT U9724 ( .A1(i_data_bus[450]), .A2(n9703), .B1(
        i_data_bus[770]), .B2(n9673), .ZN(n9153) );
  AOI22D1BWP30P140LVT U9725 ( .A1(i_data_bus[98]), .A2(n9680), .B1(
        i_data_bus[130]), .B2(n9681), .ZN(n9136) );
  AOI22D1BWP30P140LVT U9726 ( .A1(i_data_bus[66]), .A2(n9672), .B1(
        i_data_bus[898]), .B2(n9682), .ZN(n9135) );
  AOI22D1BWP30P140LVT U9727 ( .A1(i_data_bus[34]), .A2(n9670), .B1(
        i_data_bus[194]), .B2(n9679), .ZN(n9134) );
  AOI22D1BWP30P140LVT U9728 ( .A1(i_data_bus[162]), .A2(n9675), .B1(
        i_data_bus[226]), .B2(n9671), .ZN(n9133) );
  ND4D1BWP30P140LVT U9729 ( .A1(n9136), .A2(n9135), .A3(n9134), .A4(n9133), 
        .ZN(n9151) );
  OAI22D1BWP30P140LVT U9730 ( .A1(n9139), .A2(n9181), .B1(n9138), .B2(n9137), 
        .ZN(n9150) );
  AOI22D1BWP30P140LVT U9731 ( .A1(i_data_bus[802]), .A2(n9674), .B1(
        i_data_bus[738]), .B2(n9706), .ZN(n9143) );
  AOI22D1BWP30P140LVT U9732 ( .A1(i_data_bus[482]), .A2(n9656), .B1(
        i_data_bus[706]), .B2(n9704), .ZN(n9142) );
  AOI22D1BWP30P140LVT U9733 ( .A1(i_data_bus[578]), .A2(n9697), .B1(
        i_data_bus[546]), .B2(n9695), .ZN(n9141) );
  AOI22D1BWP30P140LVT U9734 ( .A1(i_data_bus[514]), .A2(n9698), .B1(
        i_data_bus[610]), .B2(n9696), .ZN(n9140) );
  ND4D1BWP30P140LVT U9735 ( .A1(n9143), .A2(n9142), .A3(n9141), .A4(n9140), 
        .ZN(n9149) );
  AOI22D1BWP30P140LVT U9736 ( .A1(i_data_bus[418]), .A2(n9709), .B1(
        i_data_bus[354]), .B2(n9691), .ZN(n9147) );
  AOI22D1BWP30P140LVT U9737 ( .A1(i_data_bus[674]), .A2(n9705), .B1(
        i_data_bus[834]), .B2(n9693), .ZN(n9146) );
  AOI22D1BWP30P140LVT U9738 ( .A1(i_data_bus[866]), .A2(n9710), .B1(
        i_data_bus[386]), .B2(n9708), .ZN(n9145) );
  AOI22D1BWP30P140LVT U9739 ( .A1(i_data_bus[290]), .A2(n9655), .B1(
        i_data_bus[642]), .B2(n9707), .ZN(n9144) );
  ND4D1BWP30P140LVT U9740 ( .A1(n9147), .A2(n9146), .A3(n9145), .A4(n9144), 
        .ZN(n9148) );
  NR4D0BWP30P140LVT U9741 ( .A1(n9151), .A2(n9150), .A3(n9149), .A4(n9148), 
        .ZN(n9152) );
  ND4D4BWP30P140LVT U9742 ( .A1(n9155), .A2(n9154), .A3(n9153), .A4(n9152), 
        .ZN(o_data_bus[2]) );
  AOI22D1BWP30P140LVT U9743 ( .A1(i_data_bus[658]), .A2(n9558), .B1(
        i_data_bus[754]), .B2(n9546), .ZN(n9176) );
  AOI22D1BWP30P140LVT U9744 ( .A1(i_data_bus[722]), .A2(n9554), .B1(
        i_data_bus[818]), .B2(n9552), .ZN(n9175) );
  AOI22D1BWP30P140LVT U9745 ( .A1(i_data_bus[178]), .A2(n9583), .B1(
        i_data_bus[306]), .B2(n9584), .ZN(n9174) );
  AOI22D1BWP30P140LVT U9746 ( .A1(i_data_bus[82]), .A2(n9549), .B1(
        i_data_bus[882]), .B2(n9556), .ZN(n9159) );
  AOI22D1BWP30P140LVT U9747 ( .A1(i_data_bus[690]), .A2(n9559), .B1(
        i_data_bus[850]), .B2(n9557), .ZN(n9158) );
  AOI22D1BWP30P140LVT U9748 ( .A1(i_data_bus[50]), .A2(n9548), .B1(
        i_data_bus[786]), .B2(n9547), .ZN(n9157) );
  AOI22D1BWP30P140LVT U9749 ( .A1(i_data_bus[114]), .A2(n9555), .B1(
        i_data_bus[18]), .B2(n9553), .ZN(n9156) );
  ND4D1BWP30P140LVT U9750 ( .A1(n9159), .A2(n9158), .A3(n9157), .A4(n9156), 
        .ZN(n9172) );
  INVD1BWP30P140LVT U9751 ( .I(n9533), .ZN(n9564) );
  MOAI22D1BWP30P140LVT U9752 ( .A1(n9160), .A2(n9564), .B1(i_data_bus[978]), 
        .B2(n9551), .ZN(n9171) );
  AOI22D1BWP30P140LVT U9753 ( .A1(i_data_bus[914]), .A2(n9581), .B1(
        i_data_bus[498]), .B2(n9580), .ZN(n9164) );
  AOI22D1BWP30P140LVT U9754 ( .A1(i_data_bus[1010]), .A2(n9571), .B1(
        i_data_bus[338]), .B2(n9570), .ZN(n9163) );
  AOI22D1BWP30P140LVT U9755 ( .A1(i_data_bus[530]), .A2(n9573), .B1(
        i_data_bus[562]), .B2(n9575), .ZN(n9162) );
  AOI22D1BWP30P140LVT U9756 ( .A1(i_data_bus[626]), .A2(n9574), .B1(
        i_data_bus[594]), .B2(n9572), .ZN(n9161) );
  ND4D1BWP30P140LVT U9757 ( .A1(n9164), .A2(n9163), .A3(n9162), .A4(n9161), 
        .ZN(n9170) );
  AOI22D1BWP30P140LVT U9758 ( .A1(i_data_bus[946]), .A2(n9587), .B1(
        i_data_bus[274]), .B2(n9586), .ZN(n9168) );
  AOI22D1BWP30P140LVT U9759 ( .A1(i_data_bus[402]), .A2(n9585), .B1(
        i_data_bus[210]), .B2(n9550), .ZN(n9167) );
  AOI22D1BWP30P140LVT U9760 ( .A1(i_data_bus[370]), .A2(n9569), .B1(
        i_data_bus[466]), .B2(n9582), .ZN(n9166) );
  AOI22D1BWP30P140LVT U9761 ( .A1(i_data_bus[242]), .A2(n9568), .B1(
        i_data_bus[434]), .B2(n9532), .ZN(n9165) );
  ND4D1BWP30P140LVT U9762 ( .A1(n9168), .A2(n9167), .A3(n9166), .A4(n9165), 
        .ZN(n9169) );
  NR4D0BWP30P140LVT U9763 ( .A1(n9172), .A2(n9171), .A3(n9170), .A4(n9169), 
        .ZN(n9173) );
  ND4D4BWP30P140LVT U9764 ( .A1(n9176), .A2(n9175), .A3(n9174), .A4(n9173), 
        .ZN(o_data_bus[242]) );
  AOI22D1BWP30P140LVT U9765 ( .A1(i_data_bus[992]), .A2(n9677), .B1(
        i_data_bus[32]), .B2(n9670), .ZN(n9198) );
  AOI22D1BWP30P140LVT U9766 ( .A1(i_data_bus[160]), .A2(n9675), .B1(
        i_data_bus[128]), .B2(n9681), .ZN(n9197) );
  AOI22D1BWP30P140LVT U9767 ( .A1(i_data_bus[480]), .A2(n9656), .B1(
        i_data_bus[448]), .B2(n9703), .ZN(n9196) );
  AOI22D1BWP30P140LVT U9768 ( .A1(i_data_bus[960]), .A2(n9678), .B1(
        i_data_bus[192]), .B2(n9679), .ZN(n9180) );
  AOI22D1BWP30P140LVT U9769 ( .A1(i_data_bus[96]), .A2(n9680), .B1(
        i_data_bus[224]), .B2(n9671), .ZN(n9179) );
  AOI22D1BWP30P140LVT U9770 ( .A1(i_data_bus[64]), .A2(n9672), .B1(
        i_data_bus[896]), .B2(n9682), .ZN(n9178) );
  AOI22D1BWP30P140LVT U9771 ( .A1(i_data_bus[928]), .A2(n9669), .B1(
        i_data_bus[0]), .B2(n9676), .ZN(n9177) );
  ND4D1BWP30P140LVT U9772 ( .A1(n9180), .A2(n9179), .A3(n9178), .A4(n9177), 
        .ZN(n9194) );
  MOAI22D1BWP30P140LVT U9773 ( .A1(n9182), .A2(n9181), .B1(i_data_bus[640]), 
        .B2(n9707), .ZN(n9193) );
  AOI22D1BWP30P140LVT U9774 ( .A1(i_data_bus[800]), .A2(n9674), .B1(
        i_data_bus[320]), .B2(n9692), .ZN(n9186) );
  AOI22D1BWP30P140LVT U9775 ( .A1(i_data_bus[384]), .A2(n9708), .B1(
        i_data_bus[768]), .B2(n9673), .ZN(n9185) );
  AOI22D1BWP30P140LVT U9776 ( .A1(i_data_bus[512]), .A2(n9698), .B1(
        i_data_bus[608]), .B2(n9696), .ZN(n9184) );
  AOI22D1BWP30P140LVT U9777 ( .A1(i_data_bus[544]), .A2(n9695), .B1(
        i_data_bus[576]), .B2(n9697), .ZN(n9183) );
  ND4D1BWP30P140LVT U9778 ( .A1(n9186), .A2(n9185), .A3(n9184), .A4(n9183), 
        .ZN(n9192) );
  AOI22D1BWP30P140LVT U9779 ( .A1(i_data_bus[352]), .A2(n9691), .B1(
        i_data_bus[672]), .B2(n9705), .ZN(n9190) );
  AOI22D1BWP30P140LVT U9780 ( .A1(i_data_bus[704]), .A2(n9704), .B1(
        i_data_bus[864]), .B2(n9710), .ZN(n9189) );
  AOI22D1BWP30P140LVT U9781 ( .A1(i_data_bus[416]), .A2(n9709), .B1(
        i_data_bus[288]), .B2(n9655), .ZN(n9188) );
  AOI22D1BWP30P140LVT U9782 ( .A1(i_data_bus[832]), .A2(n9693), .B1(
        i_data_bus[736]), .B2(n9706), .ZN(n9187) );
  ND4D1BWP30P140LVT U9783 ( .A1(n9190), .A2(n9189), .A3(n9188), .A4(n9187), 
        .ZN(n9191) );
  NR4D0BWP30P140LVT U9784 ( .A1(n9194), .A2(n9193), .A3(n9192), .A4(n9191), 
        .ZN(n9195) );
  ND4D4BWP30P140LVT U9785 ( .A1(n9198), .A2(n9197), .A3(n9196), .A4(n9195), 
        .ZN(o_data_bus[0]) );
  AOI22D1BWP30P140LVT U9786 ( .A1(i_data_bus[63]), .A2(n9548), .B1(
        i_data_bus[671]), .B2(n9558), .ZN(n9219) );
  AOI22D1BWP30P140LVT U9787 ( .A1(i_data_bus[767]), .A2(n9546), .B1(
        i_data_bus[703]), .B2(n9559), .ZN(n9218) );
  AOI22D1BWP30P140LVT U9788 ( .A1(i_data_bus[991]), .A2(n9551), .B1(
        i_data_bus[255]), .B2(n9568), .ZN(n9217) );
  AOI22D1BWP30P140LVT U9789 ( .A1(i_data_bus[95]), .A2(n9549), .B1(
        i_data_bus[127]), .B2(n9555), .ZN(n9202) );
  AOI22D1BWP30P140LVT U9790 ( .A1(i_data_bus[799]), .A2(n9547), .B1(
        i_data_bus[863]), .B2(n9557), .ZN(n9201) );
  AOI22D1BWP30P140LVT U9791 ( .A1(i_data_bus[735]), .A2(n9554), .B1(
        i_data_bus[831]), .B2(n9552), .ZN(n9200) );
  AOI22D1BWP30P140LVT U9792 ( .A1(i_data_bus[31]), .A2(n9553), .B1(
        i_data_bus[895]), .B2(n9556), .ZN(n9199) );
  ND4D1BWP30P140LVT U9793 ( .A1(n9202), .A2(n9201), .A3(n9200), .A4(n9199), 
        .ZN(n9215) );
  MOAI22D1BWP30P140LVT U9794 ( .A1(n9203), .A2(n9419), .B1(i_data_bus[511]), 
        .B2(n9580), .ZN(n9214) );
  AOI22D1BWP30P140LVT U9795 ( .A1(i_data_bus[1023]), .A2(n9571), .B1(
        i_data_bus[287]), .B2(n9586), .ZN(n9207) );
  AOI22D1BWP30P140LVT U9796 ( .A1(i_data_bus[927]), .A2(n9581), .B1(
        i_data_bus[351]), .B2(n9570), .ZN(n9206) );
  AOI22D1BWP30P140LVT U9797 ( .A1(i_data_bus[575]), .A2(n9575), .B1(
        i_data_bus[607]), .B2(n9572), .ZN(n9205) );
  AOI22D1BWP30P140LVT U9798 ( .A1(i_data_bus[639]), .A2(n9574), .B1(
        i_data_bus[543]), .B2(n9573), .ZN(n9204) );
  ND4D1BWP30P140LVT U9799 ( .A1(n9207), .A2(n9206), .A3(n9205), .A4(n9204), 
        .ZN(n9213) );
  AOI22D1BWP30P140LVT U9800 ( .A1(i_data_bus[447]), .A2(n9532), .B1(
        i_data_bus[479]), .B2(n9582), .ZN(n9211) );
  AOI22D1BWP30P140LVT U9801 ( .A1(i_data_bus[223]), .A2(n9550), .B1(
        i_data_bus[383]), .B2(n9569), .ZN(n9210) );
  AOI22D1BWP30P140LVT U9802 ( .A1(i_data_bus[959]), .A2(n9587), .B1(
        i_data_bus[159]), .B2(n9533), .ZN(n9209) );
  AOI22D1BWP30P140LVT U9803 ( .A1(i_data_bus[319]), .A2(n9584), .B1(
        i_data_bus[415]), .B2(n9585), .ZN(n9208) );
  ND4D1BWP30P140LVT U9804 ( .A1(n9211), .A2(n9210), .A3(n9209), .A4(n9208), 
        .ZN(n9212) );
  NR4D0BWP30P140LVT U9805 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), 
        .ZN(n9216) );
  ND4D4BWP30P140LVT U9806 ( .A1(n9219), .A2(n9218), .A3(n9217), .A4(n9216), 
        .ZN(o_data_bus[255]) );
  AOI22D1BWP30P140LVT U9807 ( .A1(i_data_bus[94]), .A2(n9549), .B1(
        i_data_bus[702]), .B2(n9559), .ZN(n9240) );
  AOI22D1BWP30P140LVT U9808 ( .A1(i_data_bus[62]), .A2(n9548), .B1(
        i_data_bus[126]), .B2(n9555), .ZN(n9239) );
  AOI22D1BWP30P140LVT U9809 ( .A1(i_data_bus[958]), .A2(n9587), .B1(
        i_data_bus[478]), .B2(n9582), .ZN(n9238) );
  AOI22D1BWP30P140LVT U9810 ( .A1(i_data_bus[862]), .A2(n9557), .B1(
        i_data_bus[734]), .B2(n9554), .ZN(n9223) );
  AOI22D1BWP30P140LVT U9811 ( .A1(i_data_bus[30]), .A2(n9553), .B1(
        i_data_bus[798]), .B2(n9547), .ZN(n9222) );
  AOI22D1BWP30P140LVT U9812 ( .A1(i_data_bus[670]), .A2(n9558), .B1(
        i_data_bus[830]), .B2(n9552), .ZN(n9221) );
  AOI22D1BWP30P140LVT U9813 ( .A1(i_data_bus[766]), .A2(n9546), .B1(
        i_data_bus[894]), .B2(n9556), .ZN(n9220) );
  ND4D1BWP30P140LVT U9814 ( .A1(n9223), .A2(n9222), .A3(n9221), .A4(n9220), 
        .ZN(n9236) );
  MOAI22D1BWP30P140LVT U9815 ( .A1(n9224), .A2(n9245), .B1(i_data_bus[990]), 
        .B2(n9551), .ZN(n9235) );
  AOI22D1BWP30P140LVT U9816 ( .A1(i_data_bus[222]), .A2(n9550), .B1(
        i_data_bus[382]), .B2(n9569), .ZN(n9228) );
  AOI22D1BWP30P140LVT U9817 ( .A1(i_data_bus[1022]), .A2(n9571), .B1(
        i_data_bus[446]), .B2(n9532), .ZN(n9227) );
  AOI22D1BWP30P140LVT U9818 ( .A1(i_data_bus[542]), .A2(n9573), .B1(
        i_data_bus[606]), .B2(n9572), .ZN(n9226) );
  AOI22D1BWP30P140LVT U9819 ( .A1(i_data_bus[574]), .A2(n9575), .B1(
        i_data_bus[638]), .B2(n9574), .ZN(n9225) );
  ND4D1BWP30P140LVT U9820 ( .A1(n9228), .A2(n9227), .A3(n9226), .A4(n9225), 
        .ZN(n9234) );
  AOI22D1BWP30P140LVT U9821 ( .A1(i_data_bus[926]), .A2(n9581), .B1(
        i_data_bus[286]), .B2(n9586), .ZN(n9232) );
  AOI22D1BWP30P140LVT U9822 ( .A1(i_data_bus[318]), .A2(n9584), .B1(
        i_data_bus[190]), .B2(n9583), .ZN(n9231) );
  AOI22D1BWP30P140LVT U9823 ( .A1(i_data_bus[254]), .A2(n9568), .B1(
        i_data_bus[158]), .B2(n9533), .ZN(n9230) );
  AOI22D1BWP30P140LVT U9824 ( .A1(i_data_bus[350]), .A2(n9570), .B1(
        i_data_bus[510]), .B2(n9580), .ZN(n9229) );
  ND4D1BWP30P140LVT U9825 ( .A1(n9232), .A2(n9231), .A3(n9230), .A4(n9229), 
        .ZN(n9233) );
  NR4D0BWP30P140LVT U9826 ( .A1(n9236), .A2(n9235), .A3(n9234), .A4(n9233), 
        .ZN(n9237) );
  ND4D4BWP30P140LVT U9827 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), 
        .ZN(o_data_bus[254]) );
  AOI22D1BWP30P140LVT U9828 ( .A1(i_data_bus[124]), .A2(n9555), .B1(
        i_data_bus[860]), .B2(n9557), .ZN(n9264) );
  AOI22D1BWP30P140LVT U9829 ( .A1(i_data_bus[92]), .A2(n9549), .B1(
        i_data_bus[668]), .B2(n9558), .ZN(n9263) );
  AOI22D1BWP30P140LVT U9830 ( .A1(i_data_bus[988]), .A2(n9551), .B1(
        i_data_bus[284]), .B2(n9586), .ZN(n9262) );
  AOI22D1BWP30P140LVT U9831 ( .A1(i_data_bus[28]), .A2(n9553), .B1(
        i_data_bus[732]), .B2(n9554), .ZN(n9244) );
  AOI22D1BWP30P140LVT U9832 ( .A1(i_data_bus[828]), .A2(n9552), .B1(
        i_data_bus[700]), .B2(n9559), .ZN(n9243) );
  AOI22D1BWP30P140LVT U9833 ( .A1(i_data_bus[796]), .A2(n9547), .B1(
        i_data_bus[764]), .B2(n9546), .ZN(n9242) );
  AOI22D1BWP30P140LVT U9834 ( .A1(i_data_bus[60]), .A2(n9548), .B1(
        i_data_bus[892]), .B2(n9556), .ZN(n9241) );
  ND4D1BWP30P140LVT U9835 ( .A1(n9244), .A2(n9243), .A3(n9242), .A4(n9241), 
        .ZN(n9260) );
  OAI22D1BWP30P140LVT U9836 ( .A1(n9248), .A2(n9247), .B1(n9246), .B2(n9245), 
        .ZN(n9259) );
  AOI22D1BWP30P140LVT U9837 ( .A1(i_data_bus[924]), .A2(n9581), .B1(
        i_data_bus[444]), .B2(n9532), .ZN(n9252) );
  AOI22D1BWP30P140LVT U9838 ( .A1(i_data_bus[380]), .A2(n9569), .B1(
        i_data_bus[220]), .B2(n9550), .ZN(n9251) );
  AOI22D1BWP30P140LVT U9839 ( .A1(i_data_bus[636]), .A2(n9574), .B1(
        i_data_bus[604]), .B2(n9572), .ZN(n9250) );
  AOI22D1BWP30P140LVT U9840 ( .A1(i_data_bus[540]), .A2(n9573), .B1(
        i_data_bus[572]), .B2(n9575), .ZN(n9249) );
  ND4D1BWP30P140LVT U9841 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), 
        .ZN(n9258) );
  AOI22D1BWP30P140LVT U9842 ( .A1(i_data_bus[956]), .A2(n9587), .B1(
        i_data_bus[316]), .B2(n9584), .ZN(n9256) );
  AOI22D1BWP30P140LVT U9843 ( .A1(i_data_bus[1020]), .A2(n9571), .B1(
        i_data_bus[156]), .B2(n9533), .ZN(n9255) );
  AOI22D1BWP30P140LVT U9844 ( .A1(i_data_bus[188]), .A2(n9583), .B1(
        i_data_bus[476]), .B2(n9582), .ZN(n9254) );
  AOI22D1BWP30P140LVT U9845 ( .A1(i_data_bus[252]), .A2(n9568), .B1(
        i_data_bus[508]), .B2(n9580), .ZN(n9253) );
  ND4D1BWP30P140LVT U9846 ( .A1(n9256), .A2(n9255), .A3(n9254), .A4(n9253), 
        .ZN(n9257) );
  NR4D0BWP30P140LVT U9847 ( .A1(n9260), .A2(n9259), .A3(n9258), .A4(n9257), 
        .ZN(n9261) );
  ND4D4BWP30P140LVT U9848 ( .A1(n9264), .A2(n9263), .A3(n9262), .A4(n9261), 
        .ZN(o_data_bus[252]) );
  AOI22D1BWP30P140LVT U9849 ( .A1(i_data_bus[90]), .A2(n9549), .B1(
        i_data_bus[730]), .B2(n9554), .ZN(n9285) );
  AOI22D1BWP30P140LVT U9850 ( .A1(i_data_bus[698]), .A2(n9559), .B1(
        i_data_bus[794]), .B2(n9547), .ZN(n9284) );
  AOI22D1BWP30P140LVT U9851 ( .A1(i_data_bus[1018]), .A2(n9571), .B1(
        i_data_bus[314]), .B2(n9584), .ZN(n9283) );
  AOI22D1BWP30P140LVT U9852 ( .A1(i_data_bus[58]), .A2(n9548), .B1(
        i_data_bus[826]), .B2(n9552), .ZN(n9268) );
  AOI22D1BWP30P140LVT U9853 ( .A1(i_data_bus[890]), .A2(n9556), .B1(
        i_data_bus[858]), .B2(n9557), .ZN(n9267) );
  AOI22D1BWP30P140LVT U9854 ( .A1(i_data_bus[122]), .A2(n9555), .B1(
        i_data_bus[666]), .B2(n9558), .ZN(n9266) );
  AOI22D1BWP30P140LVT U9855 ( .A1(i_data_bus[26]), .A2(n9553), .B1(
        i_data_bus[762]), .B2(n9546), .ZN(n9265) );
  ND4D1BWP30P140LVT U9856 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), 
        .ZN(n9281) );
  MOAI22D1BWP30P140LVT U9857 ( .A1(n9269), .A2(n9375), .B1(i_data_bus[250]), 
        .B2(n9568), .ZN(n9280) );
  AOI22D1BWP30P140LVT U9858 ( .A1(i_data_bus[954]), .A2(n9587), .B1(
        i_data_bus[282]), .B2(n9586), .ZN(n9273) );
  AOI22D1BWP30P140LVT U9859 ( .A1(i_data_bus[346]), .A2(n9570), .B1(
        i_data_bus[186]), .B2(n9583), .ZN(n9272) );
  AOI22D1BWP30P140LVT U9860 ( .A1(i_data_bus[538]), .A2(n9573), .B1(
        i_data_bus[570]), .B2(n9575), .ZN(n9271) );
  AOI22D1BWP30P140LVT U9861 ( .A1(i_data_bus[602]), .A2(n9572), .B1(
        i_data_bus[634]), .B2(n9574), .ZN(n9270) );
  ND4D1BWP30P140LVT U9862 ( .A1(n9273), .A2(n9272), .A3(n9271), .A4(n9270), 
        .ZN(n9279) );
  AOI22D1BWP30P140LVT U9863 ( .A1(i_data_bus[922]), .A2(n9581), .B1(
        i_data_bus[506]), .B2(n9580), .ZN(n9277) );
  AOI22D1BWP30P140LVT U9864 ( .A1(i_data_bus[154]), .A2(n9533), .B1(
        i_data_bus[474]), .B2(n9582), .ZN(n9276) );
  AOI22D1BWP30P140LVT U9865 ( .A1(i_data_bus[986]), .A2(n9551), .B1(
        i_data_bus[410]), .B2(n9585), .ZN(n9275) );
  AOI22D1BWP30P140LVT U9866 ( .A1(i_data_bus[442]), .A2(n9532), .B1(
        i_data_bus[218]), .B2(n9550), .ZN(n9274) );
  ND4D1BWP30P140LVT U9867 ( .A1(n9277), .A2(n9276), .A3(n9275), .A4(n9274), 
        .ZN(n9278) );
  NR4D0BWP30P140LVT U9868 ( .A1(n9281), .A2(n9280), .A3(n9279), .A4(n9278), 
        .ZN(n9282) );
  ND4D4BWP30P140LVT U9869 ( .A1(n9285), .A2(n9284), .A3(n9283), .A4(n9282), 
        .ZN(o_data_bus[250]) );
  AOI22D1BWP30P140LVT U9870 ( .A1(i_data_bus[695]), .A2(n9559), .B1(
        i_data_bus[791]), .B2(n9547), .ZN(n9307) );
  AOI22D1BWP30P140LVT U9871 ( .A1(i_data_bus[119]), .A2(n9555), .B1(
        i_data_bus[855]), .B2(n9557), .ZN(n9306) );
  AOI22D1BWP30P140LVT U9872 ( .A1(i_data_bus[1015]), .A2(n9571), .B1(
        i_data_bus[951]), .B2(n9587), .ZN(n9305) );
  AOI22D1BWP30P140LVT U9873 ( .A1(i_data_bus[23]), .A2(n9553), .B1(
        i_data_bus[727]), .B2(n9554), .ZN(n9289) );
  AOI22D1BWP30P140LVT U9874 ( .A1(i_data_bus[759]), .A2(n9546), .B1(
        i_data_bus[663]), .B2(n9558), .ZN(n9288) );
  AOI22D1BWP30P140LVT U9875 ( .A1(i_data_bus[87]), .A2(n9549), .B1(
        i_data_bus[887]), .B2(n9556), .ZN(n9287) );
  AOI22D1BWP30P140LVT U9876 ( .A1(i_data_bus[55]), .A2(n9548), .B1(
        i_data_bus[823]), .B2(n9552), .ZN(n9286) );
  ND4D1BWP30P140LVT U9877 ( .A1(n9289), .A2(n9288), .A3(n9287), .A4(n9286), 
        .ZN(n9303) );
  OAI22D1BWP30P140LVT U9878 ( .A1(n9291), .A2(n9566), .B1(n9290), .B2(n9375), 
        .ZN(n9302) );
  AOI22D1BWP30P140LVT U9879 ( .A1(i_data_bus[183]), .A2(n9583), .B1(
        i_data_bus[503]), .B2(n9580), .ZN(n9295) );
  AOI22D1BWP30P140LVT U9880 ( .A1(i_data_bus[215]), .A2(n9550), .B1(
        i_data_bus[343]), .B2(n9570), .ZN(n9294) );
  AOI22D1BWP30P140LVT U9881 ( .A1(i_data_bus[631]), .A2(n9574), .B1(
        i_data_bus[599]), .B2(n9572), .ZN(n9293) );
  AOI22D1BWP30P140LVT U9882 ( .A1(i_data_bus[535]), .A2(n9573), .B1(
        i_data_bus[567]), .B2(n9575), .ZN(n9292) );
  ND4D1BWP30P140LVT U9883 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), 
        .ZN(n9301) );
  AOI22D1BWP30P140LVT U9884 ( .A1(i_data_bus[279]), .A2(n9586), .B1(
        i_data_bus[407]), .B2(n9585), .ZN(n9299) );
  AOI22D1BWP30P140LVT U9885 ( .A1(i_data_bus[247]), .A2(n9568), .B1(
        i_data_bus[311]), .B2(n9584), .ZN(n9298) );
  AOI22D1BWP30P140LVT U9886 ( .A1(i_data_bus[471]), .A2(n9582), .B1(
        i_data_bus[151]), .B2(n9533), .ZN(n9297) );
  AOI22D1BWP30P140LVT U9887 ( .A1(i_data_bus[983]), .A2(n9551), .B1(
        i_data_bus[919]), .B2(n9581), .ZN(n9296) );
  ND4D1BWP30P140LVT U9888 ( .A1(n9299), .A2(n9298), .A3(n9297), .A4(n9296), 
        .ZN(n9300) );
  NR4D0BWP30P140LVT U9889 ( .A1(n9303), .A2(n9302), .A3(n9301), .A4(n9300), 
        .ZN(n9304) );
  ND4D4BWP30P140LVT U9890 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), 
        .ZN(o_data_bus[247]) );
  AOI22D1BWP30P140LVT U9891 ( .A1(i_data_bus[789]), .A2(n9547), .B1(
        i_data_bus[725]), .B2(n9554), .ZN(n9328) );
  AOI22D1BWP30P140LVT U9892 ( .A1(i_data_bus[53]), .A2(n9548), .B1(
        i_data_bus[821]), .B2(n9552), .ZN(n9327) );
  AOI22D1BWP30P140LVT U9893 ( .A1(i_data_bus[213]), .A2(n9550), .B1(
        i_data_bus[277]), .B2(n9586), .ZN(n9326) );
  AOI22D1BWP30P140LVT U9894 ( .A1(i_data_bus[21]), .A2(n9553), .B1(
        i_data_bus[853]), .B2(n9557), .ZN(n9311) );
  AOI22D1BWP30P140LVT U9895 ( .A1(i_data_bus[661]), .A2(n9558), .B1(
        i_data_bus[693]), .B2(n9559), .ZN(n9310) );
  AOI22D1BWP30P140LVT U9896 ( .A1(i_data_bus[117]), .A2(n9555), .B1(
        i_data_bus[757]), .B2(n9546), .ZN(n9309) );
  AOI22D1BWP30P140LVT U9897 ( .A1(i_data_bus[85]), .A2(n9549), .B1(
        i_data_bus[885]), .B2(n9556), .ZN(n9308) );
  ND4D1BWP30P140LVT U9898 ( .A1(n9311), .A2(n9310), .A3(n9309), .A4(n9308), 
        .ZN(n9324) );
  MOAI22D1BWP30P140LVT U9899 ( .A1(n9312), .A2(n9375), .B1(i_data_bus[181]), 
        .B2(n9583), .ZN(n9323) );
  AOI22D1BWP30P140LVT U9900 ( .A1(i_data_bus[981]), .A2(n9551), .B1(
        i_data_bus[341]), .B2(n9570), .ZN(n9316) );
  AOI22D1BWP30P140LVT U9901 ( .A1(i_data_bus[917]), .A2(n9581), .B1(
        i_data_bus[1013]), .B2(n9571), .ZN(n9315) );
  AOI22D1BWP30P140LVT U9902 ( .A1(i_data_bus[597]), .A2(n9572), .B1(
        i_data_bus[565]), .B2(n9575), .ZN(n9314) );
  AOI22D1BWP30P140LVT U9903 ( .A1(i_data_bus[629]), .A2(n9574), .B1(
        i_data_bus[533]), .B2(n9573), .ZN(n9313) );
  ND4D1BWP30P140LVT U9904 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), 
        .ZN(n9322) );
  AOI22D1BWP30P140LVT U9905 ( .A1(i_data_bus[501]), .A2(n9580), .B1(
        i_data_bus[469]), .B2(n9582), .ZN(n9320) );
  AOI22D1BWP30P140LVT U9906 ( .A1(i_data_bus[949]), .A2(n9587), .B1(
        i_data_bus[149]), .B2(n9533), .ZN(n9319) );
  AOI22D1BWP30P140LVT U9907 ( .A1(i_data_bus[437]), .A2(n9532), .B1(
        i_data_bus[245]), .B2(n9568), .ZN(n9318) );
  AOI22D1BWP30P140LVT U9908 ( .A1(i_data_bus[309]), .A2(n9584), .B1(
        i_data_bus[405]), .B2(n9585), .ZN(n9317) );
  ND4D1BWP30P140LVT U9909 ( .A1(n9320), .A2(n9319), .A3(n9318), .A4(n9317), 
        .ZN(n9321) );
  NR4D0BWP30P140LVT U9910 ( .A1(n9324), .A2(n9323), .A3(n9322), .A4(n9321), 
        .ZN(n9325) );
  ND4D4BWP30P140LVT U9911 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), 
        .ZN(o_data_bus[245]) );
  AOI22D1BWP30P140LVT U9912 ( .A1(i_data_bus[37]), .A2(n9548), .B1(
        i_data_bus[645]), .B2(n9558), .ZN(n9349) );
  AOI22D1BWP30P140LVT U9913 ( .A1(i_data_bus[69]), .A2(n9549), .B1(
        i_data_bus[805]), .B2(n9552), .ZN(n9348) );
  AOI22D1BWP30P140LVT U9914 ( .A1(i_data_bus[165]), .A2(n9583), .B1(
        i_data_bus[389]), .B2(n9585), .ZN(n9347) );
  AOI22D1BWP30P140LVT U9915 ( .A1(i_data_bus[101]), .A2(n9555), .B1(
        i_data_bus[677]), .B2(n9559), .ZN(n9332) );
  AOI22D1BWP30P140LVT U9916 ( .A1(i_data_bus[837]), .A2(n9557), .B1(
        i_data_bus[869]), .B2(n9556), .ZN(n9331) );
  AOI22D1BWP30P140LVT U9917 ( .A1(i_data_bus[5]), .A2(n9553), .B1(
        i_data_bus[773]), .B2(n9547), .ZN(n9330) );
  AOI22D1BWP30P140LVT U9918 ( .A1(i_data_bus[709]), .A2(n9554), .B1(
        i_data_bus[741]), .B2(n9546), .ZN(n9329) );
  ND4D1BWP30P140LVT U9919 ( .A1(n9332), .A2(n9331), .A3(n9330), .A4(n9329), 
        .ZN(n9345) );
  MOAI22D1BWP30P140LVT U9920 ( .A1(n9333), .A2(n9461), .B1(i_data_bus[453]), 
        .B2(n9582), .ZN(n9344) );
  AOI22D1BWP30P140LVT U9921 ( .A1(i_data_bus[933]), .A2(n9587), .B1(
        i_data_bus[261]), .B2(n9586), .ZN(n9337) );
  AOI22D1BWP30P140LVT U9922 ( .A1(i_data_bus[901]), .A2(n9581), .B1(
        i_data_bus[197]), .B2(n9550), .ZN(n9336) );
  AOI22D1BWP30P140LVT U9923 ( .A1(i_data_bus[581]), .A2(n9572), .B1(
        i_data_bus[613]), .B2(n9574), .ZN(n9335) );
  AOI22D1BWP30P140LVT U9924 ( .A1(i_data_bus[517]), .A2(n9573), .B1(
        i_data_bus[549]), .B2(n9575), .ZN(n9334) );
  ND4D1BWP30P140LVT U9925 ( .A1(n9337), .A2(n9336), .A3(n9335), .A4(n9334), 
        .ZN(n9343) );
  AOI22D1BWP30P140LVT U9926 ( .A1(i_data_bus[965]), .A2(n9551), .B1(
        i_data_bus[485]), .B2(n9580), .ZN(n9341) );
  AOI22D1BWP30P140LVT U9927 ( .A1(i_data_bus[997]), .A2(n9571), .B1(
        i_data_bus[325]), .B2(n9570), .ZN(n9340) );
  AOI22D1BWP30P140LVT U9928 ( .A1(i_data_bus[133]), .A2(n9533), .B1(
        i_data_bus[229]), .B2(n9568), .ZN(n9339) );
  AOI22D1BWP30P140LVT U9929 ( .A1(i_data_bus[357]), .A2(n9569), .B1(
        i_data_bus[421]), .B2(n9532), .ZN(n9338) );
  ND4D1BWP30P140LVT U9930 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), 
        .ZN(n9342) );
  NR4D0BWP30P140LVT U9931 ( .A1(n9345), .A2(n9344), .A3(n9343), .A4(n9342), 
        .ZN(n9346) );
  ND4D4BWP30P140LVT U9932 ( .A1(n9349), .A2(n9348), .A3(n9347), .A4(n9346), 
        .ZN(o_data_bus[229]) );
  AOI22D1BWP30P140LVT U9933 ( .A1(i_data_bus[788]), .A2(n9547), .B1(
        i_data_bus[692]), .B2(n9559), .ZN(n9370) );
  AOI22D1BWP30P140LVT U9934 ( .A1(i_data_bus[52]), .A2(n9548), .B1(
        i_data_bus[84]), .B2(n9549), .ZN(n9369) );
  AOI22D1BWP30P140LVT U9935 ( .A1(i_data_bus[244]), .A2(n9568), .B1(
        i_data_bus[436]), .B2(n9532), .ZN(n9368) );
  AOI22D1BWP30P140LVT U9936 ( .A1(i_data_bus[20]), .A2(n9553), .B1(
        i_data_bus[724]), .B2(n9554), .ZN(n9353) );
  AOI22D1BWP30P140LVT U9937 ( .A1(i_data_bus[820]), .A2(n9552), .B1(
        i_data_bus[660]), .B2(n9558), .ZN(n9352) );
  AOI22D1BWP30P140LVT U9938 ( .A1(i_data_bus[116]), .A2(n9555), .B1(
        i_data_bus[756]), .B2(n9546), .ZN(n9351) );
  AOI22D1BWP30P140LVT U9939 ( .A1(i_data_bus[852]), .A2(n9557), .B1(
        i_data_bus[884]), .B2(n9556), .ZN(n9350) );
  ND4D1BWP30P140LVT U9940 ( .A1(n9353), .A2(n9352), .A3(n9351), .A4(n9350), 
        .ZN(n9366) );
  MOAI22D1BWP30P140LVT U9941 ( .A1(n9354), .A2(n9461), .B1(i_data_bus[276]), 
        .B2(n9586), .ZN(n9365) );
  AOI22D1BWP30P140LVT U9942 ( .A1(i_data_bus[948]), .A2(n9587), .B1(
        i_data_bus[148]), .B2(n9533), .ZN(n9358) );
  AOI22D1BWP30P140LVT U9943 ( .A1(i_data_bus[980]), .A2(n9551), .B1(
        i_data_bus[404]), .B2(n9585), .ZN(n9357) );
  AOI22D1BWP30P140LVT U9944 ( .A1(i_data_bus[596]), .A2(n9572), .B1(
        i_data_bus[564]), .B2(n9575), .ZN(n9356) );
  AOI22D1BWP30P140LVT U9945 ( .A1(i_data_bus[532]), .A2(n9573), .B1(
        i_data_bus[628]), .B2(n9574), .ZN(n9355) );
  ND4D1BWP30P140LVT U9946 ( .A1(n9358), .A2(n9357), .A3(n9356), .A4(n9355), 
        .ZN(n9364) );
  AOI22D1BWP30P140LVT U9947 ( .A1(i_data_bus[340]), .A2(n9570), .B1(
        i_data_bus[500]), .B2(n9580), .ZN(n9362) );
  AOI22D1BWP30P140LVT U9948 ( .A1(i_data_bus[1012]), .A2(n9571), .B1(
        i_data_bus[180]), .B2(n9583), .ZN(n9361) );
  AOI22D1BWP30P140LVT U9949 ( .A1(i_data_bus[916]), .A2(n9581), .B1(
        i_data_bus[468]), .B2(n9582), .ZN(n9360) );
  AOI22D1BWP30P140LVT U9950 ( .A1(i_data_bus[212]), .A2(n9550), .B1(
        i_data_bus[372]), .B2(n9569), .ZN(n9359) );
  ND4D1BWP30P140LVT U9951 ( .A1(n9362), .A2(n9361), .A3(n9360), .A4(n9359), 
        .ZN(n9363) );
  NR4D0BWP30P140LVT U9952 ( .A1(n9366), .A2(n9365), .A3(n9364), .A4(n9363), 
        .ZN(n9367) );
  ND4D4BWP30P140LVT U9953 ( .A1(n9370), .A2(n9369), .A3(n9368), .A4(n9367), 
        .ZN(o_data_bus[244]) );
  AOI22D1BWP30P140LVT U9954 ( .A1(i_data_bus[657]), .A2(n9558), .B1(
        i_data_bus[753]), .B2(n9546), .ZN(n9392) );
  AOI22D1BWP30P140LVT U9955 ( .A1(i_data_bus[49]), .A2(n9548), .B1(
        i_data_bus[689]), .B2(n9559), .ZN(n9391) );
  AOI22D1BWP30P140LVT U9956 ( .A1(i_data_bus[1009]), .A2(n9571), .B1(
        i_data_bus[401]), .B2(n9585), .ZN(n9390) );
  AOI22D1BWP30P140LVT U9957 ( .A1(i_data_bus[17]), .A2(n9553), .B1(
        i_data_bus[849]), .B2(n9557), .ZN(n9374) );
  AOI22D1BWP30P140LVT U9958 ( .A1(i_data_bus[785]), .A2(n9547), .B1(
        i_data_bus[721]), .B2(n9554), .ZN(n9373) );
  AOI22D1BWP30P140LVT U9959 ( .A1(i_data_bus[881]), .A2(n9556), .B1(
        i_data_bus[817]), .B2(n9552), .ZN(n9372) );
  AOI22D1BWP30P140LVT U9960 ( .A1(i_data_bus[81]), .A2(n9549), .B1(
        i_data_bus[113]), .B2(n9555), .ZN(n9371) );
  ND4D1BWP30P140LVT U9961 ( .A1(n9374), .A2(n9373), .A3(n9372), .A4(n9371), 
        .ZN(n9388) );
  MOAI22D1BWP30P140LVT U9962 ( .A1(n9376), .A2(n9375), .B1(i_data_bus[497]), 
        .B2(n9580), .ZN(n9387) );
  AOI22D1BWP30P140LVT U9963 ( .A1(i_data_bus[241]), .A2(n9568), .B1(
        i_data_bus[273]), .B2(n9586), .ZN(n9380) );
  AOI22D1BWP30P140LVT U9964 ( .A1(i_data_bus[977]), .A2(n9551), .B1(
        i_data_bus[433]), .B2(n9532), .ZN(n9379) );
  AOI22D1BWP30P140LVT U9965 ( .A1(i_data_bus[593]), .A2(n9572), .B1(
        i_data_bus[561]), .B2(n9575), .ZN(n9378) );
  AOI22D1BWP30P140LVT U9966 ( .A1(i_data_bus[625]), .A2(n9574), .B1(
        i_data_bus[529]), .B2(n9573), .ZN(n9377) );
  ND4D1BWP30P140LVT U9967 ( .A1(n9380), .A2(n9379), .A3(n9378), .A4(n9377), 
        .ZN(n9386) );
  AOI22D1BWP30P140LVT U9968 ( .A1(i_data_bus[337]), .A2(n9570), .B1(
        i_data_bus[145]), .B2(n9533), .ZN(n9384) );
  AOI22D1BWP30P140LVT U9969 ( .A1(i_data_bus[209]), .A2(n9550), .B1(
        i_data_bus[305]), .B2(n9584), .ZN(n9383) );
  AOI22D1BWP30P140LVT U9970 ( .A1(i_data_bus[945]), .A2(n9587), .B1(
        i_data_bus[465]), .B2(n9582), .ZN(n9382) );
  AOI22D1BWP30P140LVT U9971 ( .A1(i_data_bus[913]), .A2(n9581), .B1(
        i_data_bus[177]), .B2(n9583), .ZN(n9381) );
  ND4D1BWP30P140LVT U9972 ( .A1(n9384), .A2(n9383), .A3(n9382), .A4(n9381), 
        .ZN(n9385) );
  NR4D0BWP30P140LVT U9973 ( .A1(n9388), .A2(n9387), .A3(n9386), .A4(n9385), 
        .ZN(n9389) );
  ND4D4BWP30P140LVT U9974 ( .A1(n9392), .A2(n9391), .A3(n9390), .A4(n9389), 
        .ZN(o_data_bus[241]) );
  AOI22D1BWP30P140LVT U9975 ( .A1(i_data_bus[46]), .A2(n9548), .B1(
        i_data_bus[654]), .B2(n9558), .ZN(n9414) );
  AOI22D1BWP30P140LVT U9976 ( .A1(i_data_bus[110]), .A2(n9555), .B1(
        i_data_bus[78]), .B2(n9549), .ZN(n9413) );
  AOI22D1BWP30P140LVT U9977 ( .A1(i_data_bus[942]), .A2(n9587), .B1(
        i_data_bus[174]), .B2(n9583), .ZN(n9412) );
  AOI22D1BWP30P140LVT U9978 ( .A1(i_data_bus[814]), .A2(n9552), .B1(
        i_data_bus[846]), .B2(n9557), .ZN(n9396) );
  AOI22D1BWP30P140LVT U9979 ( .A1(i_data_bus[14]), .A2(n9553), .B1(
        i_data_bus[878]), .B2(n9556), .ZN(n9395) );
  AOI22D1BWP30P140LVT U9980 ( .A1(i_data_bus[782]), .A2(n9547), .B1(
        i_data_bus[686]), .B2(n9559), .ZN(n9394) );
  AOI22D1BWP30P140LVT U9981 ( .A1(i_data_bus[750]), .A2(n9546), .B1(
        i_data_bus[718]), .B2(n9554), .ZN(n9393) );
  ND4D1BWP30P140LVT U9982 ( .A1(n9396), .A2(n9395), .A3(n9394), .A4(n9393), 
        .ZN(n9410) );
  MOAI22D1BWP30P140LVT U9983 ( .A1(n9398), .A2(n9397), .B1(i_data_bus[302]), 
        .B2(n9584), .ZN(n9409) );
  AOI22D1BWP30P140LVT U9984 ( .A1(i_data_bus[270]), .A2(n9586), .B1(
        i_data_bus[206]), .B2(n9550), .ZN(n9402) );
  AOI22D1BWP30P140LVT U9985 ( .A1(i_data_bus[910]), .A2(n9581), .B1(
        i_data_bus[334]), .B2(n9570), .ZN(n9401) );
  AOI22D1BWP30P140LVT U9986 ( .A1(i_data_bus[558]), .A2(n9575), .B1(
        i_data_bus[526]), .B2(n9573), .ZN(n9400) );
  AOI22D1BWP30P140LVT U9987 ( .A1(i_data_bus[590]), .A2(n9572), .B1(
        i_data_bus[622]), .B2(n9574), .ZN(n9399) );
  ND4D1BWP30P140LVT U9988 ( .A1(n9402), .A2(n9401), .A3(n9400), .A4(n9399), 
        .ZN(n9408) );
  AOI22D1BWP30P140LVT U9989 ( .A1(i_data_bus[366]), .A2(n9569), .B1(
        i_data_bus[462]), .B2(n9582), .ZN(n9406) );
  AOI22D1BWP30P140LVT U9990 ( .A1(i_data_bus[142]), .A2(n9533), .B1(
        i_data_bus[398]), .B2(n9585), .ZN(n9405) );
  AOI22D1BWP30P140LVT U9991 ( .A1(i_data_bus[1006]), .A2(n9571), .B1(
        i_data_bus[430]), .B2(n9532), .ZN(n9404) );
  AOI22D1BWP30P140LVT U9992 ( .A1(i_data_bus[974]), .A2(n9551), .B1(
        i_data_bus[238]), .B2(n9568), .ZN(n9403) );
  ND4D1BWP30P140LVT U9993 ( .A1(n9406), .A2(n9405), .A3(n9404), .A4(n9403), 
        .ZN(n9407) );
  NR4D0BWP30P140LVT U9994 ( .A1(n9410), .A2(n9409), .A3(n9408), .A4(n9407), 
        .ZN(n9411) );
  ND4D4BWP30P140LVT U9995 ( .A1(n9414), .A2(n9413), .A3(n9412), .A4(n9411), 
        .ZN(o_data_bus[238]) );
  AOI22D1BWP30P140LVT U9996 ( .A1(i_data_bus[45]), .A2(n9548), .B1(
        i_data_bus[717]), .B2(n9554), .ZN(n9436) );
  AOI22D1BWP30P140LVT U9997 ( .A1(i_data_bus[845]), .A2(n9557), .B1(
        i_data_bus[813]), .B2(n9552), .ZN(n9435) );
  AOI22D1BWP30P140LVT U9998 ( .A1(i_data_bus[237]), .A2(n9568), .B1(
        i_data_bus[141]), .B2(n9533), .ZN(n9434) );
  AOI22D1BWP30P140LVT U9999 ( .A1(i_data_bus[781]), .A2(n9547), .B1(
        i_data_bus[749]), .B2(n9546), .ZN(n9418) );
  AOI22D1BWP30P140LVT U10000 ( .A1(i_data_bus[77]), .A2(n9549), .B1(
        i_data_bus[685]), .B2(n9559), .ZN(n9417) );
  AOI22D1BWP30P140LVT U10001 ( .A1(i_data_bus[109]), .A2(n9555), .B1(
        i_data_bus[877]), .B2(n9556), .ZN(n9416) );
  AOI22D1BWP30P140LVT U10002 ( .A1(i_data_bus[13]), .A2(n9553), .B1(
        i_data_bus[653]), .B2(n9558), .ZN(n9415) );
  ND4D1BWP30P140LVT U10003 ( .A1(n9418), .A2(n9417), .A3(n9416), .A4(n9415), 
        .ZN(n9432) );
  MOAI22D1BWP30P140LVT U10004 ( .A1(n9420), .A2(n9419), .B1(i_data_bus[365]), 
        .B2(n9569), .ZN(n9431) );
  AOI22D1BWP30P140LVT U10005 ( .A1(i_data_bus[909]), .A2(n9581), .B1(
        i_data_bus[461]), .B2(n9582), .ZN(n9424) );
  AOI22D1BWP30P140LVT U10006 ( .A1(i_data_bus[973]), .A2(n9551), .B1(
        i_data_bus[1005]), .B2(n9571), .ZN(n9423) );
  AOI22D1BWP30P140LVT U10007 ( .A1(i_data_bus[621]), .A2(n9574), .B1(
        i_data_bus[557]), .B2(n9575), .ZN(n9422) );
  AOI22D1BWP30P140LVT U10008 ( .A1(i_data_bus[525]), .A2(n9573), .B1(
        i_data_bus[589]), .B2(n9572), .ZN(n9421) );
  ND4D1BWP30P140LVT U10009 ( .A1(n9424), .A2(n9423), .A3(n9422), .A4(n9421), 
        .ZN(n9430) );
  AOI22D1BWP30P140LVT U10010 ( .A1(i_data_bus[269]), .A2(n9586), .B1(
        i_data_bus[429]), .B2(n9532), .ZN(n9428) );
  AOI22D1BWP30P140LVT U10011 ( .A1(i_data_bus[397]), .A2(n9585), .B1(
        i_data_bus[493]), .B2(n9580), .ZN(n9427) );
  AOI22D1BWP30P140LVT U10012 ( .A1(i_data_bus[941]), .A2(n9587), .B1(
        i_data_bus[333]), .B2(n9570), .ZN(n9426) );
  AOI22D1BWP30P140LVT U10013 ( .A1(i_data_bus[205]), .A2(n9550), .B1(
        i_data_bus[301]), .B2(n9584), .ZN(n9425) );
  ND4D1BWP30P140LVT U10014 ( .A1(n9428), .A2(n9427), .A3(n9426), .A4(n9425), 
        .ZN(n9429) );
  NR4D0BWP30P140LVT U10015 ( .A1(n9432), .A2(n9431), .A3(n9430), .A4(n9429), 
        .ZN(n9433) );
  ND4D4BWP30P140LVT U10016 ( .A1(n9436), .A2(n9435), .A3(n9434), .A4(n9433), 
        .ZN(o_data_bus[237]) );
  AOI22D1BWP30P140LVT U10017 ( .A1(i_data_bus[73]), .A2(n9549), .B1(
        i_data_bus[105]), .B2(n9555), .ZN(n9456) );
  AOI22D1BWP30P140LVT U10018 ( .A1(i_data_bus[777]), .A2(n9547), .B1(
        i_data_bus[649]), .B2(n9558), .ZN(n9455) );
  AOI22D1BWP30P140LVT U10019 ( .A1(i_data_bus[969]), .A2(n9551), .B1(
        i_data_bus[329]), .B2(n9570), .ZN(n9454) );
  AOI22D1BWP30P140LVT U10020 ( .A1(i_data_bus[873]), .A2(n9556), .B1(
        i_data_bus[841]), .B2(n9557), .ZN(n9440) );
  AOI22D1BWP30P140LVT U10021 ( .A1(i_data_bus[41]), .A2(n9548), .B1(
        i_data_bus[713]), .B2(n9554), .ZN(n9439) );
  AOI22D1BWP30P140LVT U10022 ( .A1(i_data_bus[9]), .A2(n9553), .B1(
        i_data_bus[809]), .B2(n9552), .ZN(n9438) );
  AOI22D1BWP30P140LVT U10023 ( .A1(i_data_bus[745]), .A2(n9546), .B1(
        i_data_bus[681]), .B2(n9559), .ZN(n9437) );
  ND4D1BWP30P140LVT U10024 ( .A1(n9440), .A2(n9439), .A3(n9438), .A4(n9437), 
        .ZN(n9452) );
  MOAI22D1BWP30P140LVT U10025 ( .A1(n9688), .A2(n9461), .B1(i_data_bus[137]), 
        .B2(n9533), .ZN(n9451) );
  AOI22D1BWP30P140LVT U10026 ( .A1(i_data_bus[905]), .A2(n9581), .B1(
        i_data_bus[937]), .B2(n9587), .ZN(n9444) );
  AOI22D1BWP30P140LVT U10027 ( .A1(i_data_bus[1001]), .A2(n9571), .B1(
        i_data_bus[489]), .B2(n9580), .ZN(n9443) );
  AOI22D1BWP30P140LVT U10028 ( .A1(i_data_bus[617]), .A2(n9574), .B1(
        i_data_bus[553]), .B2(n9575), .ZN(n9442) );
  AOI22D1BWP30P140LVT U10029 ( .A1(i_data_bus[521]), .A2(n9573), .B1(
        i_data_bus[585]), .B2(n9572), .ZN(n9441) );
  ND4D1BWP30P140LVT U10030 ( .A1(n9444), .A2(n9443), .A3(n9442), .A4(n9441), 
        .ZN(n9450) );
  AOI22D1BWP30P140LVT U10031 ( .A1(i_data_bus[233]), .A2(n9568), .B1(
        i_data_bus[265]), .B2(n9586), .ZN(n9448) );
  AOI22D1BWP30P140LVT U10032 ( .A1(i_data_bus[425]), .A2(n9532), .B1(
        i_data_bus[457]), .B2(n9582), .ZN(n9447) );
  AOI22D1BWP30P140LVT U10033 ( .A1(i_data_bus[201]), .A2(n9550), .B1(
        i_data_bus[169]), .B2(n9583), .ZN(n9446) );
  AOI22D1BWP30P140LVT U10034 ( .A1(i_data_bus[361]), .A2(n9569), .B1(
        i_data_bus[393]), .B2(n9585), .ZN(n9445) );
  ND4D1BWP30P140LVT U10035 ( .A1(n9448), .A2(n9447), .A3(n9446), .A4(n9445), 
        .ZN(n9449) );
  NR4D0BWP30P140LVT U10036 ( .A1(n9452), .A2(n9451), .A3(n9450), .A4(n9449), 
        .ZN(n9453) );
  ND4D4BWP30P140LVT U10037 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), 
        .ZN(o_data_bus[233]) );
  AOI22D1BWP30P140LVT U10038 ( .A1(i_data_bus[744]), .A2(n9546), .B1(
        i_data_bus[680]), .B2(n9559), .ZN(n9478) );
  AOI22D1BWP30P140LVT U10039 ( .A1(i_data_bus[104]), .A2(n9555), .B1(
        i_data_bus[72]), .B2(n9549), .ZN(n9477) );
  AOI22D1BWP30P140LVT U10040 ( .A1(i_data_bus[200]), .A2(n9550), .B1(
        i_data_bus[136]), .B2(n9533), .ZN(n9476) );
  AOI22D1BWP30P140LVT U10041 ( .A1(i_data_bus[808]), .A2(n9552), .B1(
        i_data_bus[776]), .B2(n9547), .ZN(n9460) );
  AOI22D1BWP30P140LVT U10042 ( .A1(i_data_bus[8]), .A2(n9553), .B1(
        i_data_bus[40]), .B2(n9548), .ZN(n9459) );
  AOI22D1BWP30P140LVT U10043 ( .A1(i_data_bus[872]), .A2(n9556), .B1(
        i_data_bus[648]), .B2(n9558), .ZN(n9458) );
  AOI22D1BWP30P140LVT U10044 ( .A1(i_data_bus[840]), .A2(n9557), .B1(
        i_data_bus[712]), .B2(n9554), .ZN(n9457) );
  ND4D1BWP30P140LVT U10045 ( .A1(n9460), .A2(n9459), .A3(n9458), .A4(n9457), 
        .ZN(n9474) );
  MOAI22D1BWP30P140LVT U10046 ( .A1(n9462), .A2(n9461), .B1(i_data_bus[424]), 
        .B2(n9532), .ZN(n9473) );
  AOI22D1BWP30P140LVT U10047 ( .A1(i_data_bus[168]), .A2(n9583), .B1(
        i_data_bus[392]), .B2(n9585), .ZN(n9466) );
  AOI22D1BWP30P140LVT U10048 ( .A1(i_data_bus[936]), .A2(n9587), .B1(
        i_data_bus[456]), .B2(n9582), .ZN(n9465) );
  AOI22D1BWP30P140LVT U10049 ( .A1(i_data_bus[584]), .A2(n9572), .B1(
        i_data_bus[520]), .B2(n9573), .ZN(n9464) );
  AOI22D1BWP30P140LVT U10050 ( .A1(i_data_bus[616]), .A2(n9574), .B1(
        i_data_bus[552]), .B2(n9575), .ZN(n9463) );
  ND4D1BWP30P140LVT U10051 ( .A1(n9466), .A2(n9465), .A3(n9464), .A4(n9463), 
        .ZN(n9472) );
  AOI22D1BWP30P140LVT U10052 ( .A1(i_data_bus[968]), .A2(n9551), .B1(
        i_data_bus[488]), .B2(n9580), .ZN(n9470) );
  AOI22D1BWP30P140LVT U10053 ( .A1(i_data_bus[1000]), .A2(n9571), .B1(
        i_data_bus[904]), .B2(n9581), .ZN(n9469) );
  AOI22D1BWP30P140LVT U10054 ( .A1(i_data_bus[264]), .A2(n9586), .B1(
        i_data_bus[360]), .B2(n9569), .ZN(n9468) );
  AOI22D1BWP30P140LVT U10055 ( .A1(i_data_bus[328]), .A2(n9570), .B1(
        i_data_bus[232]), .B2(n9568), .ZN(n9467) );
  ND4D1BWP30P140LVT U10056 ( .A1(n9470), .A2(n9469), .A3(n9468), .A4(n9467), 
        .ZN(n9471) );
  NR4D0BWP30P140LVT U10057 ( .A1(n9474), .A2(n9473), .A3(n9472), .A4(n9471), 
        .ZN(n9475) );
  ND4D4BWP30P140LVT U10058 ( .A1(n9478), .A2(n9477), .A3(n9476), .A4(n9475), 
        .ZN(o_data_bus[232]) );
  AOI22D1BWP30P140LVT U10059 ( .A1(i_data_bus[839]), .A2(n9557), .B1(
        i_data_bus[647]), .B2(n9558), .ZN(n9500) );
  AOI22D1BWP30P140LVT U10060 ( .A1(i_data_bus[103]), .A2(n9555), .B1(
        i_data_bus[743]), .B2(n9546), .ZN(n9499) );
  AOI22D1BWP30P140LVT U10061 ( .A1(i_data_bus[967]), .A2(n9551), .B1(
        i_data_bus[295]), .B2(n9584), .ZN(n9498) );
  AOI22D1BWP30P140LVT U10062 ( .A1(i_data_bus[39]), .A2(n9548), .B1(
        i_data_bus[7]), .B2(n9553), .ZN(n9482) );
  AOI22D1BWP30P140LVT U10063 ( .A1(i_data_bus[807]), .A2(n9552), .B1(
        i_data_bus[711]), .B2(n9554), .ZN(n9481) );
  AOI22D1BWP30P140LVT U10064 ( .A1(i_data_bus[71]), .A2(n9549), .B1(
        i_data_bus[871]), .B2(n9556), .ZN(n9480) );
  AOI22D1BWP30P140LVT U10065 ( .A1(i_data_bus[679]), .A2(n9559), .B1(
        i_data_bus[775]), .B2(n9547), .ZN(n9479) );
  ND4D1BWP30P140LVT U10066 ( .A1(n9482), .A2(n9481), .A3(n9480), .A4(n9479), 
        .ZN(n9496) );
  MOAI22D1BWP30P140LVT U10067 ( .A1(n9484), .A2(n9483), .B1(i_data_bus[391]), 
        .B2(n9585), .ZN(n9495) );
  AOI22D1BWP30P140LVT U10068 ( .A1(i_data_bus[935]), .A2(n9587), .B1(
        i_data_bus[487]), .B2(n9580), .ZN(n9488) );
  AOI22D1BWP30P140LVT U10069 ( .A1(i_data_bus[455]), .A2(n9582), .B1(
        i_data_bus[327]), .B2(n9570), .ZN(n9487) );
  AOI22D1BWP30P140LVT U10070 ( .A1(i_data_bus[519]), .A2(n9573), .B1(
        i_data_bus[583]), .B2(n9572), .ZN(n9486) );
  AOI22D1BWP30P140LVT U10071 ( .A1(i_data_bus[615]), .A2(n9574), .B1(
        i_data_bus[551]), .B2(n9575), .ZN(n9485) );
  ND4D1BWP30P140LVT U10072 ( .A1(n9488), .A2(n9487), .A3(n9486), .A4(n9485), 
        .ZN(n9494) );
  AOI22D1BWP30P140LVT U10073 ( .A1(i_data_bus[263]), .A2(n9586), .B1(
        i_data_bus[135]), .B2(n9533), .ZN(n9492) );
  AOI22D1BWP30P140LVT U10074 ( .A1(i_data_bus[359]), .A2(n9569), .B1(
        i_data_bus[231]), .B2(n9568), .ZN(n9491) );
  AOI22D1BWP30P140LVT U10075 ( .A1(i_data_bus[903]), .A2(n9581), .B1(
        i_data_bus[999]), .B2(n9571), .ZN(n9490) );
  AOI22D1BWP30P140LVT U10076 ( .A1(i_data_bus[167]), .A2(n9583), .B1(
        i_data_bus[423]), .B2(n9532), .ZN(n9489) );
  ND4D1BWP30P140LVT U10077 ( .A1(n9492), .A2(n9491), .A3(n9490), .A4(n9489), 
        .ZN(n9493) );
  NR4D0BWP30P140LVT U10078 ( .A1(n9496), .A2(n9495), .A3(n9494), .A4(n9493), 
        .ZN(n9497) );
  ND4D4BWP30P140LVT U10079 ( .A1(n9500), .A2(n9499), .A3(n9498), .A4(n9497), 
        .ZN(o_data_bus[231]) );
  AOI22D1BWP30P140LVT U10080 ( .A1(i_data_bus[742]), .A2(n9546), .B1(
        i_data_bus[710]), .B2(n9554), .ZN(n9521) );
  AOI22D1BWP30P140LVT U10081 ( .A1(i_data_bus[6]), .A2(n9553), .B1(
        i_data_bus[678]), .B2(n9559), .ZN(n9520) );
  AOI22D1BWP30P140LVT U10082 ( .A1(i_data_bus[934]), .A2(n9587), .B1(
        i_data_bus[390]), .B2(n9585), .ZN(n9519) );
  AOI22D1BWP30P140LVT U10083 ( .A1(i_data_bus[70]), .A2(n9549), .B1(
        i_data_bus[870]), .B2(n9556), .ZN(n9504) );
  AOI22D1BWP30P140LVT U10084 ( .A1(i_data_bus[38]), .A2(n9548), .B1(
        i_data_bus[838]), .B2(n9557), .ZN(n9503) );
  AOI22D1BWP30P140LVT U10085 ( .A1(i_data_bus[806]), .A2(n9552), .B1(
        i_data_bus[646]), .B2(n9558), .ZN(n9502) );
  AOI22D1BWP30P140LVT U10086 ( .A1(i_data_bus[102]), .A2(n9555), .B1(
        i_data_bus[774]), .B2(n9547), .ZN(n9501) );
  ND4D1BWP30P140LVT U10087 ( .A1(n9504), .A2(n9503), .A3(n9502), .A4(n9501), 
        .ZN(n9517) );
  MOAI22D1BWP30P140LVT U10088 ( .A1(n9505), .A2(n9526), .B1(i_data_bus[262]), 
        .B2(n9586), .ZN(n9516) );
  AOI22D1BWP30P140LVT U10089 ( .A1(i_data_bus[230]), .A2(n9568), .B1(
        i_data_bus[358]), .B2(n9569), .ZN(n9509) );
  AOI22D1BWP30P140LVT U10090 ( .A1(i_data_bus[486]), .A2(n9580), .B1(
        i_data_bus[134]), .B2(n9533), .ZN(n9508) );
  AOI22D1BWP30P140LVT U10091 ( .A1(i_data_bus[582]), .A2(n9572), .B1(
        i_data_bus[550]), .B2(n9575), .ZN(n9507) );
  AOI22D1BWP30P140LVT U10092 ( .A1(i_data_bus[614]), .A2(n9574), .B1(
        i_data_bus[518]), .B2(n9573), .ZN(n9506) );
  ND4D1BWP30P140LVT U10093 ( .A1(n9509), .A2(n9508), .A3(n9507), .A4(n9506), 
        .ZN(n9515) );
  AOI22D1BWP30P140LVT U10094 ( .A1(i_data_bus[902]), .A2(n9581), .B1(
        i_data_bus[326]), .B2(n9570), .ZN(n9513) );
  AOI22D1BWP30P140LVT U10095 ( .A1(i_data_bus[998]), .A2(n9571), .B1(
        i_data_bus[198]), .B2(n9550), .ZN(n9512) );
  AOI22D1BWP30P140LVT U10096 ( .A1(i_data_bus[166]), .A2(n9583), .B1(
        i_data_bus[422]), .B2(n9532), .ZN(n9511) );
  AOI22D1BWP30P140LVT U10097 ( .A1(i_data_bus[966]), .A2(n9551), .B1(
        i_data_bus[294]), .B2(n9584), .ZN(n9510) );
  ND4D1BWP30P140LVT U10098 ( .A1(n9513), .A2(n9512), .A3(n9511), .A4(n9510), 
        .ZN(n9514) );
  NR4D0BWP30P140LVT U10099 ( .A1(n9517), .A2(n9516), .A3(n9515), .A4(n9514), 
        .ZN(n9518) );
  ND4D4BWP30P140LVT U10100 ( .A1(n9521), .A2(n9520), .A3(n9519), .A4(n9518), 
        .ZN(o_data_bus[230]) );
  AOI22D1BWP30P140LVT U10101 ( .A1(i_data_bus[4]), .A2(n9553), .B1(
        i_data_bus[836]), .B2(n9557), .ZN(n9545) );
  AOI22D1BWP30P140LVT U10102 ( .A1(i_data_bus[740]), .A2(n9546), .B1(
        i_data_bus[868]), .B2(n9556), .ZN(n9544) );
  AOI22D1BWP30P140LVT U10103 ( .A1(i_data_bus[932]), .A2(n9587), .B1(
        i_data_bus[324]), .B2(n9570), .ZN(n9543) );
  AOI22D1BWP30P140LVT U10104 ( .A1(i_data_bus[708]), .A2(n9554), .B1(
        i_data_bus[676]), .B2(n9559), .ZN(n9525) );
  AOI22D1BWP30P140LVT U10105 ( .A1(i_data_bus[772]), .A2(n9547), .B1(
        i_data_bus[804]), .B2(n9552), .ZN(n9524) );
  AOI22D1BWP30P140LVT U10106 ( .A1(i_data_bus[68]), .A2(n9549), .B1(
        i_data_bus[36]), .B2(n9548), .ZN(n9523) );
  AOI22D1BWP30P140LVT U10107 ( .A1(i_data_bus[100]), .A2(n9555), .B1(
        i_data_bus[644]), .B2(n9558), .ZN(n9522) );
  ND4D1BWP30P140LVT U10108 ( .A1(n9525), .A2(n9524), .A3(n9523), .A4(n9522), 
        .ZN(n9541) );
  MOAI22D1BWP30P140LVT U10109 ( .A1(n9527), .A2(n9526), .B1(i_data_bus[196]), 
        .B2(n9550), .ZN(n9540) );
  AOI22D1BWP30P140LVT U10110 ( .A1(i_data_bus[228]), .A2(n9568), .B1(
        i_data_bus[164]), .B2(n9583), .ZN(n9531) );
  AOI22D1BWP30P140LVT U10111 ( .A1(i_data_bus[996]), .A2(n9571), .B1(
        i_data_bus[484]), .B2(n9580), .ZN(n9530) );
  AOI22D1BWP30P140LVT U10112 ( .A1(i_data_bus[548]), .A2(n9575), .B1(
        i_data_bus[580]), .B2(n9572), .ZN(n9529) );
  AOI22D1BWP30P140LVT U10113 ( .A1(i_data_bus[612]), .A2(n9574), .B1(
        i_data_bus[516]), .B2(n9573), .ZN(n9528) );
  ND4D1BWP30P140LVT U10114 ( .A1(n9531), .A2(n9530), .A3(n9529), .A4(n9528), 
        .ZN(n9539) );
  AOI22D1BWP30P140LVT U10115 ( .A1(i_data_bus[964]), .A2(n9551), .B1(
        i_data_bus[356]), .B2(n9569), .ZN(n9537) );
  AOI22D1BWP30P140LVT U10116 ( .A1(i_data_bus[900]), .A2(n9581), .B1(
        i_data_bus[420]), .B2(n9532), .ZN(n9536) );
  AOI22D1BWP30P140LVT U10117 ( .A1(i_data_bus[292]), .A2(n9584), .B1(
        i_data_bus[388]), .B2(n9585), .ZN(n9535) );
  AOI22D1BWP30P140LVT U10118 ( .A1(i_data_bus[132]), .A2(n9533), .B1(
        i_data_bus[260]), .B2(n9586), .ZN(n9534) );
  ND4D1BWP30P140LVT U10119 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), 
        .ZN(n9538) );
  NR4D0BWP30P140LVT U10120 ( .A1(n9541), .A2(n9540), .A3(n9539), .A4(n9538), 
        .ZN(n9542) );
  ND4D4BWP30P140LVT U10121 ( .A1(n9545), .A2(n9544), .A3(n9543), .A4(n9542), 
        .ZN(o_data_bus[228]) );
  AOI22D1BWP30P140LVT U10122 ( .A1(i_data_bus[771]), .A2(n9547), .B1(
        i_data_bus[739]), .B2(n9546), .ZN(n9599) );
  AOI22D1BWP30P140LVT U10123 ( .A1(i_data_bus[67]), .A2(n9549), .B1(
        i_data_bus[35]), .B2(n9548), .ZN(n9598) );
  AOI22D1BWP30P140LVT U10124 ( .A1(i_data_bus[963]), .A2(n9551), .B1(
        i_data_bus[195]), .B2(n9550), .ZN(n9597) );
  AOI22D1BWP30P140LVT U10125 ( .A1(i_data_bus[3]), .A2(n9553), .B1(
        i_data_bus[803]), .B2(n9552), .ZN(n9563) );
  AOI22D1BWP30P140LVT U10126 ( .A1(i_data_bus[99]), .A2(n9555), .B1(
        i_data_bus[707]), .B2(n9554), .ZN(n9562) );
  AOI22D1BWP30P140LVT U10127 ( .A1(i_data_bus[835]), .A2(n9557), .B1(
        i_data_bus[867]), .B2(n9556), .ZN(n9561) );
  AOI22D1BWP30P140LVT U10128 ( .A1(i_data_bus[675]), .A2(n9559), .B1(
        i_data_bus[643]), .B2(n9558), .ZN(n9560) );
  ND4D1BWP30P140LVT U10129 ( .A1(n9563), .A2(n9562), .A3(n9561), .A4(n9560), 
        .ZN(n9595) );
  OAI22D1BWP30P140LVT U10130 ( .A1(n9567), .A2(n9566), .B1(n9565), .B2(n9564), 
        .ZN(n9594) );
  AOI22D1BWP30P140LVT U10131 ( .A1(i_data_bus[355]), .A2(n9569), .B1(
        i_data_bus[227]), .B2(n9568), .ZN(n9579) );
  AOI22D1BWP30P140LVT U10132 ( .A1(i_data_bus[995]), .A2(n9571), .B1(
        i_data_bus[323]), .B2(n9570), .ZN(n9578) );
  AOI22D1BWP30P140LVT U10133 ( .A1(i_data_bus[515]), .A2(n9573), .B1(
        i_data_bus[579]), .B2(n9572), .ZN(n9577) );
  AOI22D1BWP30P140LVT U10134 ( .A1(i_data_bus[547]), .A2(n9575), .B1(
        i_data_bus[611]), .B2(n9574), .ZN(n9576) );
  ND4D1BWP30P140LVT U10135 ( .A1(n9579), .A2(n9578), .A3(n9577), .A4(n9576), 
        .ZN(n9593) );
  AOI22D1BWP30P140LVT U10136 ( .A1(i_data_bus[899]), .A2(n9581), .B1(
        i_data_bus[483]), .B2(n9580), .ZN(n9591) );
  AOI22D1BWP30P140LVT U10137 ( .A1(i_data_bus[163]), .A2(n9583), .B1(
        i_data_bus[451]), .B2(n9582), .ZN(n9590) );
  AOI22D1BWP30P140LVT U10138 ( .A1(i_data_bus[387]), .A2(n9585), .B1(
        i_data_bus[291]), .B2(n9584), .ZN(n9589) );
  AOI22D1BWP30P140LVT U10139 ( .A1(i_data_bus[931]), .A2(n9587), .B1(
        i_data_bus[259]), .B2(n9586), .ZN(n9588) );
  ND4D1BWP30P140LVT U10140 ( .A1(n9591), .A2(n9590), .A3(n9589), .A4(n9588), 
        .ZN(n9592) );
  NR4D0BWP30P140LVT U10141 ( .A1(n9595), .A2(n9594), .A3(n9593), .A4(n9592), 
        .ZN(n9596) );
  ND4D4BWP30P140LVT U10142 ( .A1(n9599), .A2(n9598), .A3(n9597), .A4(n9596), 
        .ZN(o_data_bus[227]) );
  AOI22D1BWP30P140LVT U10143 ( .A1(i_data_bus[59]), .A2(n9670), .B1(
        i_data_bus[251]), .B2(n9671), .ZN(n9621) );
  AOI22D1BWP30P140LVT U10144 ( .A1(i_data_bus[923]), .A2(n9682), .B1(
        i_data_bus[155]), .B2(n9681), .ZN(n9620) );
  AOI22D1BWP30P140LVT U10145 ( .A1(i_data_bus[827]), .A2(n9674), .B1(
        i_data_bus[315]), .B2(n9655), .ZN(n9619) );
  AOI22D1BWP30P140LVT U10146 ( .A1(i_data_bus[123]), .A2(n9680), .B1(
        i_data_bus[187]), .B2(n9675), .ZN(n9603) );
  AOI22D1BWP30P140LVT U10147 ( .A1(i_data_bus[1019]), .A2(n9677), .B1(
        i_data_bus[27]), .B2(n9676), .ZN(n9602) );
  AOI22D1BWP30P140LVT U10148 ( .A1(i_data_bus[91]), .A2(n9672), .B1(
        i_data_bus[219]), .B2(n9679), .ZN(n9601) );
  AOI22D1BWP30P140LVT U10149 ( .A1(i_data_bus[987]), .A2(n9678), .B1(
        i_data_bus[955]), .B2(n9669), .ZN(n9600) );
  ND4D1BWP30P140LVT U10150 ( .A1(n9603), .A2(n9602), .A3(n9601), .A4(n9600), 
        .ZN(n9617) );
  MOAI22D1BWP30P140LVT U10151 ( .A1(n9605), .A2(n9604), .B1(i_data_bus[891]), 
        .B2(n9710), .ZN(n9616) );
  AOI22D1BWP30P140LVT U10152 ( .A1(i_data_bus[731]), .A2(n9704), .B1(
        i_data_bus[667]), .B2(n9707), .ZN(n9609) );
  AOI22D1BWP30P140LVT U10153 ( .A1(i_data_bus[763]), .A2(n9706), .B1(
        i_data_bus[347]), .B2(n9692), .ZN(n9608) );
  AOI22D1BWP30P140LVT U10154 ( .A1(i_data_bus[571]), .A2(n9695), .B1(
        i_data_bus[635]), .B2(n9696), .ZN(n9607) );
  AOI22D1BWP30P140LVT U10155 ( .A1(i_data_bus[603]), .A2(n9697), .B1(
        i_data_bus[539]), .B2(n9698), .ZN(n9606) );
  ND4D1BWP30P140LVT U10156 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), 
        .ZN(n9615) );
  AOI22D1BWP30P140LVT U10157 ( .A1(i_data_bus[443]), .A2(n9709), .B1(
        i_data_bus[699]), .B2(n9705), .ZN(n9613) );
  AOI22D1BWP30P140LVT U10158 ( .A1(i_data_bus[795]), .A2(n9673), .B1(
        i_data_bus[475]), .B2(n9703), .ZN(n9612) );
  AOI22D1BWP30P140LVT U10159 ( .A1(i_data_bus[507]), .A2(n9656), .B1(
        i_data_bus[283]), .B2(n9694), .ZN(n9611) );
  AOI22D1BWP30P140LVT U10160 ( .A1(i_data_bus[411]), .A2(n9708), .B1(
        i_data_bus[859]), .B2(n9693), .ZN(n9610) );
  ND4D1BWP30P140LVT U10161 ( .A1(n9613), .A2(n9612), .A3(n9611), .A4(n9610), 
        .ZN(n9614) );
  NR4D0BWP30P140LVT U10162 ( .A1(n9617), .A2(n9616), .A3(n9615), .A4(n9614), 
        .ZN(n9618) );
  ND4D4BWP30P140LVT U10163 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), 
        .ZN(o_data_bus[27]) );
  AOI22D1BWP30P140LVT U10164 ( .A1(i_data_bus[90]), .A2(n9672), .B1(
        i_data_bus[986]), .B2(n9678), .ZN(n9644) );
  AOI22D1BWP30P140LVT U10165 ( .A1(i_data_bus[1018]), .A2(n9677), .B1(
        i_data_bus[154]), .B2(n9681), .ZN(n9643) );
  AOI22D1BWP30P140LVT U10166 ( .A1(i_data_bus[442]), .A2(n9709), .B1(
        i_data_bus[698]), .B2(n9705), .ZN(n9642) );
  AOI22D1BWP30P140LVT U10167 ( .A1(i_data_bus[922]), .A2(n9682), .B1(
        i_data_bus[250]), .B2(n9671), .ZN(n9625) );
  AOI22D1BWP30P140LVT U10168 ( .A1(i_data_bus[954]), .A2(n9669), .B1(
        i_data_bus[186]), .B2(n9675), .ZN(n9624) );
  AOI22D1BWP30P140LVT U10169 ( .A1(i_data_bus[26]), .A2(n9676), .B1(
        i_data_bus[58]), .B2(n9670), .ZN(n9623) );
  AOI22D1BWP30P140LVT U10170 ( .A1(i_data_bus[122]), .A2(n9680), .B1(
        i_data_bus[218]), .B2(n9679), .ZN(n9622) );
  ND4D1BWP30P140LVT U10171 ( .A1(n9625), .A2(n9624), .A3(n9623), .A4(n9622), 
        .ZN(n9640) );
  OAI22D1BWP30P140LVT U10172 ( .A1(n9628), .A2(n9689), .B1(n9627), .B2(n9626), 
        .ZN(n9639) );
  AOI22D1BWP30P140LVT U10173 ( .A1(i_data_bus[826]), .A2(n9674), .B1(
        i_data_bus[890]), .B2(n9710), .ZN(n9632) );
  AOI22D1BWP30P140LVT U10174 ( .A1(i_data_bus[346]), .A2(n9692), .B1(
        i_data_bus[762]), .B2(n9706), .ZN(n9631) );
  AOI22D1BWP30P140LVT U10175 ( .A1(i_data_bus[538]), .A2(n9698), .B1(
        i_data_bus[570]), .B2(n9695), .ZN(n9630) );
  AOI22D1BWP30P140LVT U10176 ( .A1(i_data_bus[602]), .A2(n9697), .B1(
        i_data_bus[634]), .B2(n9696), .ZN(n9629) );
  ND4D1BWP30P140LVT U10177 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), 
        .ZN(n9638) );
  AOI22D1BWP30P140LVT U10178 ( .A1(i_data_bus[858]), .A2(n9693), .B1(
        i_data_bus[730]), .B2(n9704), .ZN(n9636) );
  AOI22D1BWP30P140LVT U10179 ( .A1(i_data_bus[666]), .A2(n9707), .B1(
        i_data_bus[474]), .B2(n9703), .ZN(n9635) );
  AOI22D1BWP30P140LVT U10180 ( .A1(i_data_bus[314]), .A2(n9655), .B1(
        i_data_bus[378]), .B2(n9691), .ZN(n9634) );
  AOI22D1BWP30P140LVT U10181 ( .A1(i_data_bus[282]), .A2(n9694), .B1(
        i_data_bus[794]), .B2(n9673), .ZN(n9633) );
  ND4D1BWP30P140LVT U10182 ( .A1(n9636), .A2(n9635), .A3(n9634), .A4(n9633), 
        .ZN(n9637) );
  NR4D0BWP30P140LVT U10183 ( .A1(n9640), .A2(n9639), .A3(n9638), .A4(n9637), 
        .ZN(n9641) );
  ND4D4BWP30P140LVT U10184 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), 
        .ZN(o_data_bus[26]) );
  AOI22D1BWP30P140LVT U10185 ( .A1(i_data_bus[907]), .A2(n9682), .B1(
        i_data_bus[971]), .B2(n9678), .ZN(n9668) );
  AOI22D1BWP30P140LVT U10186 ( .A1(i_data_bus[1003]), .A2(n9677), .B1(
        i_data_bus[75]), .B2(n9672), .ZN(n9667) );
  AOI22D1BWP30P140LVT U10187 ( .A1(i_data_bus[875]), .A2(n9710), .B1(
        i_data_bus[843]), .B2(n9693), .ZN(n9666) );
  AOI22D1BWP30P140LVT U10188 ( .A1(i_data_bus[107]), .A2(n9680), .B1(
        i_data_bus[203]), .B2(n9679), .ZN(n9648) );
  AOI22D1BWP30P140LVT U10189 ( .A1(i_data_bus[939]), .A2(n9669), .B1(
        i_data_bus[11]), .B2(n9676), .ZN(n9647) );
  AOI22D1BWP30P140LVT U10190 ( .A1(i_data_bus[171]), .A2(n9675), .B1(
        i_data_bus[235]), .B2(n9671), .ZN(n9646) );
  AOI22D1BWP30P140LVT U10191 ( .A1(i_data_bus[43]), .A2(n9670), .B1(
        i_data_bus[139]), .B2(n9681), .ZN(n9645) );
  ND4D1BWP30P140LVT U10192 ( .A1(n9648), .A2(n9647), .A3(n9646), .A4(n9645), 
        .ZN(n9664) );
  MOAI22D1BWP30P140LVT U10193 ( .A1(n9650), .A2(n9649), .B1(i_data_bus[747]), 
        .B2(n9706), .ZN(n9663) );
  AOI22D1BWP30P140LVT U10194 ( .A1(i_data_bus[651]), .A2(n9707), .B1(
        i_data_bus[683]), .B2(n9705), .ZN(n9654) );
  AOI22D1BWP30P140LVT U10195 ( .A1(i_data_bus[427]), .A2(n9709), .B1(
        i_data_bus[715]), .B2(n9704), .ZN(n9653) );
  AOI22D1BWP30P140LVT U10196 ( .A1(i_data_bus[619]), .A2(n9696), .B1(
        i_data_bus[587]), .B2(n9697), .ZN(n9652) );
  AOI22D1BWP30P140LVT U10197 ( .A1(i_data_bus[523]), .A2(n9698), .B1(
        i_data_bus[555]), .B2(n9695), .ZN(n9651) );
  ND4D1BWP30P140LVT U10198 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), 
        .ZN(n9662) );
  AOI22D1BWP30P140LVT U10199 ( .A1(i_data_bus[395]), .A2(n9708), .B1(
        i_data_bus[811]), .B2(n9674), .ZN(n9660) );
  AOI22D1BWP30P140LVT U10200 ( .A1(i_data_bus[363]), .A2(n9691), .B1(
        i_data_bus[267]), .B2(n9694), .ZN(n9659) );
  AOI22D1BWP30P140LVT U10201 ( .A1(i_data_bus[779]), .A2(n9673), .B1(
        i_data_bus[299]), .B2(n9655), .ZN(n9658) );
  AOI22D1BWP30P140LVT U10202 ( .A1(i_data_bus[491]), .A2(n9656), .B1(
        i_data_bus[331]), .B2(n9692), .ZN(n9657) );
  ND4D1BWP30P140LVT U10203 ( .A1(n9660), .A2(n9659), .A3(n9658), .A4(n9657), 
        .ZN(n9661) );
  NR4D0BWP30P140LVT U10204 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), 
        .ZN(n9665) );
  ND4D4BWP30P140LVT U10205 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), 
        .ZN(o_data_bus[11]) );
  AOI22D1BWP30P140LVT U10206 ( .A1(i_data_bus[41]), .A2(n9670), .B1(
        i_data_bus[937]), .B2(n9669), .ZN(n9722) );
  AOI22D1BWP30P140LVT U10207 ( .A1(i_data_bus[73]), .A2(n9672), .B1(
        i_data_bus[233]), .B2(n9671), .ZN(n9721) );
  AOI22D1BWP30P140LVT U10208 ( .A1(i_data_bus[809]), .A2(n9674), .B1(
        i_data_bus[777]), .B2(n9673), .ZN(n9720) );
  AOI22D1BWP30P140LVT U10209 ( .A1(i_data_bus[9]), .A2(n9676), .B1(
        i_data_bus[169]), .B2(n9675), .ZN(n9686) );
  AOI22D1BWP30P140LVT U10210 ( .A1(i_data_bus[969]), .A2(n9678), .B1(
        i_data_bus[1001]), .B2(n9677), .ZN(n9685) );
  AOI22D1BWP30P140LVT U10211 ( .A1(i_data_bus[105]), .A2(n9680), .B1(
        i_data_bus[201]), .B2(n9679), .ZN(n9684) );
  AOI22D1BWP30P140LVT U10212 ( .A1(i_data_bus[905]), .A2(n9682), .B1(
        i_data_bus[137]), .B2(n9681), .ZN(n9683) );
  ND4D1BWP30P140LVT U10213 ( .A1(n9686), .A2(n9685), .A3(n9684), .A4(n9683), 
        .ZN(n9718) );
  OAI22D1BWP30P140LVT U10214 ( .A1(n9690), .A2(n9689), .B1(n9688), .B2(n9687), 
        .ZN(n9717) );
  AOI22D1BWP30P140LVT U10215 ( .A1(i_data_bus[329]), .A2(n9692), .B1(
        i_data_bus[361]), .B2(n9691), .ZN(n9702) );
  AOI22D1BWP30P140LVT U10216 ( .A1(i_data_bus[265]), .A2(n9694), .B1(
        i_data_bus[841]), .B2(n9693), .ZN(n9701) );
  AOI22D1BWP30P140LVT U10217 ( .A1(i_data_bus[617]), .A2(n9696), .B1(
        i_data_bus[553]), .B2(n9695), .ZN(n9700) );
  AOI22D1BWP30P140LVT U10218 ( .A1(i_data_bus[521]), .A2(n9698), .B1(
        i_data_bus[585]), .B2(n9697), .ZN(n9699) );
  ND4D1BWP30P140LVT U10219 ( .A1(n9702), .A2(n9701), .A3(n9700), .A4(n9699), 
        .ZN(n9716) );
  AOI22D1BWP30P140LVT U10220 ( .A1(i_data_bus[713]), .A2(n9704), .B1(
        i_data_bus[457]), .B2(n9703), .ZN(n9714) );
  AOI22D1BWP30P140LVT U10221 ( .A1(i_data_bus[745]), .A2(n9706), .B1(
        i_data_bus[681]), .B2(n9705), .ZN(n9713) );
  AOI22D1BWP30P140LVT U10222 ( .A1(i_data_bus[393]), .A2(n9708), .B1(
        i_data_bus[649]), .B2(n9707), .ZN(n9712) );
  AOI22D1BWP30P140LVT U10223 ( .A1(i_data_bus[873]), .A2(n9710), .B1(
        i_data_bus[425]), .B2(n9709), .ZN(n9711) );
  ND4D1BWP30P140LVT U10224 ( .A1(n9714), .A2(n9713), .A3(n9712), .A4(n9711), 
        .ZN(n9715) );
  NR4D0BWP30P140LVT U10225 ( .A1(n9718), .A2(n9717), .A3(n9716), .A4(n9715), 
        .ZN(n9719) );
  ND4D4BWP30P140LVT U10226 ( .A1(n9722), .A2(n9721), .A3(n9720), .A4(n9719), 
        .ZN(o_data_bus[9]) );
  ND4D1BWP30P140LVT U10227 ( .A1(n9726), .A2(n9725), .A3(n9724), .A4(n9723), 
        .ZN(n9727) );
  NR2D1BWP30P140LVT U10228 ( .A1(n9728), .A2(n9727), .ZN(n9732) );
  ND4D4BWP30P140LVT U10229 ( .A1(n9732), .A2(n9731), .A3(n9730), .A4(n9729), 
        .ZN(o_valid[2]) );
  INVD1BWP30P140LVT U10230 ( .I(n9753), .ZN(n9733) );
  NR3D0P7BWP30P140LVT U10231 ( .A1(n11703), .A2(n9734), .A3(n9733), .ZN(n12490) );
  INR3D0BWP30P140LVT U10232 ( .A1(i_cmd[52]), .B1(n11030), .B2(n9749), .ZN(
        n12495) );
  AOI22D1BWP30P140LVT U10233 ( .A1(i_data_bus[5]), .A2(n12490), .B1(
        i_data_bus[197]), .B2(n12495), .ZN(n9740) );
  NR3D0P7BWP30P140LVT U10234 ( .A1(n11717), .A2(n9735), .A3(n9755), .ZN(n12496) );
  AN3D1BWP30P140LVT U10235 ( .A1(i_cmd[20]), .A2(i_valid[2]), .A3(n9753), .Z(
        n12478) );
  AOI22D1BWP30P140LVT U10236 ( .A1(i_data_bus[997]), .A2(n12496), .B1(
        i_data_bus[69]), .B2(n12478), .ZN(n9739) );
  INR3D0BWP30P140LVT U10237 ( .A1(i_cmd[92]), .B1(n11731), .B2(n9750), .ZN(
        n12491) );
  INR3D0BWP30P140LVT U10238 ( .A1(i_cmd[76]), .B1(n11711), .B2(n9750), .ZN(
        n12505) );
  AOI22D1BWP30P140LVT U10239 ( .A1(i_data_bus[357]), .A2(n12491), .B1(
        i_data_bus[293]), .B2(n12505), .ZN(n9738) );
  NR3D0P7BWP30P140LVT U10240 ( .A1(n11713), .A2(n9736), .A3(n9754), .ZN(n12477) );
  INR3D0BWP30P140LVT U10241 ( .A1(i_cmd[60]), .B1(n11032), .B2(n9749), .ZN(
        n12493) );
  AOI22D1BWP30P140LVT U10242 ( .A1(i_data_bus[517]), .A2(n12477), .B1(
        i_data_bus[229]), .B2(n12493), .ZN(n9737) );
  ND4D1BWP30P140LVT U10243 ( .A1(n9740), .A2(n9739), .A3(n9738), .A4(n9737), 
        .ZN(n9772) );
  INR3D0BWP30P140LVT U10244 ( .A1(i_cmd[148]), .B1(n11733), .B2(n9754), .ZN(
        n12480) );
  INVD1BWP30P140LVT U10245 ( .I(i_cmd[100]), .ZN(n9741) );
  NR3D0P7BWP30P140LVT U10246 ( .A1(n11705), .A2(n9741), .A3(n9748), .ZN(n12506) );
  AOI22D1BWP30P140LVT U10247 ( .A1(i_data_bus[581]), .A2(n12480), .B1(
        i_data_bus[389]), .B2(n12506), .ZN(n9747) );
  AN3D1BWP30P140LVT U10248 ( .A1(i_cmd[28]), .A2(i_valid[3]), .A3(n9753), .Z(
        n12489) );
  INVD1BWP30P140LVT U10249 ( .I(i_cmd[36]), .ZN(n9742) );
  NR3D0P7BWP30P140LVT U10250 ( .A1(n11721), .A2(n9742), .A3(n9749), .ZN(n12502) );
  AOI22D1BWP30P140LVT U10251 ( .A1(i_data_bus[101]), .A2(n12489), .B1(
        i_data_bus[133]), .B2(n12502), .ZN(n9746) );
  INR3D0BWP30P140LVT U10252 ( .A1(i_cmd[116]), .B1(n11706), .B2(n9748), .ZN(
        n12507) );
  INR3D0BWP30P140LVT U10253 ( .A1(i_cmd[84]), .B1(n11700), .B2(n9750), .ZN(
        n12508) );
  AOI22D1BWP30P140LVT U10254 ( .A1(i_data_bus[453]), .A2(n12507), .B1(
        i_data_bus[325]), .B2(n12508), .ZN(n9745) );
  NR3D0P7BWP30P140LVT U10255 ( .A1(n11715), .A2(n9743), .A3(n9755), .ZN(n12482) );
  INR3D0BWP30P140LVT U10256 ( .A1(i_cmd[124]), .B1(n11719), .B2(n9748), .ZN(
        n12494) );
  AOI22D1BWP30P140LVT U10257 ( .A1(i_data_bus[965]), .A2(n12482), .B1(
        i_data_bus[485]), .B2(n12494), .ZN(n9744) );
  ND4D1BWP30P140LVT U10258 ( .A1(n9747), .A2(n9746), .A3(n9745), .A4(n9744), 
        .ZN(n9771) );
  INR3D0BWP30P140LVT U10259 ( .A1(i_cmd[156]), .B1(n11697), .B2(n9754), .ZN(
        n12504) );
  INR3D0BWP30P140LVT U10260 ( .A1(i_cmd[108]), .B1(n11698), .B2(n9748), .ZN(
        n12481) );
  AOI22D1BWP30P140LVT U10261 ( .A1(i_data_bus[613]), .A2(n12504), .B1(
        i_data_bus[421]), .B2(n12481), .ZN(n9760) );
  INR3D0BWP30P140LVT U10262 ( .A1(i_cmd[44]), .B1(n11023), .B2(n9749), .ZN(
        n12501) );
  NR3D0P7BWP30P140LVT U10263 ( .A1(n11728), .A2(n9751), .A3(n9750), .ZN(n12503) );
  AOI22D1BWP30P140LVT U10264 ( .A1(i_data_bus[165]), .A2(n12501), .B1(
        i_data_bus[261]), .B2(n12503), .ZN(n9759) );
  NR3D0P7BWP30P140LVT U10265 ( .A1(n11735), .A2(n9752), .A3(n9755), .ZN(n12484) );
  AN3D1BWP30P140LVT U10266 ( .A1(i_cmd[12]), .A2(i_valid[1]), .A3(n9753), .Z(
        n12483) );
  AOI22D1BWP30P140LVT U10267 ( .A1(i_data_bus[901]), .A2(n12484), .B1(
        i_data_bus[37]), .B2(n12483), .ZN(n9758) );
  INR3D0BWP30P140LVT U10268 ( .A1(i_cmd[140]), .B1(n11701), .B2(n9754), .ZN(
        n12479) );
  NR3D0P7BWP30P140LVT U10269 ( .A1(n11740), .A2(n9756), .A3(n9755), .ZN(n12492) );
  AOI22D1BWP30P140LVT U10270 ( .A1(i_data_bus[549]), .A2(n12479), .B1(
        i_data_bus[933]), .B2(n12492), .ZN(n9757) );
  ND4D1BWP30P140LVT U10271 ( .A1(n9760), .A2(n9759), .A3(n9758), .A4(n9757), 
        .ZN(n9770) );
  INR3D0BWP30P140LVT U10272 ( .A1(i_cmd[204]), .B1(n11751), .B2(n9762), .ZN(
        n12517) );
  INR3D0BWP30P140LVT U10273 ( .A1(i_cmd[180]), .B1(n11748), .B2(n9764), .ZN(
        n12519) );
  AOI22D1BWP30P140LVT U10274 ( .A1(i_data_bus[805]), .A2(n12517), .B1(
        i_data_bus[709]), .B2(n12519), .ZN(n9768) );
  INR3D0BWP30P140LVT U10275 ( .A1(i_cmd[172]), .B1(n11756), .B2(n9764), .ZN(
        n12515) );
  INR3D0BWP30P140LVT U10276 ( .A1(i_cmd[212]), .B1(n11745), .B2(n9762), .ZN(
        n12514) );
  AOI22D1BWP30P140LVT U10277 ( .A1(i_data_bus[677]), .A2(n12515), .B1(
        i_data_bus[837]), .B2(n12514), .ZN(n9767) );
  NR3D0P7BWP30P140LVT U10278 ( .A1(n11747), .A2(n9761), .A3(n9764), .ZN(n12520) );
  INR3D0BWP30P140LVT U10279 ( .A1(i_cmd[220]), .B1(n11749), .B2(n9762), .ZN(
        n12513) );
  AOI22D1BWP30P140LVT U10280 ( .A1(i_data_bus[645]), .A2(n12520), .B1(
        i_data_bus[869]), .B2(n12513), .ZN(n9766) );
  NR3D0P7BWP30P140LVT U10281 ( .A1(n11754), .A2(n9763), .A3(n9762), .ZN(n12516) );
  INR3D0BWP30P140LVT U10282 ( .A1(i_cmd[188]), .B1(n11750), .B2(n9764), .ZN(
        n12518) );
  AOI22D1BWP30P140LVT U10283 ( .A1(i_data_bus[773]), .A2(n12516), .B1(
        i_data_bus[741]), .B2(n12518), .ZN(n9765) );
  ND4D1BWP30P140LVT U10284 ( .A1(n9768), .A2(n9767), .A3(n9766), .A4(n9765), 
        .ZN(n9769) );
  OR4D1BWP30P140LVT U10285 ( .A1(n9772), .A2(n9771), .A3(n9770), .A4(n9769), 
        .Z(o_data_bus[133]) );
  AOI22D1BWP30P140LVT U10286 ( .A1(i_data_bus[902]), .A2(n12484), .B1(
        i_data_bus[166]), .B2(n12501), .ZN(n9776) );
  AOI22D1BWP30P140LVT U10287 ( .A1(i_data_bus[390]), .A2(n12506), .B1(
        i_data_bus[454]), .B2(n12507), .ZN(n9775) );
  AOI22D1BWP30P140LVT U10288 ( .A1(i_data_bus[582]), .A2(n12480), .B1(
        i_data_bus[550]), .B2(n12479), .ZN(n9774) );
  AOI22D1BWP30P140LVT U10289 ( .A1(i_data_bus[422]), .A2(n12481), .B1(
        i_data_bus[294]), .B2(n12505), .ZN(n9773) );
  ND4D1BWP30P140LVT U10290 ( .A1(n9776), .A2(n9775), .A3(n9774), .A4(n9773), 
        .ZN(n9792) );
  AOI22D1BWP30P140LVT U10291 ( .A1(i_data_bus[70]), .A2(n12478), .B1(
        i_data_bus[102]), .B2(n12489), .ZN(n9780) );
  AOI22D1BWP30P140LVT U10292 ( .A1(i_data_bus[358]), .A2(n12491), .B1(
        i_data_bus[198]), .B2(n12495), .ZN(n9779) );
  AOI22D1BWP30P140LVT U10293 ( .A1(i_data_bus[38]), .A2(n12483), .B1(
        i_data_bus[326]), .B2(n12508), .ZN(n9778) );
  AOI22D1BWP30P140LVT U10294 ( .A1(i_data_bus[934]), .A2(n12492), .B1(
        i_data_bus[486]), .B2(n12494), .ZN(n9777) );
  ND4D1BWP30P140LVT U10295 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), 
        .ZN(n9791) );
  AOI22D1BWP30P140LVT U10296 ( .A1(i_data_bus[6]), .A2(n12490), .B1(
        i_data_bus[518]), .B2(n12477), .ZN(n9784) );
  AOI22D1BWP30P140LVT U10297 ( .A1(i_data_bus[614]), .A2(n12504), .B1(
        i_data_bus[998]), .B2(n12496), .ZN(n9783) );
  AOI22D1BWP30P140LVT U10298 ( .A1(i_data_bus[966]), .A2(n12482), .B1(
        i_data_bus[262]), .B2(n12503), .ZN(n9782) );
  AOI22D1BWP30P140LVT U10299 ( .A1(i_data_bus[230]), .A2(n12493), .B1(
        i_data_bus[134]), .B2(n12502), .ZN(n9781) );
  ND4D1BWP30P140LVT U10300 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), 
        .ZN(n9790) );
  AOI22D1BWP30P140LVT U10301 ( .A1(i_data_bus[646]), .A2(n12520), .B1(
        i_data_bus[678]), .B2(n12515), .ZN(n9788) );
  AOI22D1BWP30P140LVT U10302 ( .A1(i_data_bus[870]), .A2(n12513), .B1(
        i_data_bus[838]), .B2(n12514), .ZN(n9787) );
  AOI22D1BWP30P140LVT U10303 ( .A1(i_data_bus[710]), .A2(n12519), .B1(
        i_data_bus[774]), .B2(n12516), .ZN(n9786) );
  AOI22D1BWP30P140LVT U10304 ( .A1(i_data_bus[806]), .A2(n12517), .B1(
        i_data_bus[742]), .B2(n12518), .ZN(n9785) );
  ND4D1BWP30P140LVT U10305 ( .A1(n9788), .A2(n9787), .A3(n9786), .A4(n9785), 
        .ZN(n9789) );
  OR4D1BWP30P140LVT U10306 ( .A1(n9792), .A2(n9791), .A3(n9790), .A4(n9789), 
        .Z(o_data_bus[134]) );
  AOI22D1BWP30P140LVT U10307 ( .A1(i_data_bus[967]), .A2(n12482), .B1(
        i_data_bus[359]), .B2(n12491), .ZN(n9796) );
  AOI22D1BWP30P140LVT U10308 ( .A1(i_data_bus[615]), .A2(n12504), .B1(
        i_data_bus[519]), .B2(n12477), .ZN(n9795) );
  AOI22D1BWP30P140LVT U10309 ( .A1(i_data_bus[935]), .A2(n12492), .B1(
        i_data_bus[135]), .B2(n12502), .ZN(n9794) );
  AOI22D1BWP30P140LVT U10310 ( .A1(i_data_bus[487]), .A2(n12494), .B1(
        i_data_bus[167]), .B2(n12501), .ZN(n9793) );
  ND4D1BWP30P140LVT U10311 ( .A1(n9796), .A2(n9795), .A3(n9794), .A4(n9793), 
        .ZN(n9812) );
  AOI22D1BWP30P140LVT U10312 ( .A1(i_data_bus[103]), .A2(n12489), .B1(
        i_data_bus[7]), .B2(n12490), .ZN(n9800) );
  AOI22D1BWP30P140LVT U10313 ( .A1(i_data_bus[39]), .A2(n12483), .B1(
        i_data_bus[199]), .B2(n12495), .ZN(n9799) );
  AOI22D1BWP30P140LVT U10314 ( .A1(i_data_bus[263]), .A2(n12503), .B1(
        i_data_bus[295]), .B2(n12505), .ZN(n9798) );
  AOI22D1BWP30P140LVT U10315 ( .A1(i_data_bus[903]), .A2(n12484), .B1(
        i_data_bus[231]), .B2(n12493), .ZN(n9797) );
  ND4D1BWP30P140LVT U10316 ( .A1(n9800), .A2(n9799), .A3(n9798), .A4(n9797), 
        .ZN(n9811) );
  AOI22D1BWP30P140LVT U10317 ( .A1(i_data_bus[999]), .A2(n12496), .B1(
        i_data_bus[71]), .B2(n12478), .ZN(n9804) );
  AOI22D1BWP30P140LVT U10318 ( .A1(i_data_bus[423]), .A2(n12481), .B1(
        i_data_bus[327]), .B2(n12508), .ZN(n9803) );
  AOI22D1BWP30P140LVT U10319 ( .A1(i_data_bus[455]), .A2(n12507), .B1(
        i_data_bus[391]), .B2(n12506), .ZN(n9802) );
  AOI22D1BWP30P140LVT U10320 ( .A1(i_data_bus[551]), .A2(n12479), .B1(
        i_data_bus[583]), .B2(n12480), .ZN(n9801) );
  ND4D1BWP30P140LVT U10321 ( .A1(n9804), .A2(n9803), .A3(n9802), .A4(n9801), 
        .ZN(n9810) );
  AOI22D1BWP30P140LVT U10322 ( .A1(i_data_bus[871]), .A2(n12513), .B1(
        i_data_bus[711]), .B2(n12519), .ZN(n9808) );
  AOI22D1BWP30P140LVT U10323 ( .A1(i_data_bus[839]), .A2(n12514), .B1(
        i_data_bus[647]), .B2(n12520), .ZN(n9807) );
  AOI22D1BWP30P140LVT U10324 ( .A1(i_data_bus[679]), .A2(n12515), .B1(
        i_data_bus[775]), .B2(n12516), .ZN(n9806) );
  AOI22D1BWP30P140LVT U10325 ( .A1(i_data_bus[807]), .A2(n12517), .B1(
        i_data_bus[743]), .B2(n12518), .ZN(n9805) );
  ND4D1BWP30P140LVT U10326 ( .A1(n9808), .A2(n9807), .A3(n9806), .A4(n9805), 
        .ZN(n9809) );
  OR4D1BWP30P140LVT U10327 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), 
        .Z(o_data_bus[135]) );
  AOI22D1BWP30P140LVT U10328 ( .A1(i_data_bus[424]), .A2(n12481), .B1(
        i_data_bus[360]), .B2(n12491), .ZN(n9816) );
  AOI22D1BWP30P140LVT U10329 ( .A1(i_data_bus[552]), .A2(n12479), .B1(
        i_data_bus[40]), .B2(n12483), .ZN(n9815) );
  AOI22D1BWP30P140LVT U10330 ( .A1(i_data_bus[104]), .A2(n12489), .B1(
        i_data_bus[1000]), .B2(n12496), .ZN(n9814) );
  AOI22D1BWP30P140LVT U10331 ( .A1(i_data_bus[520]), .A2(n12477), .B1(
        i_data_bus[72]), .B2(n12478), .ZN(n9813) );
  ND4D1BWP30P140LVT U10332 ( .A1(n9816), .A2(n9815), .A3(n9814), .A4(n9813), 
        .ZN(n9832) );
  AOI22D1BWP30P140LVT U10333 ( .A1(i_data_bus[936]), .A2(n12492), .B1(
        i_data_bus[328]), .B2(n12508), .ZN(n9820) );
  AOI22D1BWP30P140LVT U10334 ( .A1(i_data_bus[8]), .A2(n12490), .B1(
        i_data_bus[488]), .B2(n12494), .ZN(n9819) );
  AOI22D1BWP30P140LVT U10335 ( .A1(i_data_bus[968]), .A2(n12482), .B1(
        i_data_bus[296]), .B2(n12505), .ZN(n9818) );
  AOI22D1BWP30P140LVT U10336 ( .A1(i_data_bus[264]), .A2(n12503), .B1(
        i_data_bus[136]), .B2(n12502), .ZN(n9817) );
  ND4D1BWP30P140LVT U10337 ( .A1(n9820), .A2(n9819), .A3(n9818), .A4(n9817), 
        .ZN(n9831) );
  AOI22D1BWP30P140LVT U10338 ( .A1(i_data_bus[456]), .A2(n12507), .B1(
        i_data_bus[200]), .B2(n12495), .ZN(n9824) );
  AOI22D1BWP30P140LVT U10339 ( .A1(i_data_bus[584]), .A2(n12480), .B1(
        i_data_bus[392]), .B2(n12506), .ZN(n9823) );
  AOI22D1BWP30P140LVT U10340 ( .A1(i_data_bus[904]), .A2(n12484), .B1(
        i_data_bus[168]), .B2(n12501), .ZN(n9822) );
  AOI22D1BWP30P140LVT U10341 ( .A1(i_data_bus[616]), .A2(n12504), .B1(
        i_data_bus[232]), .B2(n12493), .ZN(n9821) );
  ND4D1BWP30P140LVT U10342 ( .A1(n9824), .A2(n9823), .A3(n9822), .A4(n9821), 
        .ZN(n9830) );
  AOI22D1BWP30P140LVT U10343 ( .A1(i_data_bus[680]), .A2(n12515), .B1(
        i_data_bus[872]), .B2(n12513), .ZN(n9828) );
  AOI22D1BWP30P140LVT U10344 ( .A1(i_data_bus[840]), .A2(n12514), .B1(
        i_data_bus[776]), .B2(n12516), .ZN(n9827) );
  AOI22D1BWP30P140LVT U10345 ( .A1(i_data_bus[744]), .A2(n12518), .B1(
        i_data_bus[808]), .B2(n12517), .ZN(n9826) );
  AOI22D1BWP30P140LVT U10346 ( .A1(i_data_bus[712]), .A2(n12519), .B1(
        i_data_bus[648]), .B2(n12520), .ZN(n9825) );
  ND4D1BWP30P140LVT U10347 ( .A1(n9828), .A2(n9827), .A3(n9826), .A4(n9825), 
        .ZN(n9829) );
  OR4D1BWP30P140LVT U10348 ( .A1(n9832), .A2(n9831), .A3(n9830), .A4(n9829), 
        .Z(o_data_bus[136]) );
  AOI22D1BWP30P140LVT U10349 ( .A1(i_data_bus[553]), .A2(n12479), .B1(
        i_data_bus[361]), .B2(n12491), .ZN(n9836) );
  AOI22D1BWP30P140LVT U10350 ( .A1(i_data_bus[201]), .A2(n12495), .B1(
        i_data_bus[329]), .B2(n12508), .ZN(n9835) );
  AOI22D1BWP30P140LVT U10351 ( .A1(i_data_bus[233]), .A2(n12493), .B1(
        i_data_bus[137]), .B2(n12502), .ZN(n9834) );
  AOI22D1BWP30P140LVT U10352 ( .A1(i_data_bus[297]), .A2(n12505), .B1(
        i_data_bus[457]), .B2(n12507), .ZN(n9833) );
  ND4D1BWP30P140LVT U10353 ( .A1(n9836), .A2(n9835), .A3(n9834), .A4(n9833), 
        .ZN(n9852) );
  AOI22D1BWP30P140LVT U10354 ( .A1(i_data_bus[9]), .A2(n12490), .B1(
        i_data_bus[585]), .B2(n12480), .ZN(n9840) );
  AOI22D1BWP30P140LVT U10355 ( .A1(i_data_bus[73]), .A2(n12478), .B1(
        i_data_bus[969]), .B2(n12482), .ZN(n9839) );
  AOI22D1BWP30P140LVT U10356 ( .A1(i_data_bus[489]), .A2(n12494), .B1(
        i_data_bus[393]), .B2(n12506), .ZN(n9838) );
  AOI22D1BWP30P140LVT U10357 ( .A1(i_data_bus[105]), .A2(n12489), .B1(
        i_data_bus[1001]), .B2(n12496), .ZN(n9837) );
  ND4D1BWP30P140LVT U10358 ( .A1(n9840), .A2(n9839), .A3(n9838), .A4(n9837), 
        .ZN(n9851) );
  AOI22D1BWP30P140LVT U10359 ( .A1(i_data_bus[41]), .A2(n12483), .B1(
        i_data_bus[265]), .B2(n12503), .ZN(n9844) );
  AOI22D1BWP30P140LVT U10360 ( .A1(i_data_bus[905]), .A2(n12484), .B1(
        i_data_bus[937]), .B2(n12492), .ZN(n9843) );
  AOI22D1BWP30P140LVT U10361 ( .A1(i_data_bus[521]), .A2(n12477), .B1(
        i_data_bus[617]), .B2(n12504), .ZN(n9842) );
  AOI22D1BWP30P140LVT U10362 ( .A1(i_data_bus[169]), .A2(n12501), .B1(
        i_data_bus[425]), .B2(n12481), .ZN(n9841) );
  ND4D1BWP30P140LVT U10363 ( .A1(n9844), .A2(n9843), .A3(n9842), .A4(n9841), 
        .ZN(n9850) );
  AOI22D1BWP30P140LVT U10364 ( .A1(i_data_bus[745]), .A2(n12518), .B1(
        i_data_bus[873]), .B2(n12513), .ZN(n9848) );
  AOI22D1BWP30P140LVT U10365 ( .A1(i_data_bus[681]), .A2(n12515), .B1(
        i_data_bus[649]), .B2(n12520), .ZN(n9847) );
  AOI22D1BWP30P140LVT U10366 ( .A1(i_data_bus[777]), .A2(n12516), .B1(
        i_data_bus[841]), .B2(n12514), .ZN(n9846) );
  AOI22D1BWP30P140LVT U10367 ( .A1(i_data_bus[713]), .A2(n12519), .B1(
        i_data_bus[809]), .B2(n12517), .ZN(n9845) );
  ND4D1BWP30P140LVT U10368 ( .A1(n9848), .A2(n9847), .A3(n9846), .A4(n9845), 
        .ZN(n9849) );
  OR4D1BWP30P140LVT U10369 ( .A1(n9852), .A2(n9851), .A3(n9850), .A4(n9849), 
        .Z(o_data_bus[137]) );
  AOI22D1BWP30P140LVT U10370 ( .A1(i_data_bus[906]), .A2(n12484), .B1(
        i_data_bus[522]), .B2(n12477), .ZN(n9856) );
  AOI22D1BWP30P140LVT U10371 ( .A1(i_data_bus[618]), .A2(n12504), .B1(
        i_data_bus[426]), .B2(n12481), .ZN(n9855) );
  AOI22D1BWP30P140LVT U10372 ( .A1(i_data_bus[970]), .A2(n12482), .B1(
        i_data_bus[266]), .B2(n12503), .ZN(n9854) );
  AOI22D1BWP30P140LVT U10373 ( .A1(i_data_bus[106]), .A2(n12489), .B1(
        i_data_bus[586]), .B2(n12480), .ZN(n9853) );
  ND4D1BWP30P140LVT U10374 ( .A1(n9856), .A2(n9855), .A3(n9854), .A4(n9853), 
        .ZN(n9872) );
  AOI22D1BWP30P140LVT U10375 ( .A1(i_data_bus[74]), .A2(n12478), .B1(
        i_data_bus[394]), .B2(n12506), .ZN(n9860) );
  AOI22D1BWP30P140LVT U10376 ( .A1(i_data_bus[202]), .A2(n12495), .B1(
        i_data_bus[234]), .B2(n12493), .ZN(n9859) );
  AOI22D1BWP30P140LVT U10377 ( .A1(i_data_bus[554]), .A2(n12479), .B1(
        i_data_bus[298]), .B2(n12505), .ZN(n9858) );
  AOI22D1BWP30P140LVT U10378 ( .A1(i_data_bus[42]), .A2(n12483), .B1(
        i_data_bus[362]), .B2(n12491), .ZN(n9857) );
  ND4D1BWP30P140LVT U10379 ( .A1(n9860), .A2(n9859), .A3(n9858), .A4(n9857), 
        .ZN(n9871) );
  AOI22D1BWP30P140LVT U10380 ( .A1(i_data_bus[10]), .A2(n12490), .B1(
        i_data_bus[138]), .B2(n12502), .ZN(n9864) );
  AOI22D1BWP30P140LVT U10381 ( .A1(i_data_bus[1002]), .A2(n12496), .B1(
        i_data_bus[170]), .B2(n12501), .ZN(n9863) );
  AOI22D1BWP30P140LVT U10382 ( .A1(i_data_bus[330]), .A2(n12508), .B1(
        i_data_bus[458]), .B2(n12507), .ZN(n9862) );
  AOI22D1BWP30P140LVT U10383 ( .A1(i_data_bus[938]), .A2(n12492), .B1(
        i_data_bus[490]), .B2(n12494), .ZN(n9861) );
  ND4D1BWP30P140LVT U10384 ( .A1(n9864), .A2(n9863), .A3(n9862), .A4(n9861), 
        .ZN(n9870) );
  AOI22D1BWP30P140LVT U10385 ( .A1(i_data_bus[650]), .A2(n12520), .B1(
        i_data_bus[842]), .B2(n12514), .ZN(n9868) );
  AOI22D1BWP30P140LVT U10386 ( .A1(i_data_bus[778]), .A2(n12516), .B1(
        i_data_bus[874]), .B2(n12513), .ZN(n9867) );
  AOI22D1BWP30P140LVT U10387 ( .A1(i_data_bus[714]), .A2(n12519), .B1(
        i_data_bus[810]), .B2(n12517), .ZN(n9866) );
  AOI22D1BWP30P140LVT U10388 ( .A1(i_data_bus[746]), .A2(n12518), .B1(
        i_data_bus[682]), .B2(n12515), .ZN(n9865) );
  ND4D1BWP30P140LVT U10389 ( .A1(n9868), .A2(n9867), .A3(n9866), .A4(n9865), 
        .ZN(n9869) );
  OR4D1BWP30P140LVT U10390 ( .A1(n9872), .A2(n9871), .A3(n9870), .A4(n9869), 
        .Z(o_data_bus[138]) );
  AOI22D1BWP30P140LVT U10391 ( .A1(i_data_bus[523]), .A2(n12477), .B1(
        i_data_bus[235]), .B2(n12493), .ZN(n9876) );
  AOI22D1BWP30P140LVT U10392 ( .A1(i_data_bus[203]), .A2(n12495), .B1(
        i_data_bus[171]), .B2(n12501), .ZN(n9875) );
  AOI22D1BWP30P140LVT U10393 ( .A1(i_data_bus[971]), .A2(n12482), .B1(
        i_data_bus[587]), .B2(n12480), .ZN(n9874) );
  AOI22D1BWP30P140LVT U10394 ( .A1(i_data_bus[907]), .A2(n12484), .B1(
        i_data_bus[619]), .B2(n12504), .ZN(n9873) );
  ND4D1BWP30P140LVT U10395 ( .A1(n9876), .A2(n9875), .A3(n9874), .A4(n9873), 
        .ZN(n9892) );
  AOI22D1BWP30P140LVT U10396 ( .A1(i_data_bus[107]), .A2(n12489), .B1(
        i_data_bus[427]), .B2(n12481), .ZN(n9880) );
  AOI22D1BWP30P140LVT U10397 ( .A1(i_data_bus[75]), .A2(n12478), .B1(
        i_data_bus[139]), .B2(n12502), .ZN(n9879) );
  AOI22D1BWP30P140LVT U10398 ( .A1(i_data_bus[555]), .A2(n12479), .B1(
        i_data_bus[299]), .B2(n12505), .ZN(n9878) );
  AOI22D1BWP30P140LVT U10399 ( .A1(i_data_bus[939]), .A2(n12492), .B1(
        i_data_bus[267]), .B2(n12503), .ZN(n9877) );
  ND4D1BWP30P140LVT U10400 ( .A1(n9880), .A2(n9879), .A3(n9878), .A4(n9877), 
        .ZN(n9891) );
  AOI22D1BWP30P140LVT U10401 ( .A1(i_data_bus[43]), .A2(n12483), .B1(
        i_data_bus[363]), .B2(n12491), .ZN(n9884) );
  AOI22D1BWP30P140LVT U10402 ( .A1(i_data_bus[11]), .A2(n12490), .B1(
        i_data_bus[459]), .B2(n12507), .ZN(n9883) );
  AOI22D1BWP30P140LVT U10403 ( .A1(i_data_bus[1003]), .A2(n12496), .B1(
        i_data_bus[491]), .B2(n12494), .ZN(n9882) );
  AOI22D1BWP30P140LVT U10404 ( .A1(i_data_bus[395]), .A2(n12506), .B1(
        i_data_bus[331]), .B2(n12508), .ZN(n9881) );
  ND4D1BWP30P140LVT U10405 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), 
        .ZN(n9890) );
  AOI22D1BWP30P140LVT U10406 ( .A1(i_data_bus[811]), .A2(n12517), .B1(
        i_data_bus[779]), .B2(n12516), .ZN(n9888) );
  AOI22D1BWP30P140LVT U10407 ( .A1(i_data_bus[843]), .A2(n12514), .B1(
        i_data_bus[683]), .B2(n12515), .ZN(n9887) );
  AOI22D1BWP30P140LVT U10408 ( .A1(i_data_bus[651]), .A2(n12520), .B1(
        i_data_bus[715]), .B2(n12519), .ZN(n9886) );
  AOI22D1BWP30P140LVT U10409 ( .A1(i_data_bus[875]), .A2(n12513), .B1(
        i_data_bus[747]), .B2(n12518), .ZN(n9885) );
  ND4D1BWP30P140LVT U10410 ( .A1(n9888), .A2(n9887), .A3(n9886), .A4(n9885), 
        .ZN(n9889) );
  OR4D1BWP30P140LVT U10411 ( .A1(n9892), .A2(n9891), .A3(n9890), .A4(n9889), 
        .Z(o_data_bus[139]) );
  AOI22D1BWP30P140LVT U10412 ( .A1(i_data_bus[524]), .A2(n12477), .B1(
        i_data_bus[268]), .B2(n12503), .ZN(n9896) );
  AOI22D1BWP30P140LVT U10413 ( .A1(i_data_bus[460]), .A2(n12507), .B1(
        i_data_bus[332]), .B2(n12508), .ZN(n9895) );
  AOI22D1BWP30P140LVT U10414 ( .A1(i_data_bus[620]), .A2(n12504), .B1(
        i_data_bus[972]), .B2(n12482), .ZN(n9894) );
  AOI22D1BWP30P140LVT U10415 ( .A1(i_data_bus[492]), .A2(n12494), .B1(
        i_data_bus[172]), .B2(n12501), .ZN(n9893) );
  ND4D1BWP30P140LVT U10416 ( .A1(n9896), .A2(n9895), .A3(n9894), .A4(n9893), 
        .ZN(n9912) );
  AOI22D1BWP30P140LVT U10417 ( .A1(i_data_bus[76]), .A2(n12478), .B1(
        i_data_bus[204]), .B2(n12495), .ZN(n9900) );
  AOI22D1BWP30P140LVT U10418 ( .A1(i_data_bus[44]), .A2(n12483), .B1(
        i_data_bus[908]), .B2(n12484), .ZN(n9899) );
  AOI22D1BWP30P140LVT U10419 ( .A1(i_data_bus[12]), .A2(n12490), .B1(
        i_data_bus[396]), .B2(n12506), .ZN(n9898) );
  AOI22D1BWP30P140LVT U10420 ( .A1(i_data_bus[108]), .A2(n12489), .B1(
        i_data_bus[140]), .B2(n12502), .ZN(n9897) );
  ND4D1BWP30P140LVT U10421 ( .A1(n9900), .A2(n9899), .A3(n9898), .A4(n9897), 
        .ZN(n9911) );
  AOI22D1BWP30P140LVT U10422 ( .A1(i_data_bus[588]), .A2(n12480), .B1(
        i_data_bus[428]), .B2(n12481), .ZN(n9904) );
  AOI22D1BWP30P140LVT U10423 ( .A1(i_data_bus[556]), .A2(n12479), .B1(
        i_data_bus[364]), .B2(n12491), .ZN(n9903) );
  AOI22D1BWP30P140LVT U10424 ( .A1(i_data_bus[1004]), .A2(n12496), .B1(
        i_data_bus[300]), .B2(n12505), .ZN(n9902) );
  AOI22D1BWP30P140LVT U10425 ( .A1(i_data_bus[940]), .A2(n12492), .B1(
        i_data_bus[236]), .B2(n12493), .ZN(n9901) );
  ND4D1BWP30P140LVT U10426 ( .A1(n9904), .A2(n9903), .A3(n9902), .A4(n9901), 
        .ZN(n9910) );
  AOI22D1BWP30P140LVT U10427 ( .A1(i_data_bus[716]), .A2(n12519), .B1(
        i_data_bus[844]), .B2(n12514), .ZN(n9908) );
  AOI22D1BWP30P140LVT U10428 ( .A1(i_data_bus[780]), .A2(n12516), .B1(
        i_data_bus[748]), .B2(n12518), .ZN(n9907) );
  AOI22D1BWP30P140LVT U10429 ( .A1(i_data_bus[812]), .A2(n12517), .B1(
        i_data_bus[652]), .B2(n12520), .ZN(n9906) );
  AOI22D1BWP30P140LVT U10430 ( .A1(i_data_bus[684]), .A2(n12515), .B1(
        i_data_bus[876]), .B2(n12513), .ZN(n9905) );
  ND4D1BWP30P140LVT U10431 ( .A1(n9908), .A2(n9907), .A3(n9906), .A4(n9905), 
        .ZN(n9909) );
  OR4D1BWP30P140LVT U10432 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), 
        .Z(o_data_bus[140]) );
  AOI22D1BWP30P140LVT U10433 ( .A1(i_data_bus[397]), .A2(n12506), .B1(
        i_data_bus[461]), .B2(n12507), .ZN(n9916) );
  AOI22D1BWP30P140LVT U10434 ( .A1(i_data_bus[941]), .A2(n12492), .B1(
        i_data_bus[141]), .B2(n12502), .ZN(n9915) );
  AOI22D1BWP30P140LVT U10435 ( .A1(i_data_bus[525]), .A2(n12477), .B1(
        i_data_bus[557]), .B2(n12479), .ZN(n9914) );
  AOI22D1BWP30P140LVT U10436 ( .A1(i_data_bus[973]), .A2(n12482), .B1(
        i_data_bus[429]), .B2(n12481), .ZN(n9913) );
  ND4D1BWP30P140LVT U10437 ( .A1(n9916), .A2(n9915), .A3(n9914), .A4(n9913), 
        .ZN(n9932) );
  AOI22D1BWP30P140LVT U10438 ( .A1(i_data_bus[493]), .A2(n12494), .B1(
        i_data_bus[333]), .B2(n12508), .ZN(n9920) );
  AOI22D1BWP30P140LVT U10439 ( .A1(i_data_bus[621]), .A2(n12504), .B1(
        i_data_bus[109]), .B2(n12489), .ZN(n9919) );
  AOI22D1BWP30P140LVT U10440 ( .A1(i_data_bus[301]), .A2(n12505), .B1(
        i_data_bus[173]), .B2(n12501), .ZN(n9918) );
  AOI22D1BWP30P140LVT U10441 ( .A1(i_data_bus[589]), .A2(n12480), .B1(
        i_data_bus[269]), .B2(n12503), .ZN(n9917) );
  ND4D1BWP30P140LVT U10442 ( .A1(n9920), .A2(n9919), .A3(n9918), .A4(n9917), 
        .ZN(n9931) );
  AOI22D1BWP30P140LVT U10443 ( .A1(i_data_bus[45]), .A2(n12483), .B1(
        i_data_bus[1005]), .B2(n12496), .ZN(n9924) );
  AOI22D1BWP30P140LVT U10444 ( .A1(i_data_bus[13]), .A2(n12490), .B1(
        i_data_bus[205]), .B2(n12495), .ZN(n9923) );
  AOI22D1BWP30P140LVT U10445 ( .A1(i_data_bus[909]), .A2(n12484), .B1(
        i_data_bus[365]), .B2(n12491), .ZN(n9922) );
  AOI22D1BWP30P140LVT U10446 ( .A1(i_data_bus[77]), .A2(n12478), .B1(
        i_data_bus[237]), .B2(n12493), .ZN(n9921) );
  ND4D1BWP30P140LVT U10447 ( .A1(n9924), .A2(n9923), .A3(n9922), .A4(n9921), 
        .ZN(n9930) );
  AOI22D1BWP30P140LVT U10448 ( .A1(i_data_bus[749]), .A2(n12518), .B1(
        i_data_bus[845]), .B2(n12514), .ZN(n9928) );
  AOI22D1BWP30P140LVT U10449 ( .A1(i_data_bus[813]), .A2(n12517), .B1(
        i_data_bus[717]), .B2(n12519), .ZN(n9927) );
  AOI22D1BWP30P140LVT U10450 ( .A1(i_data_bus[685]), .A2(n12515), .B1(
        i_data_bus[653]), .B2(n12520), .ZN(n9926) );
  AOI22D1BWP30P140LVT U10451 ( .A1(i_data_bus[877]), .A2(n12513), .B1(
        i_data_bus[781]), .B2(n12516), .ZN(n9925) );
  ND4D1BWP30P140LVT U10452 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), 
        .ZN(n9929) );
  OR4D1BWP30P140LVT U10453 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), 
        .Z(o_data_bus[141]) );
  AOI22D1BWP30P140LVT U10454 ( .A1(i_data_bus[942]), .A2(n12492), .B1(
        i_data_bus[430]), .B2(n12481), .ZN(n9936) );
  AOI22D1BWP30P140LVT U10455 ( .A1(i_data_bus[270]), .A2(n12503), .B1(
        i_data_bus[142]), .B2(n12502), .ZN(n9935) );
  AOI22D1BWP30P140LVT U10456 ( .A1(i_data_bus[334]), .A2(n12508), .B1(
        i_data_bus[398]), .B2(n12506), .ZN(n9934) );
  AOI22D1BWP30P140LVT U10457 ( .A1(i_data_bus[622]), .A2(n12504), .B1(
        i_data_bus[302]), .B2(n12505), .ZN(n9933) );
  ND4D1BWP30P140LVT U10458 ( .A1(n9936), .A2(n9935), .A3(n9934), .A4(n9933), 
        .ZN(n9952) );
  AOI22D1BWP30P140LVT U10459 ( .A1(i_data_bus[558]), .A2(n12479), .B1(
        i_data_bus[174]), .B2(n12501), .ZN(n9940) );
  AOI22D1BWP30P140LVT U10460 ( .A1(i_data_bus[78]), .A2(n12478), .B1(
        i_data_bus[462]), .B2(n12507), .ZN(n9939) );
  AOI22D1BWP30P140LVT U10461 ( .A1(i_data_bus[590]), .A2(n12480), .B1(
        i_data_bus[494]), .B2(n12494), .ZN(n9938) );
  AOI22D1BWP30P140LVT U10462 ( .A1(i_data_bus[366]), .A2(n12491), .B1(
        i_data_bus[238]), .B2(n12493), .ZN(n9937) );
  ND4D1BWP30P140LVT U10463 ( .A1(n9940), .A2(n9939), .A3(n9938), .A4(n9937), 
        .ZN(n9951) );
  AOI22D1BWP30P140LVT U10464 ( .A1(i_data_bus[1006]), .A2(n12496), .B1(
        i_data_bus[526]), .B2(n12477), .ZN(n9944) );
  AOI22D1BWP30P140LVT U10465 ( .A1(i_data_bus[14]), .A2(n12490), .B1(
        i_data_bus[974]), .B2(n12482), .ZN(n9943) );
  AOI22D1BWP30P140LVT U10466 ( .A1(i_data_bus[910]), .A2(n12484), .B1(
        i_data_bus[46]), .B2(n12483), .ZN(n9942) );
  AOI22D1BWP30P140LVT U10467 ( .A1(i_data_bus[110]), .A2(n12489), .B1(
        i_data_bus[206]), .B2(n12495), .ZN(n9941) );
  ND4D1BWP30P140LVT U10468 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), 
        .ZN(n9950) );
  AOI22D1BWP30P140LVT U10469 ( .A1(i_data_bus[814]), .A2(n12517), .B1(
        i_data_bus[878]), .B2(n12513), .ZN(n9948) );
  AOI22D1BWP30P140LVT U10470 ( .A1(i_data_bus[750]), .A2(n12518), .B1(
        i_data_bus[718]), .B2(n12519), .ZN(n9947) );
  AOI22D1BWP30P140LVT U10471 ( .A1(i_data_bus[686]), .A2(n12515), .B1(
        i_data_bus[654]), .B2(n12520), .ZN(n9946) );
  AOI22D1BWP30P140LVT U10472 ( .A1(i_data_bus[846]), .A2(n12514), .B1(
        i_data_bus[782]), .B2(n12516), .ZN(n9945) );
  ND4D1BWP30P140LVT U10473 ( .A1(n9948), .A2(n9947), .A3(n9946), .A4(n9945), 
        .ZN(n9949) );
  OR4D1BWP30P140LVT U10474 ( .A1(n9952), .A2(n9951), .A3(n9950), .A4(n9949), 
        .Z(o_data_bus[142]) );
  AOI22D1BWP30P140LVT U10475 ( .A1(i_data_bus[79]), .A2(n12478), .B1(
        i_data_bus[911]), .B2(n12484), .ZN(n9956) );
  AOI22D1BWP30P140LVT U10476 ( .A1(i_data_bus[975]), .A2(n12482), .B1(
        i_data_bus[591]), .B2(n12480), .ZN(n9955) );
  AOI22D1BWP30P140LVT U10477 ( .A1(i_data_bus[559]), .A2(n12479), .B1(
        i_data_bus[495]), .B2(n12494), .ZN(n9954) );
  AOI22D1BWP30P140LVT U10478 ( .A1(i_data_bus[1007]), .A2(n12496), .B1(
        i_data_bus[207]), .B2(n12495), .ZN(n9953) );
  ND4D1BWP30P140LVT U10479 ( .A1(n9956), .A2(n9955), .A3(n9954), .A4(n9953), 
        .ZN(n9972) );
  AOI22D1BWP30P140LVT U10480 ( .A1(i_data_bus[399]), .A2(n12506), .B1(
        i_data_bus[367]), .B2(n12491), .ZN(n9960) );
  AOI22D1BWP30P140LVT U10481 ( .A1(i_data_bus[47]), .A2(n12483), .B1(
        i_data_bus[15]), .B2(n12490), .ZN(n9959) );
  AOI22D1BWP30P140LVT U10482 ( .A1(i_data_bus[111]), .A2(n12489), .B1(
        i_data_bus[143]), .B2(n12502), .ZN(n9958) );
  AOI22D1BWP30P140LVT U10483 ( .A1(i_data_bus[943]), .A2(n12492), .B1(
        i_data_bus[271]), .B2(n12503), .ZN(n9957) );
  ND4D1BWP30P140LVT U10484 ( .A1(n9960), .A2(n9959), .A3(n9958), .A4(n9957), 
        .ZN(n9971) );
  AOI22D1BWP30P140LVT U10485 ( .A1(i_data_bus[623]), .A2(n12504), .B1(
        i_data_bus[463]), .B2(n12507), .ZN(n9964) );
  AOI22D1BWP30P140LVT U10486 ( .A1(i_data_bus[239]), .A2(n12493), .B1(
        i_data_bus[335]), .B2(n12508), .ZN(n9963) );
  AOI22D1BWP30P140LVT U10487 ( .A1(i_data_bus[527]), .A2(n12477), .B1(
        i_data_bus[175]), .B2(n12501), .ZN(n9962) );
  AOI22D1BWP30P140LVT U10488 ( .A1(i_data_bus[431]), .A2(n12481), .B1(
        i_data_bus[303]), .B2(n12505), .ZN(n9961) );
  ND4D1BWP30P140LVT U10489 ( .A1(n9964), .A2(n9963), .A3(n9962), .A4(n9961), 
        .ZN(n9970) );
  AOI22D1BWP30P140LVT U10490 ( .A1(i_data_bus[847]), .A2(n12514), .B1(
        i_data_bus[655]), .B2(n12520), .ZN(n9968) );
  AOI22D1BWP30P140LVT U10491 ( .A1(i_data_bus[719]), .A2(n12519), .B1(
        i_data_bus[879]), .B2(n12513), .ZN(n9967) );
  AOI22D1BWP30P140LVT U10492 ( .A1(i_data_bus[751]), .A2(n12518), .B1(
        i_data_bus[815]), .B2(n12517), .ZN(n9966) );
  AOI22D1BWP30P140LVT U10493 ( .A1(i_data_bus[783]), .A2(n12516), .B1(
        i_data_bus[687]), .B2(n12515), .ZN(n9965) );
  ND4D1BWP30P140LVT U10494 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), 
        .ZN(n9969) );
  OR4D1BWP30P140LVT U10495 ( .A1(n9972), .A2(n9971), .A3(n9970), .A4(n9969), 
        .Z(o_data_bus[143]) );
  AOI22D1BWP30P140LVT U10496 ( .A1(i_data_bus[48]), .A2(n12483), .B1(
        i_data_bus[240]), .B2(n12493), .ZN(n9976) );
  AOI22D1BWP30P140LVT U10497 ( .A1(i_data_bus[592]), .A2(n12480), .B1(
        i_data_bus[304]), .B2(n12505), .ZN(n9975) );
  AOI22D1BWP30P140LVT U10498 ( .A1(i_data_bus[528]), .A2(n12477), .B1(
        i_data_bus[112]), .B2(n12489), .ZN(n9974) );
  AOI22D1BWP30P140LVT U10499 ( .A1(i_data_bus[912]), .A2(n12484), .B1(
        i_data_bus[208]), .B2(n12495), .ZN(n9973) );
  ND4D1BWP30P140LVT U10500 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), 
        .ZN(n9992) );
  AOI22D1BWP30P140LVT U10501 ( .A1(i_data_bus[80]), .A2(n12478), .B1(
        i_data_bus[624]), .B2(n12504), .ZN(n9980) );
  AOI22D1BWP30P140LVT U10502 ( .A1(i_data_bus[976]), .A2(n12482), .B1(
        i_data_bus[464]), .B2(n12507), .ZN(n9979) );
  AOI22D1BWP30P140LVT U10503 ( .A1(i_data_bus[944]), .A2(n12492), .B1(
        i_data_bus[496]), .B2(n12494), .ZN(n9978) );
  AOI22D1BWP30P140LVT U10504 ( .A1(i_data_bus[1008]), .A2(n12496), .B1(
        i_data_bus[432]), .B2(n12481), .ZN(n9977) );
  ND4D1BWP30P140LVT U10505 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), 
        .ZN(n9991) );
  AOI22D1BWP30P140LVT U10506 ( .A1(i_data_bus[560]), .A2(n12479), .B1(
        i_data_bus[272]), .B2(n12503), .ZN(n9984) );
  AOI22D1BWP30P140LVT U10507 ( .A1(i_data_bus[336]), .A2(n12508), .B1(
        i_data_bus[400]), .B2(n12506), .ZN(n9983) );
  AOI22D1BWP30P140LVT U10508 ( .A1(i_data_bus[144]), .A2(n12502), .B1(
        i_data_bus[176]), .B2(n12501), .ZN(n9982) );
  AOI22D1BWP30P140LVT U10509 ( .A1(i_data_bus[16]), .A2(n12490), .B1(
        i_data_bus[368]), .B2(n12491), .ZN(n9981) );
  ND4D1BWP30P140LVT U10510 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), 
        .ZN(n9990) );
  AOI22D1BWP30P140LVT U10511 ( .A1(i_data_bus[784]), .A2(n12516), .B1(
        i_data_bus[816]), .B2(n12517), .ZN(n9988) );
  AOI22D1BWP30P140LVT U10512 ( .A1(i_data_bus[720]), .A2(n12519), .B1(
        i_data_bus[848]), .B2(n12514), .ZN(n9987) );
  AOI22D1BWP30P140LVT U10513 ( .A1(i_data_bus[880]), .A2(n12513), .B1(
        i_data_bus[752]), .B2(n12518), .ZN(n9986) );
  AOI22D1BWP30P140LVT U10514 ( .A1(i_data_bus[656]), .A2(n12520), .B1(
        i_data_bus[688]), .B2(n12515), .ZN(n9985) );
  ND4D1BWP30P140LVT U10515 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), 
        .ZN(n9989) );
  OR4D1BWP30P140LVT U10516 ( .A1(n9992), .A2(n9991), .A3(n9990), .A4(n9989), 
        .Z(o_data_bus[144]) );
  AOI22D1BWP30P140LVT U10517 ( .A1(i_data_bus[465]), .A2(n12507), .B1(
        i_data_bus[369]), .B2(n12491), .ZN(n9996) );
  AOI22D1BWP30P140LVT U10518 ( .A1(i_data_bus[945]), .A2(n12492), .B1(
        i_data_bus[337]), .B2(n12508), .ZN(n9995) );
  AOI22D1BWP30P140LVT U10519 ( .A1(i_data_bus[241]), .A2(n12493), .B1(
        i_data_bus[273]), .B2(n12503), .ZN(n9994) );
  AOI22D1BWP30P140LVT U10520 ( .A1(i_data_bus[1009]), .A2(n12496), .B1(
        i_data_bus[401]), .B2(n12506), .ZN(n9993) );
  ND4D1BWP30P140LVT U10521 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), 
        .ZN(n10012) );
  AOI22D1BWP30P140LVT U10522 ( .A1(i_data_bus[17]), .A2(n12490), .B1(
        i_data_bus[529]), .B2(n12477), .ZN(n10000) );
  AOI22D1BWP30P140LVT U10523 ( .A1(i_data_bus[433]), .A2(n12481), .B1(
        i_data_bus[177]), .B2(n12501), .ZN(n9999) );
  AOI22D1BWP30P140LVT U10524 ( .A1(i_data_bus[593]), .A2(n12480), .B1(
        i_data_bus[305]), .B2(n12505), .ZN(n9998) );
  AOI22D1BWP30P140LVT U10525 ( .A1(i_data_bus[113]), .A2(n12489), .B1(
        i_data_bus[561]), .B2(n12479), .ZN(n9997) );
  ND4D1BWP30P140LVT U10526 ( .A1(n10000), .A2(n9999), .A3(n9998), .A4(n9997), 
        .ZN(n10011) );
  AOI22D1BWP30P140LVT U10527 ( .A1(i_data_bus[145]), .A2(n12502), .B1(
        i_data_bus[497]), .B2(n12494), .ZN(n10004) );
  AOI22D1BWP30P140LVT U10528 ( .A1(i_data_bus[625]), .A2(n12504), .B1(
        i_data_bus[209]), .B2(n12495), .ZN(n10003) );
  AOI22D1BWP30P140LVT U10529 ( .A1(i_data_bus[49]), .A2(n12483), .B1(
        i_data_bus[81]), .B2(n12478), .ZN(n10002) );
  AOI22D1BWP30P140LVT U10530 ( .A1(i_data_bus[913]), .A2(n12484), .B1(
        i_data_bus[977]), .B2(n12482), .ZN(n10001) );
  ND4D1BWP30P140LVT U10531 ( .A1(n10004), .A2(n10003), .A3(n10002), .A4(n10001), .ZN(n10010) );
  AOI22D1BWP30P140LVT U10532 ( .A1(i_data_bus[785]), .A2(n12516), .B1(
        i_data_bus[817]), .B2(n12517), .ZN(n10008) );
  AOI22D1BWP30P140LVT U10533 ( .A1(i_data_bus[881]), .A2(n12513), .B1(
        i_data_bus[753]), .B2(n12518), .ZN(n10007) );
  AOI22D1BWP30P140LVT U10534 ( .A1(i_data_bus[689]), .A2(n12515), .B1(
        i_data_bus[721]), .B2(n12519), .ZN(n10006) );
  AOI22D1BWP30P140LVT U10535 ( .A1(i_data_bus[849]), .A2(n12514), .B1(
        i_data_bus[657]), .B2(n12520), .ZN(n10005) );
  ND4D1BWP30P140LVT U10536 ( .A1(n10008), .A2(n10007), .A3(n10006), .A4(n10005), .ZN(n10009) );
  OR4D1BWP30P140LVT U10537 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .Z(o_data_bus[145]) );
  AOI22D1BWP30P140LVT U10538 ( .A1(i_data_bus[914]), .A2(n12484), .B1(
        i_data_bus[434]), .B2(n12481), .ZN(n10016) );
  AOI22D1BWP30P140LVT U10539 ( .A1(i_data_bus[562]), .A2(n12479), .B1(
        i_data_bus[338]), .B2(n12508), .ZN(n10015) );
  AOI22D1BWP30P140LVT U10540 ( .A1(i_data_bus[978]), .A2(n12482), .B1(
        i_data_bus[306]), .B2(n12505), .ZN(n10014) );
  AOI22D1BWP30P140LVT U10541 ( .A1(i_data_bus[50]), .A2(n12483), .B1(
        i_data_bus[146]), .B2(n12502), .ZN(n10013) );
  ND4D1BWP30P140LVT U10542 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(n10032) );
  AOI22D1BWP30P140LVT U10543 ( .A1(i_data_bus[18]), .A2(n12490), .B1(
        i_data_bus[178]), .B2(n12501), .ZN(n10020) );
  AOI22D1BWP30P140LVT U10544 ( .A1(i_data_bus[594]), .A2(n12480), .B1(
        i_data_bus[210]), .B2(n12495), .ZN(n10019) );
  AOI22D1BWP30P140LVT U10545 ( .A1(i_data_bus[626]), .A2(n12504), .B1(
        i_data_bus[370]), .B2(n12491), .ZN(n10018) );
  AOI22D1BWP30P140LVT U10546 ( .A1(i_data_bus[1010]), .A2(n12496), .B1(
        i_data_bus[82]), .B2(n12478), .ZN(n10017) );
  ND4D1BWP30P140LVT U10547 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(n10031) );
  AOI22D1BWP30P140LVT U10548 ( .A1(i_data_bus[114]), .A2(n12489), .B1(
        i_data_bus[402]), .B2(n12506), .ZN(n10024) );
  AOI22D1BWP30P140LVT U10549 ( .A1(i_data_bus[242]), .A2(n12493), .B1(
        i_data_bus[274]), .B2(n12503), .ZN(n10023) );
  AOI22D1BWP30P140LVT U10550 ( .A1(i_data_bus[946]), .A2(n12492), .B1(
        i_data_bus[498]), .B2(n12494), .ZN(n10022) );
  AOI22D1BWP30P140LVT U10551 ( .A1(i_data_bus[530]), .A2(n12477), .B1(
        i_data_bus[466]), .B2(n12507), .ZN(n10021) );
  ND4D1BWP30P140LVT U10552 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(n10030) );
  AOI22D1BWP30P140LVT U10553 ( .A1(i_data_bus[658]), .A2(n12520), .B1(
        i_data_bus[754]), .B2(n12518), .ZN(n10028) );
  AOI22D1BWP30P140LVT U10554 ( .A1(i_data_bus[882]), .A2(n12513), .B1(
        i_data_bus[850]), .B2(n12514), .ZN(n10027) );
  AOI22D1BWP30P140LVT U10555 ( .A1(i_data_bus[690]), .A2(n12515), .B1(
        i_data_bus[786]), .B2(n12516), .ZN(n10026) );
  AOI22D1BWP30P140LVT U10556 ( .A1(i_data_bus[722]), .A2(n12519), .B1(
        i_data_bus[818]), .B2(n12517), .ZN(n10025) );
  ND4D1BWP30P140LVT U10557 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(n10029) );
  OR4D1BWP30P140LVT U10558 ( .A1(n10032), .A2(n10031), .A3(n10030), .A4(n10029), .Z(o_data_bus[146]) );
  AOI22D1BWP30P140LVT U10559 ( .A1(i_data_bus[339]), .A2(n12508), .B1(
        i_data_bus[275]), .B2(n12503), .ZN(n10036) );
  AOI22D1BWP30P140LVT U10560 ( .A1(i_data_bus[531]), .A2(n12477), .B1(
        i_data_bus[19]), .B2(n12490), .ZN(n10035) );
  AOI22D1BWP30P140LVT U10561 ( .A1(i_data_bus[947]), .A2(n12492), .B1(
        i_data_bus[499]), .B2(n12494), .ZN(n10034) );
  AOI22D1BWP30P140LVT U10562 ( .A1(i_data_bus[563]), .A2(n12479), .B1(
        i_data_bus[371]), .B2(n12491), .ZN(n10033) );
  ND4D1BWP30P140LVT U10563 ( .A1(n10036), .A2(n10035), .A3(n10034), .A4(n10033), .ZN(n10052) );
  AOI22D1BWP30P140LVT U10564 ( .A1(i_data_bus[979]), .A2(n12482), .B1(
        i_data_bus[627]), .B2(n12504), .ZN(n10040) );
  AOI22D1BWP30P140LVT U10565 ( .A1(i_data_bus[211]), .A2(n12495), .B1(
        i_data_bus[147]), .B2(n12502), .ZN(n10039) );
  AOI22D1BWP30P140LVT U10566 ( .A1(i_data_bus[595]), .A2(n12480), .B1(
        i_data_bus[179]), .B2(n12501), .ZN(n10038) );
  AOI22D1BWP30P140LVT U10567 ( .A1(i_data_bus[51]), .A2(n12483), .B1(
        i_data_bus[243]), .B2(n12493), .ZN(n10037) );
  ND4D1BWP30P140LVT U10568 ( .A1(n10040), .A2(n10039), .A3(n10038), .A4(n10037), .ZN(n10051) );
  AOI22D1BWP30P140LVT U10569 ( .A1(i_data_bus[915]), .A2(n12484), .B1(
        i_data_bus[403]), .B2(n12506), .ZN(n10044) );
  AOI22D1BWP30P140LVT U10570 ( .A1(i_data_bus[83]), .A2(n12478), .B1(
        i_data_bus[435]), .B2(n12481), .ZN(n10043) );
  AOI22D1BWP30P140LVT U10571 ( .A1(i_data_bus[1011]), .A2(n12496), .B1(
        i_data_bus[307]), .B2(n12505), .ZN(n10042) );
  AOI22D1BWP30P140LVT U10572 ( .A1(i_data_bus[115]), .A2(n12489), .B1(
        i_data_bus[467]), .B2(n12507), .ZN(n10041) );
  ND4D1BWP30P140LVT U10573 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(n10050) );
  AOI22D1BWP30P140LVT U10574 ( .A1(i_data_bus[755]), .A2(n12518), .B1(
        i_data_bus[691]), .B2(n12515), .ZN(n10048) );
  AOI22D1BWP30P140LVT U10575 ( .A1(i_data_bus[787]), .A2(n12516), .B1(
        i_data_bus[851]), .B2(n12514), .ZN(n10047) );
  AOI22D1BWP30P140LVT U10576 ( .A1(i_data_bus[819]), .A2(n12517), .B1(
        i_data_bus[723]), .B2(n12519), .ZN(n10046) );
  AOI22D1BWP30P140LVT U10577 ( .A1(i_data_bus[659]), .A2(n12520), .B1(
        i_data_bus[883]), .B2(n12513), .ZN(n10045) );
  ND4D1BWP30P140LVT U10578 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(n10049) );
  OR4D1BWP30P140LVT U10579 ( .A1(n10052), .A2(n10051), .A3(n10050), .A4(n10049), .Z(o_data_bus[147]) );
  AOI22D1BWP30P140LVT U10580 ( .A1(i_data_bus[980]), .A2(n12482), .B1(
        i_data_bus[1012]), .B2(n12496), .ZN(n10056) );
  AOI22D1BWP30P140LVT U10581 ( .A1(i_data_bus[244]), .A2(n12493), .B1(
        i_data_bus[180]), .B2(n12501), .ZN(n10055) );
  AOI22D1BWP30P140LVT U10582 ( .A1(i_data_bus[20]), .A2(n12490), .B1(
        i_data_bus[372]), .B2(n12491), .ZN(n10054) );
  AOI22D1BWP30P140LVT U10583 ( .A1(i_data_bus[628]), .A2(n12504), .B1(
        i_data_bus[404]), .B2(n12506), .ZN(n10053) );
  ND4D1BWP30P140LVT U10584 ( .A1(n10056), .A2(n10055), .A3(n10054), .A4(n10053), .ZN(n10072) );
  AOI22D1BWP30P140LVT U10585 ( .A1(i_data_bus[52]), .A2(n12483), .B1(
        i_data_bus[500]), .B2(n12494), .ZN(n10060) );
  AOI22D1BWP30P140LVT U10586 ( .A1(i_data_bus[340]), .A2(n12508), .B1(
        i_data_bus[276]), .B2(n12503), .ZN(n10059) );
  AOI22D1BWP30P140LVT U10587 ( .A1(i_data_bus[948]), .A2(n12492), .B1(
        i_data_bus[148]), .B2(n12502), .ZN(n10058) );
  AOI22D1BWP30P140LVT U10588 ( .A1(i_data_bus[596]), .A2(n12480), .B1(
        i_data_bus[436]), .B2(n12481), .ZN(n10057) );
  ND4D1BWP30P140LVT U10589 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(n10071) );
  AOI22D1BWP30P140LVT U10590 ( .A1(i_data_bus[532]), .A2(n12477), .B1(
        i_data_bus[308]), .B2(n12505), .ZN(n10064) );
  AOI22D1BWP30P140LVT U10591 ( .A1(i_data_bus[564]), .A2(n12479), .B1(
        i_data_bus[212]), .B2(n12495), .ZN(n10063) );
  AOI22D1BWP30P140LVT U10592 ( .A1(i_data_bus[84]), .A2(n12478), .B1(
        i_data_bus[116]), .B2(n12489), .ZN(n10062) );
  AOI22D1BWP30P140LVT U10593 ( .A1(i_data_bus[916]), .A2(n12484), .B1(
        i_data_bus[468]), .B2(n12507), .ZN(n10061) );
  ND4D1BWP30P140LVT U10594 ( .A1(n10064), .A2(n10063), .A3(n10062), .A4(n10061), .ZN(n10070) );
  AOI22D1BWP30P140LVT U10595 ( .A1(i_data_bus[884]), .A2(n12513), .B1(
        i_data_bus[692]), .B2(n12515), .ZN(n10068) );
  AOI22D1BWP30P140LVT U10596 ( .A1(i_data_bus[724]), .A2(n12519), .B1(
        i_data_bus[820]), .B2(n12517), .ZN(n10067) );
  AOI22D1BWP30P140LVT U10597 ( .A1(i_data_bus[852]), .A2(n12514), .B1(
        i_data_bus[660]), .B2(n12520), .ZN(n10066) );
  AOI22D1BWP30P140LVT U10598 ( .A1(i_data_bus[788]), .A2(n12516), .B1(
        i_data_bus[756]), .B2(n12518), .ZN(n10065) );
  ND4D1BWP30P140LVT U10599 ( .A1(n10068), .A2(n10067), .A3(n10066), .A4(n10065), .ZN(n10069) );
  OR4D1BWP30P140LVT U10600 ( .A1(n10072), .A2(n10071), .A3(n10070), .A4(n10069), .Z(o_data_bus[148]) );
  AOI22D1BWP30P140LVT U10601 ( .A1(i_data_bus[917]), .A2(n12484), .B1(
        i_data_bus[565]), .B2(n12479), .ZN(n10076) );
  AOI22D1BWP30P140LVT U10602 ( .A1(i_data_bus[1013]), .A2(n12496), .B1(
        i_data_bus[149]), .B2(n12502), .ZN(n10075) );
  AOI22D1BWP30P140LVT U10603 ( .A1(i_data_bus[117]), .A2(n12489), .B1(
        i_data_bus[629]), .B2(n12504), .ZN(n10074) );
  AOI22D1BWP30P140LVT U10604 ( .A1(i_data_bus[277]), .A2(n12503), .B1(
        i_data_bus[373]), .B2(n12491), .ZN(n10073) );
  ND4D1BWP30P140LVT U10605 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(n10092) );
  AOI22D1BWP30P140LVT U10606 ( .A1(i_data_bus[53]), .A2(n12483), .B1(
        i_data_bus[533]), .B2(n12477), .ZN(n10080) );
  AOI22D1BWP30P140LVT U10607 ( .A1(i_data_bus[437]), .A2(n12481), .B1(
        i_data_bus[501]), .B2(n12494), .ZN(n10079) );
  AOI22D1BWP30P140LVT U10608 ( .A1(i_data_bus[341]), .A2(n12508), .B1(
        i_data_bus[309]), .B2(n12505), .ZN(n10078) );
  AOI22D1BWP30P140LVT U10609 ( .A1(i_data_bus[597]), .A2(n12480), .B1(
        i_data_bus[181]), .B2(n12501), .ZN(n10077) );
  ND4D1BWP30P140LVT U10610 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(n10091) );
  AOI22D1BWP30P140LVT U10611 ( .A1(i_data_bus[85]), .A2(n12478), .B1(
        i_data_bus[245]), .B2(n12493), .ZN(n10084) );
  AOI22D1BWP30P140LVT U10612 ( .A1(i_data_bus[21]), .A2(n12490), .B1(
        i_data_bus[469]), .B2(n12507), .ZN(n10083) );
  AOI22D1BWP30P140LVT U10613 ( .A1(i_data_bus[981]), .A2(n12482), .B1(
        i_data_bus[213]), .B2(n12495), .ZN(n10082) );
  AOI22D1BWP30P140LVT U10614 ( .A1(i_data_bus[949]), .A2(n12492), .B1(
        i_data_bus[405]), .B2(n12506), .ZN(n10081) );
  ND4D1BWP30P140LVT U10615 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(n10090) );
  AOI22D1BWP30P140LVT U10616 ( .A1(i_data_bus[853]), .A2(n12514), .B1(
        i_data_bus[693]), .B2(n12515), .ZN(n10088) );
  AOI22D1BWP30P140LVT U10617 ( .A1(i_data_bus[661]), .A2(n12520), .B1(
        i_data_bus[725]), .B2(n12519), .ZN(n10087) );
  AOI22D1BWP30P140LVT U10618 ( .A1(i_data_bus[821]), .A2(n12517), .B1(
        i_data_bus[885]), .B2(n12513), .ZN(n10086) );
  AOI22D1BWP30P140LVT U10619 ( .A1(i_data_bus[757]), .A2(n12518), .B1(
        i_data_bus[789]), .B2(n12516), .ZN(n10085) );
  ND4D1BWP30P140LVT U10620 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(n10089) );
  OR4D1BWP30P140LVT U10621 ( .A1(n10092), .A2(n10091), .A3(n10090), .A4(n10089), .Z(o_data_bus[149]) );
  AOI22D1BWP30P140LVT U10622 ( .A1(i_data_bus[118]), .A2(n12489), .B1(
        i_data_bus[470]), .B2(n12507), .ZN(n10096) );
  AOI22D1BWP30P140LVT U10623 ( .A1(i_data_bus[1014]), .A2(n12496), .B1(
        i_data_bus[982]), .B2(n12482), .ZN(n10095) );
  AOI22D1BWP30P140LVT U10624 ( .A1(i_data_bus[534]), .A2(n12477), .B1(
        i_data_bus[150]), .B2(n12502), .ZN(n10094) );
  AOI22D1BWP30P140LVT U10625 ( .A1(i_data_bus[22]), .A2(n12490), .B1(
        i_data_bus[214]), .B2(n12495), .ZN(n10093) );
  ND4D1BWP30P140LVT U10626 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(n10112) );
  AOI22D1BWP30P140LVT U10627 ( .A1(i_data_bus[54]), .A2(n12483), .B1(
        i_data_bus[502]), .B2(n12494), .ZN(n10100) );
  AOI22D1BWP30P140LVT U10628 ( .A1(i_data_bus[566]), .A2(n12479), .B1(
        i_data_bus[310]), .B2(n12505), .ZN(n10099) );
  AOI22D1BWP30P140LVT U10629 ( .A1(i_data_bus[598]), .A2(n12480), .B1(
        i_data_bus[246]), .B2(n12493), .ZN(n10098) );
  AOI22D1BWP30P140LVT U10630 ( .A1(i_data_bus[438]), .A2(n12481), .B1(
        i_data_bus[278]), .B2(n12503), .ZN(n10097) );
  ND4D1BWP30P140LVT U10631 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(n10111) );
  AOI22D1BWP30P140LVT U10632 ( .A1(i_data_bus[86]), .A2(n12478), .B1(
        i_data_bus[630]), .B2(n12504), .ZN(n10104) );
  AOI22D1BWP30P140LVT U10633 ( .A1(i_data_bus[918]), .A2(n12484), .B1(
        i_data_bus[182]), .B2(n12501), .ZN(n10103) );
  AOI22D1BWP30P140LVT U10634 ( .A1(i_data_bus[406]), .A2(n12506), .B1(
        i_data_bus[342]), .B2(n12508), .ZN(n10102) );
  AOI22D1BWP30P140LVT U10635 ( .A1(i_data_bus[950]), .A2(n12492), .B1(
        i_data_bus[374]), .B2(n12491), .ZN(n10101) );
  ND4D1BWP30P140LVT U10636 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(n10110) );
  AOI22D1BWP30P140LVT U10637 ( .A1(i_data_bus[694]), .A2(n12515), .B1(
        i_data_bus[758]), .B2(n12518), .ZN(n10108) );
  AOI22D1BWP30P140LVT U10638 ( .A1(i_data_bus[822]), .A2(n12517), .B1(
        i_data_bus[886]), .B2(n12513), .ZN(n10107) );
  AOI22D1BWP30P140LVT U10639 ( .A1(i_data_bus[790]), .A2(n12516), .B1(
        i_data_bus[854]), .B2(n12514), .ZN(n10106) );
  AOI22D1BWP30P140LVT U10640 ( .A1(i_data_bus[726]), .A2(n12519), .B1(
        i_data_bus[662]), .B2(n12520), .ZN(n10105) );
  ND4D1BWP30P140LVT U10641 ( .A1(n10108), .A2(n10107), .A3(n10106), .A4(n10105), .ZN(n10109) );
  OR4D1BWP30P140LVT U10642 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .Z(o_data_bus[150]) );
  AOI22D1BWP30P140LVT U10643 ( .A1(i_data_bus[567]), .A2(n12479), .B1(
        i_data_bus[151]), .B2(n12502), .ZN(n10116) );
  AOI22D1BWP30P140LVT U10644 ( .A1(i_data_bus[919]), .A2(n12484), .B1(
        i_data_bus[503]), .B2(n12494), .ZN(n10115) );
  AOI22D1BWP30P140LVT U10645 ( .A1(i_data_bus[87]), .A2(n12478), .B1(
        i_data_bus[535]), .B2(n12477), .ZN(n10114) );
  AOI22D1BWP30P140LVT U10646 ( .A1(i_data_bus[599]), .A2(n12480), .B1(
        i_data_bus[407]), .B2(n12506), .ZN(n10113) );
  ND4D1BWP30P140LVT U10647 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(n10132) );
  AOI22D1BWP30P140LVT U10648 ( .A1(i_data_bus[279]), .A2(n12503), .B1(
        i_data_bus[215]), .B2(n12495), .ZN(n10120) );
  AOI22D1BWP30P140LVT U10649 ( .A1(i_data_bus[951]), .A2(n12492), .B1(
        i_data_bus[183]), .B2(n12501), .ZN(n10119) );
  AOI22D1BWP30P140LVT U10650 ( .A1(i_data_bus[471]), .A2(n12507), .B1(
        i_data_bus[375]), .B2(n12491), .ZN(n10118) );
  AOI22D1BWP30P140LVT U10651 ( .A1(i_data_bus[119]), .A2(n12489), .B1(
        i_data_bus[343]), .B2(n12508), .ZN(n10117) );
  ND4D1BWP30P140LVT U10652 ( .A1(n10120), .A2(n10119), .A3(n10118), .A4(n10117), .ZN(n10131) );
  AOI22D1BWP30P140LVT U10653 ( .A1(i_data_bus[247]), .A2(n12493), .B1(
        i_data_bus[439]), .B2(n12481), .ZN(n10124) );
  AOI22D1BWP30P140LVT U10654 ( .A1(i_data_bus[1015]), .A2(n12496), .B1(
        i_data_bus[311]), .B2(n12505), .ZN(n10123) );
  AOI22D1BWP30P140LVT U10655 ( .A1(i_data_bus[23]), .A2(n12490), .B1(
        i_data_bus[55]), .B2(n12483), .ZN(n10122) );
  AOI22D1BWP30P140LVT U10656 ( .A1(i_data_bus[631]), .A2(n12504), .B1(
        i_data_bus[983]), .B2(n12482), .ZN(n10121) );
  ND4D1BWP30P140LVT U10657 ( .A1(n10124), .A2(n10123), .A3(n10122), .A4(n10121), .ZN(n10130) );
  AOI22D1BWP30P140LVT U10658 ( .A1(i_data_bus[887]), .A2(n12513), .B1(
        i_data_bus[855]), .B2(n12514), .ZN(n10128) );
  AOI22D1BWP30P140LVT U10659 ( .A1(i_data_bus[695]), .A2(n12515), .B1(
        i_data_bus[663]), .B2(n12520), .ZN(n10127) );
  AOI22D1BWP30P140LVT U10660 ( .A1(i_data_bus[759]), .A2(n12518), .B1(
        i_data_bus[823]), .B2(n12517), .ZN(n10126) );
  AOI22D1BWP30P140LVT U10661 ( .A1(i_data_bus[727]), .A2(n12519), .B1(
        i_data_bus[791]), .B2(n12516), .ZN(n10125) );
  ND4D1BWP30P140LVT U10662 ( .A1(n10128), .A2(n10127), .A3(n10126), .A4(n10125), .ZN(n10129) );
  OR4D1BWP30P140LVT U10663 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .Z(o_data_bus[151]) );
  AOI22D1BWP30P140LVT U10664 ( .A1(i_data_bus[24]), .A2(n12490), .B1(
        i_data_bus[344]), .B2(n12508), .ZN(n10136) );
  AOI22D1BWP30P140LVT U10665 ( .A1(i_data_bus[88]), .A2(n12478), .B1(
        i_data_bus[248]), .B2(n12493), .ZN(n10135) );
  AOI22D1BWP30P140LVT U10666 ( .A1(i_data_bus[920]), .A2(n12484), .B1(
        i_data_bus[472]), .B2(n12507), .ZN(n10134) );
  AOI22D1BWP30P140LVT U10667 ( .A1(i_data_bus[280]), .A2(n12503), .B1(
        i_data_bus[504]), .B2(n12494), .ZN(n10133) );
  ND4D1BWP30P140LVT U10668 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(n10152) );
  AOI22D1BWP30P140LVT U10669 ( .A1(i_data_bus[984]), .A2(n12482), .B1(
        i_data_bus[184]), .B2(n12501), .ZN(n10140) );
  AOI22D1BWP30P140LVT U10670 ( .A1(i_data_bus[536]), .A2(n12477), .B1(
        i_data_bus[440]), .B2(n12481), .ZN(n10139) );
  AOI22D1BWP30P140LVT U10671 ( .A1(i_data_bus[568]), .A2(n12479), .B1(
        i_data_bus[376]), .B2(n12491), .ZN(n10138) );
  AOI22D1BWP30P140LVT U10672 ( .A1(i_data_bus[632]), .A2(n12504), .B1(
        i_data_bus[600]), .B2(n12480), .ZN(n10137) );
  ND4D1BWP30P140LVT U10673 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(n10151) );
  AOI22D1BWP30P140LVT U10674 ( .A1(i_data_bus[952]), .A2(n12492), .B1(
        i_data_bus[56]), .B2(n12483), .ZN(n10144) );
  AOI22D1BWP30P140LVT U10675 ( .A1(i_data_bus[120]), .A2(n12489), .B1(
        i_data_bus[152]), .B2(n12502), .ZN(n10143) );
  AOI22D1BWP30P140LVT U10676 ( .A1(i_data_bus[408]), .A2(n12506), .B1(
        i_data_bus[216]), .B2(n12495), .ZN(n10142) );
  AOI22D1BWP30P140LVT U10677 ( .A1(i_data_bus[1016]), .A2(n12496), .B1(
        i_data_bus[312]), .B2(n12505), .ZN(n10141) );
  ND4D1BWP30P140LVT U10678 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(n10150) );
  AOI22D1BWP30P140LVT U10679 ( .A1(i_data_bus[792]), .A2(n12516), .B1(
        i_data_bus[728]), .B2(n12519), .ZN(n10148) );
  AOI22D1BWP30P140LVT U10680 ( .A1(i_data_bus[856]), .A2(n12514), .B1(
        i_data_bus[888]), .B2(n12513), .ZN(n10147) );
  AOI22D1BWP30P140LVT U10681 ( .A1(i_data_bus[696]), .A2(n12515), .B1(
        i_data_bus[760]), .B2(n12518), .ZN(n10146) );
  AOI22D1BWP30P140LVT U10682 ( .A1(i_data_bus[824]), .A2(n12517), .B1(
        i_data_bus[664]), .B2(n12520), .ZN(n10145) );
  ND4D1BWP30P140LVT U10683 ( .A1(n10148), .A2(n10147), .A3(n10146), .A4(n10145), .ZN(n10149) );
  OR4D1BWP30P140LVT U10684 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .Z(o_data_bus[152]) );
  AOI22D1BWP30P140LVT U10685 ( .A1(i_data_bus[985]), .A2(n12482), .B1(
        i_data_bus[409]), .B2(n12506), .ZN(n10156) );
  AOI22D1BWP30P140LVT U10686 ( .A1(i_data_bus[377]), .A2(n12491), .B1(
        i_data_bus[441]), .B2(n12481), .ZN(n10155) );
  AOI22D1BWP30P140LVT U10687 ( .A1(i_data_bus[281]), .A2(n12503), .B1(
        i_data_bus[217]), .B2(n12495), .ZN(n10154) );
  AOI22D1BWP30P140LVT U10688 ( .A1(i_data_bus[1017]), .A2(n12496), .B1(
        i_data_bus[89]), .B2(n12478), .ZN(n10153) );
  ND4D1BWP30P140LVT U10689 ( .A1(n10156), .A2(n10155), .A3(n10154), .A4(n10153), .ZN(n10172) );
  AOI22D1BWP30P140LVT U10690 ( .A1(i_data_bus[601]), .A2(n12480), .B1(
        i_data_bus[313]), .B2(n12505), .ZN(n10160) );
  AOI22D1BWP30P140LVT U10691 ( .A1(i_data_bus[185]), .A2(n12501), .B1(
        i_data_bus[505]), .B2(n12494), .ZN(n10159) );
  AOI22D1BWP30P140LVT U10692 ( .A1(i_data_bus[57]), .A2(n12483), .B1(
        i_data_bus[121]), .B2(n12489), .ZN(n10158) );
  AOI22D1BWP30P140LVT U10693 ( .A1(i_data_bus[537]), .A2(n12477), .B1(
        i_data_bus[473]), .B2(n12507), .ZN(n10157) );
  ND4D1BWP30P140LVT U10694 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(n10171) );
  AOI22D1BWP30P140LVT U10695 ( .A1(i_data_bus[25]), .A2(n12490), .B1(
        i_data_bus[249]), .B2(n12493), .ZN(n10164) );
  AOI22D1BWP30P140LVT U10696 ( .A1(i_data_bus[569]), .A2(n12479), .B1(
        i_data_bus[153]), .B2(n12502), .ZN(n10163) );
  AOI22D1BWP30P140LVT U10697 ( .A1(i_data_bus[633]), .A2(n12504), .B1(
        i_data_bus[953]), .B2(n12492), .ZN(n10162) );
  AOI22D1BWP30P140LVT U10698 ( .A1(i_data_bus[921]), .A2(n12484), .B1(
        i_data_bus[345]), .B2(n12508), .ZN(n10161) );
  ND4D1BWP30P140LVT U10699 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(n10170) );
  AOI22D1BWP30P140LVT U10700 ( .A1(i_data_bus[825]), .A2(n12517), .B1(
        i_data_bus[729]), .B2(n12519), .ZN(n10168) );
  AOI22D1BWP30P140LVT U10701 ( .A1(i_data_bus[761]), .A2(n12518), .B1(
        i_data_bus[889]), .B2(n12513), .ZN(n10167) );
  AOI22D1BWP30P140LVT U10702 ( .A1(i_data_bus[665]), .A2(n12520), .B1(
        i_data_bus[793]), .B2(n12516), .ZN(n10166) );
  AOI22D1BWP30P140LVT U10703 ( .A1(i_data_bus[697]), .A2(n12515), .B1(
        i_data_bus[857]), .B2(n12514), .ZN(n10165) );
  ND4D1BWP30P140LVT U10704 ( .A1(n10168), .A2(n10167), .A3(n10166), .A4(n10165), .ZN(n10169) );
  OR4D1BWP30P140LVT U10705 ( .A1(n10172), .A2(n10171), .A3(n10170), .A4(n10169), .Z(o_data_bus[153]) );
  AOI22D1BWP30P140LVT U10706 ( .A1(i_data_bus[602]), .A2(n12480), .B1(
        i_data_bus[506]), .B2(n12494), .ZN(n10176) );
  AOI22D1BWP30P140LVT U10707 ( .A1(i_data_bus[122]), .A2(n12489), .B1(
        i_data_bus[186]), .B2(n12501), .ZN(n10175) );
  AOI22D1BWP30P140LVT U10708 ( .A1(i_data_bus[90]), .A2(n12478), .B1(
        i_data_bus[218]), .B2(n12495), .ZN(n10174) );
  AOI22D1BWP30P140LVT U10709 ( .A1(i_data_bus[570]), .A2(n12479), .B1(
        i_data_bus[410]), .B2(n12506), .ZN(n10173) );
  ND4D1BWP30P140LVT U10710 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(n10192) );
  AOI22D1BWP30P140LVT U10711 ( .A1(i_data_bus[922]), .A2(n12484), .B1(
        i_data_bus[250]), .B2(n12493), .ZN(n10180) );
  AOI22D1BWP30P140LVT U10712 ( .A1(i_data_bus[954]), .A2(n12492), .B1(
        i_data_bus[634]), .B2(n12504), .ZN(n10179) );
  AOI22D1BWP30P140LVT U10713 ( .A1(i_data_bus[346]), .A2(n12508), .B1(
        i_data_bus[282]), .B2(n12503), .ZN(n10178) );
  AOI22D1BWP30P140LVT U10714 ( .A1(i_data_bus[1018]), .A2(n12496), .B1(
        i_data_bus[58]), .B2(n12483), .ZN(n10177) );
  ND4D1BWP30P140LVT U10715 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(n10191) );
  AOI22D1BWP30P140LVT U10716 ( .A1(i_data_bus[986]), .A2(n12482), .B1(
        i_data_bus[314]), .B2(n12505), .ZN(n10184) );
  AOI22D1BWP30P140LVT U10717 ( .A1(i_data_bus[154]), .A2(n12502), .B1(
        i_data_bus[378]), .B2(n12491), .ZN(n10183) );
  AOI22D1BWP30P140LVT U10718 ( .A1(i_data_bus[538]), .A2(n12477), .B1(
        i_data_bus[442]), .B2(n12481), .ZN(n10182) );
  AOI22D1BWP30P140LVT U10719 ( .A1(i_data_bus[26]), .A2(n12490), .B1(
        i_data_bus[474]), .B2(n12507), .ZN(n10181) );
  ND4D1BWP30P140LVT U10720 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(n10190) );
  AOI22D1BWP30P140LVT U10721 ( .A1(i_data_bus[826]), .A2(n12517), .B1(
        i_data_bus[890]), .B2(n12513), .ZN(n10188) );
  AOI22D1BWP30P140LVT U10722 ( .A1(i_data_bus[794]), .A2(n12516), .B1(
        i_data_bus[666]), .B2(n12520), .ZN(n10187) );
  AOI22D1BWP30P140LVT U10723 ( .A1(i_data_bus[858]), .A2(n12514), .B1(
        i_data_bus[762]), .B2(n12518), .ZN(n10186) );
  AOI22D1BWP30P140LVT U10724 ( .A1(i_data_bus[698]), .A2(n12515), .B1(
        i_data_bus[730]), .B2(n12519), .ZN(n10185) );
  ND4D1BWP30P140LVT U10725 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(n10189) );
  OR4D1BWP30P140LVT U10726 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .Z(o_data_bus[154]) );
  AOI22D1BWP30P140LVT U10727 ( .A1(i_data_bus[539]), .A2(n12477), .B1(
        i_data_bus[475]), .B2(n12507), .ZN(n10196) );
  AOI22D1BWP30P140LVT U10728 ( .A1(i_data_bus[635]), .A2(n12504), .B1(
        i_data_bus[27]), .B2(n12490), .ZN(n10195) );
  AOI22D1BWP30P140LVT U10729 ( .A1(i_data_bus[155]), .A2(n12502), .B1(
        i_data_bus[251]), .B2(n12493), .ZN(n10194) );
  AOI22D1BWP30P140LVT U10730 ( .A1(i_data_bus[379]), .A2(n12491), .B1(
        i_data_bus[347]), .B2(n12508), .ZN(n10193) );
  ND4D1BWP30P140LVT U10731 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(n10212) );
  AOI22D1BWP30P140LVT U10732 ( .A1(i_data_bus[59]), .A2(n12483), .B1(
        i_data_bus[315]), .B2(n12505), .ZN(n10200) );
  AOI22D1BWP30P140LVT U10733 ( .A1(i_data_bus[603]), .A2(n12480), .B1(
        i_data_bus[923]), .B2(n12484), .ZN(n10199) );
  AOI22D1BWP30P140LVT U10734 ( .A1(i_data_bus[571]), .A2(n12479), .B1(
        i_data_bus[283]), .B2(n12503), .ZN(n10198) );
  AOI22D1BWP30P140LVT U10735 ( .A1(i_data_bus[987]), .A2(n12482), .B1(
        i_data_bus[187]), .B2(n12501), .ZN(n10197) );
  ND4D1BWP30P140LVT U10736 ( .A1(n10200), .A2(n10199), .A3(n10198), .A4(n10197), .ZN(n10211) );
  AOI22D1BWP30P140LVT U10737 ( .A1(i_data_bus[123]), .A2(n12489), .B1(
        i_data_bus[1019]), .B2(n12496), .ZN(n10204) );
  AOI22D1BWP30P140LVT U10738 ( .A1(i_data_bus[955]), .A2(n12492), .B1(
        i_data_bus[411]), .B2(n12506), .ZN(n10203) );
  AOI22D1BWP30P140LVT U10739 ( .A1(i_data_bus[91]), .A2(n12478), .B1(
        i_data_bus[443]), .B2(n12481), .ZN(n10202) );
  AOI22D1BWP30P140LVT U10740 ( .A1(i_data_bus[507]), .A2(n12494), .B1(
        i_data_bus[219]), .B2(n12495), .ZN(n10201) );
  ND4D1BWP30P140LVT U10741 ( .A1(n10204), .A2(n10203), .A3(n10202), .A4(n10201), .ZN(n10210) );
  AOI22D1BWP30P140LVT U10742 ( .A1(i_data_bus[763]), .A2(n12518), .B1(
        i_data_bus[699]), .B2(n12515), .ZN(n10208) );
  AOI22D1BWP30P140LVT U10743 ( .A1(i_data_bus[795]), .A2(n12516), .B1(
        i_data_bus[859]), .B2(n12514), .ZN(n10207) );
  AOI22D1BWP30P140LVT U10744 ( .A1(i_data_bus[827]), .A2(n12517), .B1(
        i_data_bus[667]), .B2(n12520), .ZN(n10206) );
  AOI22D1BWP30P140LVT U10745 ( .A1(i_data_bus[731]), .A2(n12519), .B1(
        i_data_bus[891]), .B2(n12513), .ZN(n10205) );
  ND4D1BWP30P140LVT U10746 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(n10209) );
  OR4D1BWP30P140LVT U10747 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .Z(o_data_bus[155]) );
  AOI22D1BWP30P140LVT U10748 ( .A1(i_data_bus[1020]), .A2(n12496), .B1(
        i_data_bus[508]), .B2(n12494), .ZN(n10216) );
  AOI22D1BWP30P140LVT U10749 ( .A1(i_data_bus[92]), .A2(n12478), .B1(
        i_data_bus[412]), .B2(n12506), .ZN(n10215) );
  AOI22D1BWP30P140LVT U10750 ( .A1(i_data_bus[604]), .A2(n12480), .B1(
        i_data_bus[348]), .B2(n12508), .ZN(n10214) );
  AOI22D1BWP30P140LVT U10751 ( .A1(i_data_bus[540]), .A2(n12477), .B1(
        i_data_bus[220]), .B2(n12495), .ZN(n10213) );
  ND4D1BWP30P140LVT U10752 ( .A1(n10216), .A2(n10215), .A3(n10214), .A4(n10213), .ZN(n10232) );
  AOI22D1BWP30P140LVT U10753 ( .A1(i_data_bus[636]), .A2(n12504), .B1(
        i_data_bus[252]), .B2(n12493), .ZN(n10220) );
  AOI22D1BWP30P140LVT U10754 ( .A1(i_data_bus[476]), .A2(n12507), .B1(
        i_data_bus[316]), .B2(n12505), .ZN(n10219) );
  AOI22D1BWP30P140LVT U10755 ( .A1(i_data_bus[956]), .A2(n12492), .B1(
        i_data_bus[284]), .B2(n12503), .ZN(n10218) );
  AOI22D1BWP30P140LVT U10756 ( .A1(i_data_bus[28]), .A2(n12490), .B1(
        i_data_bus[572]), .B2(n12479), .ZN(n10217) );
  ND4D1BWP30P140LVT U10757 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(n10231) );
  AOI22D1BWP30P140LVT U10758 ( .A1(i_data_bus[988]), .A2(n12482), .B1(
        i_data_bus[380]), .B2(n12491), .ZN(n10224) );
  AOI22D1BWP30P140LVT U10759 ( .A1(i_data_bus[60]), .A2(n12483), .B1(
        i_data_bus[156]), .B2(n12502), .ZN(n10223) );
  AOI22D1BWP30P140LVT U10760 ( .A1(i_data_bus[924]), .A2(n12484), .B1(
        i_data_bus[444]), .B2(n12481), .ZN(n10222) );
  AOI22D1BWP30P140LVT U10761 ( .A1(i_data_bus[124]), .A2(n12489), .B1(
        i_data_bus[188]), .B2(n12501), .ZN(n10221) );
  ND4D1BWP30P140LVT U10762 ( .A1(n10224), .A2(n10223), .A3(n10222), .A4(n10221), .ZN(n10230) );
  AOI22D1BWP30P140LVT U10763 ( .A1(i_data_bus[732]), .A2(n12519), .B1(
        i_data_bus[764]), .B2(n12518), .ZN(n10228) );
  AOI22D1BWP30P140LVT U10764 ( .A1(i_data_bus[796]), .A2(n12516), .B1(
        i_data_bus[700]), .B2(n12515), .ZN(n10227) );
  AOI22D1BWP30P140LVT U10765 ( .A1(i_data_bus[828]), .A2(n12517), .B1(
        i_data_bus[860]), .B2(n12514), .ZN(n10226) );
  AOI22D1BWP30P140LVT U10766 ( .A1(i_data_bus[892]), .A2(n12513), .B1(
        i_data_bus[668]), .B2(n12520), .ZN(n10225) );
  ND4D1BWP30P140LVT U10767 ( .A1(n10228), .A2(n10227), .A3(n10226), .A4(n10225), .ZN(n10229) );
  OR4D1BWP30P140LVT U10768 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .Z(o_data_bus[156]) );
  AOI22D1BWP30P140LVT U10769 ( .A1(i_data_bus[637]), .A2(n12504), .B1(
        i_data_bus[541]), .B2(n12477), .ZN(n10236) );
  AOI22D1BWP30P140LVT U10770 ( .A1(i_data_bus[29]), .A2(n12490), .B1(
        i_data_bus[285]), .B2(n12503), .ZN(n10235) );
  AOI22D1BWP30P140LVT U10771 ( .A1(i_data_bus[477]), .A2(n12507), .B1(
        i_data_bus[413]), .B2(n12506), .ZN(n10234) );
  AOI22D1BWP30P140LVT U10772 ( .A1(i_data_bus[957]), .A2(n12492), .B1(
        i_data_bus[93]), .B2(n12478), .ZN(n10233) );
  ND4D1BWP30P140LVT U10773 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(n10252) );
  AOI22D1BWP30P140LVT U10774 ( .A1(i_data_bus[61]), .A2(n12483), .B1(
        i_data_bus[157]), .B2(n12502), .ZN(n10240) );
  AOI22D1BWP30P140LVT U10775 ( .A1(i_data_bus[125]), .A2(n12489), .B1(
        i_data_bus[445]), .B2(n12481), .ZN(n10239) );
  AOI22D1BWP30P140LVT U10776 ( .A1(i_data_bus[1021]), .A2(n12496), .B1(
        i_data_bus[349]), .B2(n12508), .ZN(n10238) );
  AOI22D1BWP30P140LVT U10777 ( .A1(i_data_bus[381]), .A2(n12491), .B1(
        i_data_bus[253]), .B2(n12493), .ZN(n10237) );
  ND4D1BWP30P140LVT U10778 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(n10251) );
  AOI22D1BWP30P140LVT U10779 ( .A1(i_data_bus[925]), .A2(n12484), .B1(
        i_data_bus[189]), .B2(n12501), .ZN(n10244) );
  AOI22D1BWP30P140LVT U10780 ( .A1(i_data_bus[573]), .A2(n12479), .B1(
        i_data_bus[317]), .B2(n12505), .ZN(n10243) );
  AOI22D1BWP30P140LVT U10781 ( .A1(i_data_bus[509]), .A2(n12494), .B1(
        i_data_bus[221]), .B2(n12495), .ZN(n10242) );
  AOI22D1BWP30P140LVT U10782 ( .A1(i_data_bus[989]), .A2(n12482), .B1(
        i_data_bus[605]), .B2(n12480), .ZN(n10241) );
  ND4D1BWP30P140LVT U10783 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(n10250) );
  AOI22D1BWP30P140LVT U10784 ( .A1(i_data_bus[765]), .A2(n12518), .B1(
        i_data_bus[797]), .B2(n12516), .ZN(n10248) );
  AOI22D1BWP30P140LVT U10785 ( .A1(i_data_bus[733]), .A2(n12519), .B1(
        i_data_bus[829]), .B2(n12517), .ZN(n10247) );
  AOI22D1BWP30P140LVT U10786 ( .A1(i_data_bus[861]), .A2(n12514), .B1(
        i_data_bus[893]), .B2(n12513), .ZN(n10246) );
  AOI22D1BWP30P140LVT U10787 ( .A1(i_data_bus[701]), .A2(n12515), .B1(
        i_data_bus[669]), .B2(n12520), .ZN(n10245) );
  ND4D1BWP30P140LVT U10788 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(n10249) );
  OR4D1BWP30P140LVT U10789 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .Z(o_data_bus[157]) );
  AOI22D1BWP30P140LVT U10790 ( .A1(i_data_bus[926]), .A2(n12484), .B1(
        i_data_bus[350]), .B2(n12508), .ZN(n10256) );
  AOI22D1BWP30P140LVT U10791 ( .A1(i_data_bus[318]), .A2(n12505), .B1(
        i_data_bus[158]), .B2(n12502), .ZN(n10255) );
  AOI22D1BWP30P140LVT U10792 ( .A1(i_data_bus[62]), .A2(n12483), .B1(
        i_data_bus[30]), .B2(n12490), .ZN(n10254) );
  AOI22D1BWP30P140LVT U10793 ( .A1(i_data_bus[958]), .A2(n12492), .B1(
        i_data_bus[94]), .B2(n12478), .ZN(n10253) );
  ND4D1BWP30P140LVT U10794 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(n10272) );
  AOI22D1BWP30P140LVT U10795 ( .A1(i_data_bus[1022]), .A2(n12496), .B1(
        i_data_bus[286]), .B2(n12503), .ZN(n10260) );
  AOI22D1BWP30P140LVT U10796 ( .A1(i_data_bus[990]), .A2(n12482), .B1(
        i_data_bus[382]), .B2(n12491), .ZN(n10259) );
  AOI22D1BWP30P140LVT U10797 ( .A1(i_data_bus[606]), .A2(n12480), .B1(
        i_data_bus[478]), .B2(n12507), .ZN(n10258) );
  AOI22D1BWP30P140LVT U10798 ( .A1(i_data_bus[222]), .A2(n12495), .B1(
        i_data_bus[446]), .B2(n12481), .ZN(n10257) );
  ND4D1BWP30P140LVT U10799 ( .A1(n10260), .A2(n10259), .A3(n10258), .A4(n10257), .ZN(n10271) );
  AOI22D1BWP30P140LVT U10800 ( .A1(i_data_bus[574]), .A2(n12479), .B1(
        i_data_bus[510]), .B2(n12494), .ZN(n10264) );
  AOI22D1BWP30P140LVT U10801 ( .A1(i_data_bus[190]), .A2(n12501), .B1(
        i_data_bus[414]), .B2(n12506), .ZN(n10263) );
  AOI22D1BWP30P140LVT U10802 ( .A1(i_data_bus[542]), .A2(n12477), .B1(
        i_data_bus[126]), .B2(n12489), .ZN(n10262) );
  AOI22D1BWP30P140LVT U10803 ( .A1(i_data_bus[638]), .A2(n12504), .B1(
        i_data_bus[254]), .B2(n12493), .ZN(n10261) );
  ND4D1BWP30P140LVT U10804 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(n10270) );
  AOI22D1BWP30P140LVT U10805 ( .A1(i_data_bus[862]), .A2(n12514), .B1(
        i_data_bus[702]), .B2(n12515), .ZN(n10268) );
  AOI22D1BWP30P140LVT U10806 ( .A1(i_data_bus[670]), .A2(n12520), .B1(
        i_data_bus[734]), .B2(n12519), .ZN(n10267) );
  AOI22D1BWP30P140LVT U10807 ( .A1(i_data_bus[830]), .A2(n12517), .B1(
        i_data_bus[894]), .B2(n12513), .ZN(n10266) );
  AOI22D1BWP30P140LVT U10808 ( .A1(i_data_bus[798]), .A2(n12516), .B1(
        i_data_bus[766]), .B2(n12518), .ZN(n10265) );
  ND4D1BWP30P140LVT U10809 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(n10269) );
  OR4D1BWP30P140LVT U10810 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .Z(o_data_bus[158]) );
  AOI22D1BWP30P140LVT U10811 ( .A1(i_data_bus[159]), .A2(n12502), .B1(
        i_data_bus[479]), .B2(n12507), .ZN(n10276) );
  AOI22D1BWP30P140LVT U10812 ( .A1(i_data_bus[95]), .A2(n12478), .B1(
        i_data_bus[543]), .B2(n12477), .ZN(n10275) );
  AOI22D1BWP30P140LVT U10813 ( .A1(i_data_bus[319]), .A2(n12505), .B1(
        i_data_bus[255]), .B2(n12493), .ZN(n10274) );
  AOI22D1BWP30P140LVT U10814 ( .A1(i_data_bus[287]), .A2(n12503), .B1(
        i_data_bus[191]), .B2(n12501), .ZN(n10273) );
  ND4D1BWP30P140LVT U10815 ( .A1(n10276), .A2(n10275), .A3(n10274), .A4(n10273), .ZN(n10292) );
  AOI22D1BWP30P140LVT U10816 ( .A1(i_data_bus[927]), .A2(n12484), .B1(
        i_data_bus[959]), .B2(n12492), .ZN(n10280) );
  AOI22D1BWP30P140LVT U10817 ( .A1(i_data_bus[415]), .A2(n12506), .B1(
        i_data_bus[383]), .B2(n12491), .ZN(n10279) );
  AOI22D1BWP30P140LVT U10818 ( .A1(i_data_bus[1023]), .A2(n12496), .B1(
        i_data_bus[447]), .B2(n12481), .ZN(n10278) );
  AOI22D1BWP30P140LVT U10819 ( .A1(i_data_bus[575]), .A2(n12479), .B1(
        i_data_bus[639]), .B2(n12504), .ZN(n10277) );
  ND4D1BWP30P140LVT U10820 ( .A1(n10280), .A2(n10279), .A3(n10278), .A4(n10277), .ZN(n10291) );
  AOI22D1BWP30P140LVT U10821 ( .A1(i_data_bus[31]), .A2(n12490), .B1(
        i_data_bus[127]), .B2(n12489), .ZN(n10284) );
  AOI22D1BWP30P140LVT U10822 ( .A1(i_data_bus[991]), .A2(n12482), .B1(
        i_data_bus[351]), .B2(n12508), .ZN(n10283) );
  AOI22D1BWP30P140LVT U10823 ( .A1(i_data_bus[63]), .A2(n12483), .B1(
        i_data_bus[223]), .B2(n12495), .ZN(n10282) );
  AOI22D1BWP30P140LVT U10824 ( .A1(i_data_bus[607]), .A2(n12480), .B1(
        i_data_bus[511]), .B2(n12494), .ZN(n10281) );
  ND4D1BWP30P140LVT U10825 ( .A1(n10284), .A2(n10283), .A3(n10282), .A4(n10281), .ZN(n10290) );
  AOI22D1BWP30P140LVT U10826 ( .A1(i_data_bus[767]), .A2(n12518), .B1(
        i_data_bus[831]), .B2(n12517), .ZN(n10288) );
  AOI22D1BWP30P140LVT U10827 ( .A1(i_data_bus[863]), .A2(n12514), .B1(
        i_data_bus[703]), .B2(n12515), .ZN(n10287) );
  AOI22D1BWP30P140LVT U10828 ( .A1(i_data_bus[799]), .A2(n12516), .B1(
        i_data_bus[671]), .B2(n12520), .ZN(n10286) );
  AOI22D1BWP30P140LVT U10829 ( .A1(i_data_bus[735]), .A2(n12519), .B1(
        i_data_bus[895]), .B2(n12513), .ZN(n10285) );
  ND4D1BWP30P140LVT U10830 ( .A1(n10288), .A2(n10287), .A3(n10286), .A4(n10285), .ZN(n10289) );
  OR4D1BWP30P140LVT U10831 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .Z(o_data_bus[159]) );
  NR3D0P7BWP30P140LVT U10832 ( .A1(n11717), .A2(n10293), .A3(n10296), .ZN(
        n10955) );
  NR3D0P7BWP30P140LVT U10833 ( .A1(n11715), .A2(n10294), .A3(n10296), .ZN(
        n10953) );
  AOI22D1BWP30P140LVT U10834 ( .A1(i_data_bus[992]), .A2(n10955), .B1(
        i_data_bus[960]), .B2(n10953), .ZN(n10301) );
  NR3D0P7BWP30P140LVT U10835 ( .A1(n11740), .A2(n10295), .A3(n10296), .ZN(
        n10954) );
  NR3D0P7BWP30P140LVT U10836 ( .A1(n11735), .A2(n10297), .A3(n10296), .ZN(
        n10952) );
  AOI22D1BWP30P140LVT U10837 ( .A1(i_data_bus[928]), .A2(n10954), .B1(
        i_data_bus[896]), .B2(n10952), .ZN(n10300) );
  INR3D0BWP30P140LVT U10838 ( .A1(i_cmd[94]), .B1(n11731), .B2(n10309), .ZN(
        n10978) );
  INR3D0BWP30P140LVT U10839 ( .A1(i_cmd[174]), .B1(n11756), .B2(n10308), .ZN(
        n10977) );
  AOI22D1BWP30P140LVT U10840 ( .A1(i_data_bus[352]), .A2(n10978), .B1(
        i_data_bus[672]), .B2(n10977), .ZN(n10299) );
  INR3D0BWP30P140LVT U10841 ( .A1(i_cmd[158]), .B1(n11697), .B2(n10316), .ZN(
        n10971) );
  INR3D0BWP30P140LVT U10842 ( .A1(i_cmd[206]), .B1(n11751), .B2(n10319), .ZN(
        n10970) );
  AOI22D1BWP30P140LVT U10843 ( .A1(i_data_bus[608]), .A2(n10971), .B1(
        i_data_bus[800]), .B2(n10970), .ZN(n10298) );
  ND4D1BWP30P140LVT U10844 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n10298), .ZN(n10331) );
  INR3D0BWP30P140LVT U10845 ( .A1(i_cmd[150]), .B1(n11733), .B2(n10316), .ZN(
        n10981) );
  INVD1BWP30P140LVT U10846 ( .I(i_cmd[70]), .ZN(n10302) );
  NR3D0P7BWP30P140LVT U10847 ( .A1(n11728), .A2(n10302), .A3(n10309), .ZN(
        n10968) );
  AOI22D1BWP30P140LVT U10848 ( .A1(i_data_bus[576]), .A2(n10981), .B1(
        i_data_bus[256]), .B2(n10968), .ZN(n10307) );
  INR3D0BWP30P140LVT U10849 ( .A1(i_cmd[118]), .B1(n11706), .B2(n10322), .ZN(
        n10992) );
  INR3D0BWP30P140LVT U10850 ( .A1(i_cmd[86]), .B1(n11700), .B2(n10309), .ZN(
        n10964) );
  AOI22D1BWP30P140LVT U10851 ( .A1(i_data_bus[448]), .A2(n10992), .B1(
        i_data_bus[320]), .B2(n10964), .ZN(n10306) );
  INR3D0BWP30P140LVT U10852 ( .A1(i_cmd[110]), .B1(n11698), .B2(n10322), .ZN(
        n10969) );
  INVD1BWP30P140LVT U10853 ( .I(i_cmd[166]), .ZN(n10303) );
  NR3D0P7BWP30P140LVT U10854 ( .A1(n11747), .A2(n10303), .A3(n10308), .ZN(
        n10965) );
  AOI22D1BWP30P140LVT U10855 ( .A1(i_data_bus[416]), .A2(n10969), .B1(
        i_data_bus[640]), .B2(n10965), .ZN(n10305) );
  INR3D0BWP30P140LVT U10856 ( .A1(i_cmd[190]), .B1(n11750), .B2(n10308), .ZN(
        n10988) );
  INR3D0BWP30P140LVT U10857 ( .A1(i_cmd[62]), .B1(n11032), .B2(n10323), .ZN(
        n10990) );
  AOI22D1BWP30P140LVT U10858 ( .A1(i_data_bus[736]), .A2(n10988), .B1(
        i_data_bus[224]), .B2(n10990), .ZN(n10304) );
  ND4D1BWP30P140LVT U10859 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(n10330) );
  INR3D0BWP30P140LVT U10860 ( .A1(i_cmd[14]), .B1(n11737), .B2(n10320), .ZN(
        n10979) );
  INR3D0BWP30P140LVT U10861 ( .A1(i_cmd[182]), .B1(n11748), .B2(n10308), .ZN(
        n10995) );
  AOI22D1BWP30P140LVT U10862 ( .A1(i_data_bus[32]), .A2(n10979), .B1(
        i_data_bus[704]), .B2(n10995), .ZN(n10315) );
  INR3D0BWP30P140LVT U10863 ( .A1(i_cmd[142]), .B1(n11701), .B2(n10316), .ZN(
        n10958) );
  INR3D0BWP30P140LVT U10864 ( .A1(i_cmd[78]), .B1(n11711), .B2(n10309), .ZN(
        n10980) );
  AOI22D1BWP30P140LVT U10865 ( .A1(i_data_bus[544]), .A2(n10958), .B1(
        i_data_bus[288]), .B2(n10980), .ZN(n10314) );
  NR3D0P7BWP30P140LVT U10866 ( .A1(n11705), .A2(n10310), .A3(n10322), .ZN(
        n10994) );
  INR3D0BWP30P140LVT U10867 ( .A1(i_cmd[214]), .B1(n11745), .B2(n10319), .ZN(
        n10993) );
  AOI22D1BWP30P140LVT U10868 ( .A1(i_data_bus[384]), .A2(n10994), .B1(
        i_data_bus[832]), .B2(n10993), .ZN(n10313) );
  INVD1BWP30P140LVT U10869 ( .I(i_cmd[6]), .ZN(n10311) );
  NR3D0P7BWP30P140LVT U10870 ( .A1(n11703), .A2(n10311), .A3(n10320), .ZN(
        n10967) );
  INR3D0BWP30P140LVT U10871 ( .A1(i_cmd[54]), .B1(n11030), .B2(n10323), .ZN(
        n10983) );
  AOI22D1BWP30P140LVT U10872 ( .A1(i_data_bus[0]), .A2(n10967), .B1(
        i_data_bus[192]), .B2(n10983), .ZN(n10312) );
  ND4D1BWP30P140LVT U10873 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(n10329) );
  NR3D0P7BWP30P140LVT U10874 ( .A1(n11713), .A2(n10317), .A3(n10316), .ZN(
        n10957) );
  INVD1BWP30P140LVT U10875 ( .I(i_cmd[198]), .ZN(n10318) );
  NR3D0P7BWP30P140LVT U10876 ( .A1(n11754), .A2(n10318), .A3(n10319), .ZN(
        n10956) );
  AOI22D1BWP30P140LVT U10877 ( .A1(i_data_bus[512]), .A2(n10957), .B1(
        i_data_bus[768]), .B2(n10956), .ZN(n10327) );
  INR3D0BWP30P140LVT U10878 ( .A1(i_cmd[30]), .B1(n11726), .B2(n10320), .ZN(
        n10991) );
  INR3D0BWP30P140LVT U10879 ( .A1(i_cmd[222]), .B1(n11749), .B2(n10319), .ZN(
        n10982) );
  AOI22D1BWP30P140LVT U10880 ( .A1(i_data_bus[96]), .A2(n10991), .B1(
        i_data_bus[864]), .B2(n10982), .ZN(n10326) );
  INR3D0BWP30P140LVT U10881 ( .A1(i_cmd[22]), .B1(n11699), .B2(n10320), .ZN(
        n10959) );
  NR3D0P7BWP30P140LVT U10882 ( .A1(n11721), .A2(n10321), .A3(n10323), .ZN(
        n10966) );
  AOI22D1BWP30P140LVT U10883 ( .A1(i_data_bus[64]), .A2(n10959), .B1(
        i_data_bus[128]), .B2(n10966), .ZN(n10325) );
  INR3D0BWP30P140LVT U10884 ( .A1(i_cmd[126]), .B1(n11719), .B2(n10322), .ZN(
        n10989) );
  INR3D0BWP30P140LVT U10885 ( .A1(i_cmd[46]), .B1(n11023), .B2(n10323), .ZN(
        n10976) );
  AOI22D1BWP30P140LVT U10886 ( .A1(i_data_bus[480]), .A2(n10989), .B1(
        i_data_bus[160]), .B2(n10976), .ZN(n10324) );
  ND4D1BWP30P140LVT U10887 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10324), .ZN(n10328) );
  OR4D1BWP30P140LVT U10888 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .Z(o_data_bus[192]) );
  AOI22D1BWP30P140LVT U10889 ( .A1(i_data_bus[897]), .A2(n10952), .B1(
        i_data_bus[993]), .B2(n10955), .ZN(n10335) );
  AOI22D1BWP30P140LVT U10890 ( .A1(i_data_bus[961]), .A2(n10953), .B1(
        i_data_bus[929]), .B2(n10954), .ZN(n10334) );
  AOI22D1BWP30P140LVT U10891 ( .A1(i_data_bus[193]), .A2(n10983), .B1(
        i_data_bus[833]), .B2(n10993), .ZN(n10333) );
  AOI22D1BWP30P140LVT U10892 ( .A1(i_data_bus[609]), .A2(n10971), .B1(
        i_data_bus[353]), .B2(n10978), .ZN(n10332) );
  ND4D1BWP30P140LVT U10893 ( .A1(n10335), .A2(n10334), .A3(n10333), .A4(n10332), .ZN(n10351) );
  AOI22D1BWP30P140LVT U10894 ( .A1(i_data_bus[65]), .A2(n10959), .B1(
        i_data_bus[417]), .B2(n10969), .ZN(n10339) );
  AOI22D1BWP30P140LVT U10895 ( .A1(i_data_bus[289]), .A2(n10980), .B1(
        i_data_bus[321]), .B2(n10964), .ZN(n10338) );
  AOI22D1BWP30P140LVT U10896 ( .A1(i_data_bus[97]), .A2(n10991), .B1(
        i_data_bus[769]), .B2(n10956), .ZN(n10337) );
  AOI22D1BWP30P140LVT U10897 ( .A1(i_data_bus[513]), .A2(n10957), .B1(
        i_data_bus[673]), .B2(n10977), .ZN(n10336) );
  ND4D1BWP30P140LVT U10898 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(n10350) );
  AOI22D1BWP30P140LVT U10899 ( .A1(i_data_bus[1]), .A2(n10967), .B1(
        i_data_bus[257]), .B2(n10968), .ZN(n10343) );
  AOI22D1BWP30P140LVT U10900 ( .A1(i_data_bus[33]), .A2(n10979), .B1(
        i_data_bus[449]), .B2(n10992), .ZN(n10342) );
  AOI22D1BWP30P140LVT U10901 ( .A1(i_data_bus[705]), .A2(n10995), .B1(
        i_data_bus[865]), .B2(n10982), .ZN(n10341) );
  AOI22D1BWP30P140LVT U10902 ( .A1(i_data_bus[577]), .A2(n10981), .B1(
        i_data_bus[161]), .B2(n10976), .ZN(n10340) );
  ND4D1BWP30P140LVT U10903 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(n10349) );
  AOI22D1BWP30P140LVT U10904 ( .A1(i_data_bus[641]), .A2(n10965), .B1(
        i_data_bus[481]), .B2(n10989), .ZN(n10347) );
  AOI22D1BWP30P140LVT U10905 ( .A1(i_data_bus[385]), .A2(n10994), .B1(
        i_data_bus[737]), .B2(n10988), .ZN(n10346) );
  AOI22D1BWP30P140LVT U10906 ( .A1(i_data_bus[801]), .A2(n10970), .B1(
        i_data_bus[225]), .B2(n10990), .ZN(n10345) );
  AOI22D1BWP30P140LVT U10907 ( .A1(i_data_bus[545]), .A2(n10958), .B1(
        i_data_bus[129]), .B2(n10966), .ZN(n10344) );
  ND4D1BWP30P140LVT U10908 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(n10348) );
  OR4D1BWP30P140LVT U10909 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .Z(o_data_bus[193]) );
  AOI22D1BWP30P140LVT U10910 ( .A1(i_data_bus[962]), .A2(n10953), .B1(
        i_data_bus[930]), .B2(n10954), .ZN(n10355) );
  AOI22D1BWP30P140LVT U10911 ( .A1(i_data_bus[898]), .A2(n10952), .B1(
        i_data_bus[994]), .B2(n10955), .ZN(n10354) );
  AOI22D1BWP30P140LVT U10912 ( .A1(i_data_bus[674]), .A2(n10977), .B1(
        i_data_bus[770]), .B2(n10956), .ZN(n10353) );
  AOI22D1BWP30P140LVT U10913 ( .A1(i_data_bus[98]), .A2(n10991), .B1(
        i_data_bus[226]), .B2(n10990), .ZN(n10352) );
  ND4D1BWP30P140LVT U10914 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(n10371) );
  AOI22D1BWP30P140LVT U10915 ( .A1(i_data_bus[546]), .A2(n10958), .B1(
        i_data_bus[706]), .B2(n10995), .ZN(n10359) );
  AOI22D1BWP30P140LVT U10916 ( .A1(i_data_bus[610]), .A2(n10971), .B1(
        i_data_bus[834]), .B2(n10993), .ZN(n10358) );
  AOI22D1BWP30P140LVT U10917 ( .A1(i_data_bus[66]), .A2(n10959), .B1(
        i_data_bus[514]), .B2(n10957), .ZN(n10357) );
  AOI22D1BWP30P140LVT U10918 ( .A1(i_data_bus[34]), .A2(n10979), .B1(
        i_data_bus[354]), .B2(n10978), .ZN(n10356) );
  ND4D1BWP30P140LVT U10919 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(n10370) );
  AOI22D1BWP30P140LVT U10920 ( .A1(i_data_bus[290]), .A2(n10980), .B1(
        i_data_bus[802]), .B2(n10970), .ZN(n10363) );
  AOI22D1BWP30P140LVT U10921 ( .A1(i_data_bus[162]), .A2(n10976), .B1(
        i_data_bus[258]), .B2(n10968), .ZN(n10362) );
  AOI22D1BWP30P140LVT U10922 ( .A1(i_data_bus[194]), .A2(n10983), .B1(
        i_data_bus[322]), .B2(n10964), .ZN(n10361) );
  AOI22D1BWP30P140LVT U10923 ( .A1(i_data_bus[2]), .A2(n10967), .B1(
        i_data_bus[418]), .B2(n10969), .ZN(n10360) );
  ND4D1BWP30P140LVT U10924 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(n10369) );
  AOI22D1BWP30P140LVT U10925 ( .A1(i_data_bus[578]), .A2(n10981), .B1(
        i_data_bus[866]), .B2(n10982), .ZN(n10367) );
  AOI22D1BWP30P140LVT U10926 ( .A1(i_data_bus[386]), .A2(n10994), .B1(
        i_data_bus[738]), .B2(n10988), .ZN(n10366) );
  AOI22D1BWP30P140LVT U10927 ( .A1(i_data_bus[450]), .A2(n10992), .B1(
        i_data_bus[130]), .B2(n10966), .ZN(n10365) );
  AOI22D1BWP30P140LVT U10928 ( .A1(i_data_bus[482]), .A2(n10989), .B1(
        i_data_bus[642]), .B2(n10965), .ZN(n10364) );
  ND4D1BWP30P140LVT U10929 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(n10368) );
  OR4D1BWP30P140LVT U10930 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .Z(o_data_bus[194]) );
  AOI22D1BWP30P140LVT U10931 ( .A1(i_data_bus[963]), .A2(n10953), .B1(
        i_data_bus[995]), .B2(n10955), .ZN(n10375) );
  AOI22D1BWP30P140LVT U10932 ( .A1(i_data_bus[899]), .A2(n10952), .B1(
        i_data_bus[931]), .B2(n10954), .ZN(n10374) );
  AOI22D1BWP30P140LVT U10933 ( .A1(i_data_bus[3]), .A2(n10967), .B1(
        i_data_bus[323]), .B2(n10964), .ZN(n10373) );
  AOI22D1BWP30P140LVT U10934 ( .A1(i_data_bus[99]), .A2(n10991), .B1(
        i_data_bus[387]), .B2(n10994), .ZN(n10372) );
  ND4D1BWP30P140LVT U10935 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(n10391) );
  AOI22D1BWP30P140LVT U10936 ( .A1(i_data_bus[67]), .A2(n10959), .B1(
        i_data_bus[483]), .B2(n10989), .ZN(n10379) );
  AOI22D1BWP30P140LVT U10937 ( .A1(i_data_bus[163]), .A2(n10976), .B1(
        i_data_bus[707]), .B2(n10995), .ZN(n10378) );
  AOI22D1BWP30P140LVT U10938 ( .A1(i_data_bus[547]), .A2(n10958), .B1(
        i_data_bus[643]), .B2(n10965), .ZN(n10377) );
  AOI22D1BWP30P140LVT U10939 ( .A1(i_data_bus[771]), .A2(n10956), .B1(
        i_data_bus[867]), .B2(n10982), .ZN(n10376) );
  ND4D1BWP30P140LVT U10940 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(n10390) );
  AOI22D1BWP30P140LVT U10941 ( .A1(i_data_bus[675]), .A2(n10977), .B1(
        i_data_bus[451]), .B2(n10992), .ZN(n10383) );
  AOI22D1BWP30P140LVT U10942 ( .A1(i_data_bus[739]), .A2(n10988), .B1(
        i_data_bus[227]), .B2(n10990), .ZN(n10382) );
  AOI22D1BWP30P140LVT U10943 ( .A1(i_data_bus[355]), .A2(n10978), .B1(
        i_data_bus[803]), .B2(n10970), .ZN(n10381) );
  AOI22D1BWP30P140LVT U10944 ( .A1(i_data_bus[611]), .A2(n10971), .B1(
        i_data_bus[259]), .B2(n10968), .ZN(n10380) );
  ND4D1BWP30P140LVT U10945 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(n10389) );
  AOI22D1BWP30P140LVT U10946 ( .A1(i_data_bus[579]), .A2(n10981), .B1(
        i_data_bus[835]), .B2(n10993), .ZN(n10387) );
  AOI22D1BWP30P140LVT U10947 ( .A1(i_data_bus[515]), .A2(n10957), .B1(
        i_data_bus[35]), .B2(n10979), .ZN(n10386) );
  AOI22D1BWP30P140LVT U10948 ( .A1(i_data_bus[419]), .A2(n10969), .B1(
        i_data_bus[291]), .B2(n10980), .ZN(n10385) );
  AOI22D1BWP30P140LVT U10949 ( .A1(i_data_bus[131]), .A2(n10966), .B1(
        i_data_bus[195]), .B2(n10983), .ZN(n10384) );
  ND4D1BWP30P140LVT U10950 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(n10388) );
  OR4D1BWP30P140LVT U10951 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .Z(o_data_bus[195]) );
  AOI22D1BWP30P140LVT U10952 ( .A1(i_data_bus[964]), .A2(n10953), .B1(
        i_data_bus[996]), .B2(n10955), .ZN(n10395) );
  AOI22D1BWP30P140LVT U10953 ( .A1(i_data_bus[932]), .A2(n10954), .B1(
        i_data_bus[900]), .B2(n10952), .ZN(n10394) );
  AOI22D1BWP30P140LVT U10954 ( .A1(i_data_bus[740]), .A2(n10988), .B1(
        i_data_bus[676]), .B2(n10977), .ZN(n10393) );
  AOI22D1BWP30P140LVT U10955 ( .A1(i_data_bus[100]), .A2(n10991), .B1(
        i_data_bus[196]), .B2(n10983), .ZN(n10392) );
  ND4D1BWP30P140LVT U10956 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(n10411) );
  AOI22D1BWP30P140LVT U10957 ( .A1(i_data_bus[548]), .A2(n10958), .B1(
        i_data_bus[420]), .B2(n10969), .ZN(n10399) );
  AOI22D1BWP30P140LVT U10958 ( .A1(i_data_bus[708]), .A2(n10995), .B1(
        i_data_bus[228]), .B2(n10990), .ZN(n10398) );
  AOI22D1BWP30P140LVT U10959 ( .A1(i_data_bus[4]), .A2(n10967), .B1(
        i_data_bus[260]), .B2(n10968), .ZN(n10397) );
  AOI22D1BWP30P140LVT U10960 ( .A1(i_data_bus[292]), .A2(n10980), .B1(
        i_data_bus[644]), .B2(n10965), .ZN(n10396) );
  ND4D1BWP30P140LVT U10961 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(n10410) );
  AOI22D1BWP30P140LVT U10962 ( .A1(i_data_bus[324]), .A2(n10964), .B1(
        i_data_bus[356]), .B2(n10978), .ZN(n10403) );
  AOI22D1BWP30P140LVT U10963 ( .A1(i_data_bus[612]), .A2(n10971), .B1(
        i_data_bus[772]), .B2(n10956), .ZN(n10402) );
  AOI22D1BWP30P140LVT U10964 ( .A1(i_data_bus[132]), .A2(n10966), .B1(
        i_data_bus[388]), .B2(n10994), .ZN(n10401) );
  AOI22D1BWP30P140LVT U10965 ( .A1(i_data_bus[580]), .A2(n10981), .B1(
        i_data_bus[804]), .B2(n10970), .ZN(n10400) );
  ND4D1BWP30P140LVT U10966 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(n10409) );
  AOI22D1BWP30P140LVT U10967 ( .A1(i_data_bus[452]), .A2(n10992), .B1(
        i_data_bus[868]), .B2(n10982), .ZN(n10407) );
  AOI22D1BWP30P140LVT U10968 ( .A1(i_data_bus[164]), .A2(n10976), .B1(
        i_data_bus[836]), .B2(n10993), .ZN(n10406) );
  AOI22D1BWP30P140LVT U10969 ( .A1(i_data_bus[68]), .A2(n10959), .B1(
        i_data_bus[36]), .B2(n10979), .ZN(n10405) );
  AOI22D1BWP30P140LVT U10970 ( .A1(i_data_bus[516]), .A2(n10957), .B1(
        i_data_bus[484]), .B2(n10989), .ZN(n10404) );
  ND4D1BWP30P140LVT U10971 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(n10408) );
  OR4D1BWP30P140LVT U10972 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .Z(o_data_bus[196]) );
  AOI22D1BWP30P140LVT U10973 ( .A1(i_data_bus[933]), .A2(n10954), .B1(
        i_data_bus[997]), .B2(n10955), .ZN(n10415) );
  AOI22D1BWP30P140LVT U10974 ( .A1(i_data_bus[901]), .A2(n10952), .B1(
        i_data_bus[965]), .B2(n10953), .ZN(n10414) );
  AOI22D1BWP30P140LVT U10975 ( .A1(i_data_bus[517]), .A2(n10957), .B1(
        i_data_bus[261]), .B2(n10968), .ZN(n10413) );
  AOI22D1BWP30P140LVT U10976 ( .A1(i_data_bus[165]), .A2(n10976), .B1(
        i_data_bus[293]), .B2(n10980), .ZN(n10412) );
  ND4D1BWP30P140LVT U10977 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(n10431) );
  AOI22D1BWP30P140LVT U10978 ( .A1(i_data_bus[613]), .A2(n10971), .B1(
        i_data_bus[837]), .B2(n10993), .ZN(n10419) );
  AOI22D1BWP30P140LVT U10979 ( .A1(i_data_bus[805]), .A2(n10970), .B1(
        i_data_bus[741]), .B2(n10988), .ZN(n10418) );
  AOI22D1BWP30P140LVT U10980 ( .A1(i_data_bus[69]), .A2(n10959), .B1(
        i_data_bus[485]), .B2(n10989), .ZN(n10417) );
  AOI22D1BWP30P140LVT U10981 ( .A1(i_data_bus[709]), .A2(n10995), .B1(
        i_data_bus[133]), .B2(n10966), .ZN(n10416) );
  ND4D1BWP30P140LVT U10982 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(n10430) );
  AOI22D1BWP30P140LVT U10983 ( .A1(i_data_bus[869]), .A2(n10982), .B1(
        i_data_bus[325]), .B2(n10964), .ZN(n10423) );
  AOI22D1BWP30P140LVT U10984 ( .A1(i_data_bus[197]), .A2(n10983), .B1(
        i_data_bus[645]), .B2(n10965), .ZN(n10422) );
  AOI22D1BWP30P140LVT U10985 ( .A1(i_data_bus[581]), .A2(n10981), .B1(
        i_data_bus[773]), .B2(n10956), .ZN(n10421) );
  AOI22D1BWP30P140LVT U10986 ( .A1(i_data_bus[453]), .A2(n10992), .B1(
        i_data_bus[389]), .B2(n10994), .ZN(n10420) );
  ND4D1BWP30P140LVT U10987 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(n10429) );
  AOI22D1BWP30P140LVT U10988 ( .A1(i_data_bus[37]), .A2(n10979), .B1(
        i_data_bus[101]), .B2(n10991), .ZN(n10427) );
  AOI22D1BWP30P140LVT U10989 ( .A1(i_data_bus[357]), .A2(n10978), .B1(
        i_data_bus[229]), .B2(n10990), .ZN(n10426) );
  AOI22D1BWP30P140LVT U10990 ( .A1(i_data_bus[5]), .A2(n10967), .B1(
        i_data_bus[421]), .B2(n10969), .ZN(n10425) );
  AOI22D1BWP30P140LVT U10991 ( .A1(i_data_bus[549]), .A2(n10958), .B1(
        i_data_bus[677]), .B2(n10977), .ZN(n10424) );
  ND4D1BWP30P140LVT U10992 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(n10428) );
  OR4D1BWP30P140LVT U10993 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .Z(o_data_bus[197]) );
  AOI22D1BWP30P140LVT U10994 ( .A1(i_data_bus[324]), .A2(n12508), .B1(
        i_data_bus[388]), .B2(n12506), .ZN(n10435) );
  AOI22D1BWP30P140LVT U10995 ( .A1(i_data_bus[516]), .A2(n12477), .B1(
        i_data_bus[36]), .B2(n12483), .ZN(n10434) );
  AOI22D1BWP30P140LVT U10996 ( .A1(i_data_bus[132]), .A2(n12502), .B1(
        i_data_bus[484]), .B2(n12494), .ZN(n10433) );
  AOI22D1BWP30P140LVT U10997 ( .A1(i_data_bus[580]), .A2(n12480), .B1(
        i_data_bus[420]), .B2(n12481), .ZN(n10432) );
  ND4D1BWP30P140LVT U10998 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(n10451) );
  AOI22D1BWP30P140LVT U10999 ( .A1(i_data_bus[4]), .A2(n12490), .B1(
        i_data_bus[452]), .B2(n12507), .ZN(n10439) );
  AOI22D1BWP30P140LVT U11000 ( .A1(i_data_bus[932]), .A2(n12492), .B1(
        i_data_bus[228]), .B2(n12493), .ZN(n10438) );
  AOI22D1BWP30P140LVT U11001 ( .A1(i_data_bus[100]), .A2(n12489), .B1(
        i_data_bus[164]), .B2(n12501), .ZN(n10437) );
  AOI22D1BWP30P140LVT U11002 ( .A1(i_data_bus[964]), .A2(n12482), .B1(
        i_data_bus[356]), .B2(n12491), .ZN(n10436) );
  ND4D1BWP30P140LVT U11003 ( .A1(n10439), .A2(n10438), .A3(n10437), .A4(n10436), .ZN(n10450) );
  AOI22D1BWP30P140LVT U11004 ( .A1(i_data_bus[68]), .A2(n12478), .B1(
        i_data_bus[292]), .B2(n12505), .ZN(n10443) );
  AOI22D1BWP30P140LVT U11005 ( .A1(i_data_bus[612]), .A2(n12504), .B1(
        i_data_bus[900]), .B2(n12484), .ZN(n10442) );
  AOI22D1BWP30P140LVT U11006 ( .A1(i_data_bus[548]), .A2(n12479), .B1(
        i_data_bus[196]), .B2(n12495), .ZN(n10441) );
  AOI22D1BWP30P140LVT U11007 ( .A1(i_data_bus[996]), .A2(n12496), .B1(
        i_data_bus[260]), .B2(n12503), .ZN(n10440) );
  ND4D1BWP30P140LVT U11008 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(n10449) );
  AOI22D1BWP30P140LVT U11009 ( .A1(i_data_bus[868]), .A2(n12513), .B1(
        i_data_bus[644]), .B2(n12520), .ZN(n10447) );
  AOI22D1BWP30P140LVT U11010 ( .A1(i_data_bus[772]), .A2(n12516), .B1(
        i_data_bus[836]), .B2(n12514), .ZN(n10446) );
  AOI22D1BWP30P140LVT U11011 ( .A1(i_data_bus[740]), .A2(n12518), .B1(
        i_data_bus[676]), .B2(n12515), .ZN(n10445) );
  AOI22D1BWP30P140LVT U11012 ( .A1(i_data_bus[708]), .A2(n12519), .B1(
        i_data_bus[804]), .B2(n12517), .ZN(n10444) );
  ND4D1BWP30P140LVT U11013 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(n10448) );
  OR4D1BWP30P140LVT U11014 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .Z(o_data_bus[132]) );
  AOI22D1BWP30P140LVT U11015 ( .A1(i_data_bus[934]), .A2(n10954), .B1(
        i_data_bus[902]), .B2(n10952), .ZN(n10455) );
  AOI22D1BWP30P140LVT U11016 ( .A1(i_data_bus[966]), .A2(n10953), .B1(
        i_data_bus[998]), .B2(n10955), .ZN(n10454) );
  AOI22D1BWP30P140LVT U11017 ( .A1(i_data_bus[6]), .A2(n10967), .B1(
        i_data_bus[806]), .B2(n10970), .ZN(n10453) );
  AOI22D1BWP30P140LVT U11018 ( .A1(i_data_bus[742]), .A2(n10988), .B1(
        i_data_bus[326]), .B2(n10964), .ZN(n10452) );
  ND4D1BWP30P140LVT U11019 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(n10471) );
  AOI22D1BWP30P140LVT U11020 ( .A1(i_data_bus[70]), .A2(n10959), .B1(
        i_data_bus[678]), .B2(n10977), .ZN(n10459) );
  AOI22D1BWP30P140LVT U11021 ( .A1(i_data_bus[550]), .A2(n10958), .B1(
        i_data_bus[710]), .B2(n10995), .ZN(n10458) );
  AOI22D1BWP30P140LVT U11022 ( .A1(i_data_bus[38]), .A2(n10979), .B1(
        i_data_bus[134]), .B2(n10966), .ZN(n10457) );
  AOI22D1BWP30P140LVT U11023 ( .A1(i_data_bus[486]), .A2(n10989), .B1(
        i_data_bus[230]), .B2(n10990), .ZN(n10456) );
  ND4D1BWP30P140LVT U11024 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(n10470) );
  AOI22D1BWP30P140LVT U11025 ( .A1(i_data_bus[838]), .A2(n10993), .B1(
        i_data_bus[166]), .B2(n10976), .ZN(n10463) );
  AOI22D1BWP30P140LVT U11026 ( .A1(i_data_bus[582]), .A2(n10981), .B1(
        i_data_bus[454]), .B2(n10992), .ZN(n10462) );
  AOI22D1BWP30P140LVT U11027 ( .A1(i_data_bus[870]), .A2(n10982), .B1(
        i_data_bus[294]), .B2(n10980), .ZN(n10461) );
  AOI22D1BWP30P140LVT U11028 ( .A1(i_data_bus[102]), .A2(n10991), .B1(
        i_data_bus[358]), .B2(n10978), .ZN(n10460) );
  ND4D1BWP30P140LVT U11029 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(n10469) );
  AOI22D1BWP30P140LVT U11030 ( .A1(i_data_bus[646]), .A2(n10965), .B1(
        i_data_bus[774]), .B2(n10956), .ZN(n10467) );
  AOI22D1BWP30P140LVT U11031 ( .A1(i_data_bus[390]), .A2(n10994), .B1(
        i_data_bus[198]), .B2(n10983), .ZN(n10466) );
  AOI22D1BWP30P140LVT U11032 ( .A1(i_data_bus[614]), .A2(n10971), .B1(
        i_data_bus[262]), .B2(n10968), .ZN(n10465) );
  AOI22D1BWP30P140LVT U11033 ( .A1(i_data_bus[518]), .A2(n10957), .B1(
        i_data_bus[422]), .B2(n10969), .ZN(n10464) );
  ND4D1BWP30P140LVT U11034 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(n10468) );
  OR4D1BWP30P140LVT U11035 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .Z(o_data_bus[198]) );
  AOI22D1BWP30P140LVT U11036 ( .A1(i_data_bus[903]), .A2(n10952), .B1(
        i_data_bus[935]), .B2(n10954), .ZN(n10475) );
  AOI22D1BWP30P140LVT U11037 ( .A1(i_data_bus[967]), .A2(n10953), .B1(
        i_data_bus[999]), .B2(n10955), .ZN(n10474) );
  AOI22D1BWP30P140LVT U11038 ( .A1(i_data_bus[615]), .A2(n10971), .B1(
        i_data_bus[487]), .B2(n10989), .ZN(n10473) );
  AOI22D1BWP30P140LVT U11039 ( .A1(i_data_bus[167]), .A2(n10976), .B1(
        i_data_bus[423]), .B2(n10969), .ZN(n10472) );
  ND4D1BWP30P140LVT U11040 ( .A1(n10475), .A2(n10474), .A3(n10473), .A4(n10472), .ZN(n10491) );
  AOI22D1BWP30P140LVT U11041 ( .A1(i_data_bus[7]), .A2(n10967), .B1(
        i_data_bus[327]), .B2(n10964), .ZN(n10479) );
  AOI22D1BWP30P140LVT U11042 ( .A1(i_data_bus[519]), .A2(n10957), .B1(
        i_data_bus[455]), .B2(n10992), .ZN(n10478) );
  AOI22D1BWP30P140LVT U11043 ( .A1(i_data_bus[103]), .A2(n10991), .B1(
        i_data_bus[839]), .B2(n10993), .ZN(n10477) );
  AOI22D1BWP30P140LVT U11044 ( .A1(i_data_bus[71]), .A2(n10959), .B1(
        i_data_bus[775]), .B2(n10956), .ZN(n10476) );
  ND4D1BWP30P140LVT U11045 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(n10490) );
  AOI22D1BWP30P140LVT U11046 ( .A1(i_data_bus[39]), .A2(n10979), .B1(
        i_data_bus[295]), .B2(n10980), .ZN(n10483) );
  AOI22D1BWP30P140LVT U11047 ( .A1(i_data_bus[391]), .A2(n10994), .B1(
        i_data_bus[199]), .B2(n10983), .ZN(n10482) );
  AOI22D1BWP30P140LVT U11048 ( .A1(i_data_bus[583]), .A2(n10981), .B1(
        i_data_bus[359]), .B2(n10978), .ZN(n10481) );
  AOI22D1BWP30P140LVT U11049 ( .A1(i_data_bus[679]), .A2(n10977), .B1(
        i_data_bus[807]), .B2(n10970), .ZN(n10480) );
  ND4D1BWP30P140LVT U11050 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(n10489) );
  AOI22D1BWP30P140LVT U11051 ( .A1(i_data_bus[263]), .A2(n10968), .B1(
        i_data_bus[711]), .B2(n10995), .ZN(n10487) );
  AOI22D1BWP30P140LVT U11052 ( .A1(i_data_bus[871]), .A2(n10982), .B1(
        i_data_bus[231]), .B2(n10990), .ZN(n10486) );
  AOI22D1BWP30P140LVT U11053 ( .A1(i_data_bus[743]), .A2(n10988), .B1(
        i_data_bus[135]), .B2(n10966), .ZN(n10485) );
  AOI22D1BWP30P140LVT U11054 ( .A1(i_data_bus[551]), .A2(n10958), .B1(
        i_data_bus[647]), .B2(n10965), .ZN(n10484) );
  ND4D1BWP30P140LVT U11055 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(n10488) );
  OR4D1BWP30P140LVT U11056 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .Z(o_data_bus[199]) );
  AOI22D1BWP30P140LVT U11057 ( .A1(i_data_bus[936]), .A2(n10954), .B1(
        i_data_bus[904]), .B2(n10952), .ZN(n10495) );
  AOI22D1BWP30P140LVT U11058 ( .A1(i_data_bus[968]), .A2(n10953), .B1(
        i_data_bus[1000]), .B2(n10955), .ZN(n10494) );
  AOI22D1BWP30P140LVT U11059 ( .A1(i_data_bus[264]), .A2(n10968), .B1(
        i_data_bus[392]), .B2(n10994), .ZN(n10493) );
  AOI22D1BWP30P140LVT U11060 ( .A1(i_data_bus[488]), .A2(n10989), .B1(
        i_data_bus[232]), .B2(n10990), .ZN(n10492) );
  ND4D1BWP30P140LVT U11061 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(n10511) );
  AOI22D1BWP30P140LVT U11062 ( .A1(i_data_bus[72]), .A2(n10959), .B1(
        i_data_bus[168]), .B2(n10976), .ZN(n10499) );
  AOI22D1BWP30P140LVT U11063 ( .A1(i_data_bus[8]), .A2(n10967), .B1(
        i_data_bus[872]), .B2(n10982), .ZN(n10498) );
  AOI22D1BWP30P140LVT U11064 ( .A1(i_data_bus[520]), .A2(n10957), .B1(
        i_data_bus[200]), .B2(n10983), .ZN(n10497) );
  AOI22D1BWP30P140LVT U11065 ( .A1(i_data_bus[456]), .A2(n10992), .B1(
        i_data_bus[296]), .B2(n10980), .ZN(n10496) );
  ND4D1BWP30P140LVT U11066 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(n10510) );
  AOI22D1BWP30P140LVT U11067 ( .A1(i_data_bus[840]), .A2(n10993), .B1(
        i_data_bus[648]), .B2(n10965), .ZN(n10503) );
  AOI22D1BWP30P140LVT U11068 ( .A1(i_data_bus[328]), .A2(n10964), .B1(
        i_data_bus[360]), .B2(n10978), .ZN(n10502) );
  AOI22D1BWP30P140LVT U11069 ( .A1(i_data_bus[424]), .A2(n10969), .B1(
        i_data_bus[712]), .B2(n10995), .ZN(n10501) );
  AOI22D1BWP30P140LVT U11070 ( .A1(i_data_bus[680]), .A2(n10977), .B1(
        i_data_bus[776]), .B2(n10956), .ZN(n10500) );
  ND4D1BWP30P140LVT U11071 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(n10509) );
  AOI22D1BWP30P140LVT U11072 ( .A1(i_data_bus[744]), .A2(n10988), .B1(
        i_data_bus[808]), .B2(n10970), .ZN(n10507) );
  AOI22D1BWP30P140LVT U11073 ( .A1(i_data_bus[616]), .A2(n10971), .B1(
        i_data_bus[40]), .B2(n10979), .ZN(n10506) );
  AOI22D1BWP30P140LVT U11074 ( .A1(i_data_bus[104]), .A2(n10991), .B1(
        i_data_bus[552]), .B2(n10958), .ZN(n10505) );
  AOI22D1BWP30P140LVT U11075 ( .A1(i_data_bus[584]), .A2(n10981), .B1(
        i_data_bus[136]), .B2(n10966), .ZN(n10504) );
  ND4D1BWP30P140LVT U11076 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(n10508) );
  OR4D1BWP30P140LVT U11077 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .Z(o_data_bus[200]) );
  AOI22D1BWP30P140LVT U11078 ( .A1(i_data_bus[969]), .A2(n10953), .B1(
        i_data_bus[1001]), .B2(n10955), .ZN(n10515) );
  AOI22D1BWP30P140LVT U11079 ( .A1(i_data_bus[905]), .A2(n10952), .B1(
        i_data_bus[937]), .B2(n10954), .ZN(n10514) );
  AOI22D1BWP30P140LVT U11080 ( .A1(i_data_bus[9]), .A2(n10967), .B1(
        i_data_bus[105]), .B2(n10991), .ZN(n10513) );
  AOI22D1BWP30P140LVT U11081 ( .A1(i_data_bus[489]), .A2(n10989), .B1(
        i_data_bus[425]), .B2(n10969), .ZN(n10512) );
  ND4D1BWP30P140LVT U11082 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(n10531) );
  AOI22D1BWP30P140LVT U11083 ( .A1(i_data_bus[265]), .A2(n10968), .B1(
        i_data_bus[777]), .B2(n10956), .ZN(n10519) );
  AOI22D1BWP30P140LVT U11084 ( .A1(i_data_bus[41]), .A2(n10979), .B1(
        i_data_bus[137]), .B2(n10966), .ZN(n10518) );
  AOI22D1BWP30P140LVT U11085 ( .A1(i_data_bus[585]), .A2(n10981), .B1(
        i_data_bus[329]), .B2(n10964), .ZN(n10517) );
  AOI22D1BWP30P140LVT U11086 ( .A1(i_data_bus[713]), .A2(n10995), .B1(
        i_data_bus[457]), .B2(n10992), .ZN(n10516) );
  ND4D1BWP30P140LVT U11087 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(n10530) );
  AOI22D1BWP30P140LVT U11088 ( .A1(i_data_bus[201]), .A2(n10983), .B1(
        i_data_bus[393]), .B2(n10994), .ZN(n10523) );
  AOI22D1BWP30P140LVT U11089 ( .A1(i_data_bus[745]), .A2(n10988), .B1(
        i_data_bus[809]), .B2(n10970), .ZN(n10522) );
  AOI22D1BWP30P140LVT U11090 ( .A1(i_data_bus[841]), .A2(n10993), .B1(
        i_data_bus[649]), .B2(n10965), .ZN(n10521) );
  AOI22D1BWP30P140LVT U11091 ( .A1(i_data_bus[617]), .A2(n10971), .B1(
        i_data_bus[233]), .B2(n10990), .ZN(n10520) );
  ND4D1BWP30P140LVT U11092 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(n10529) );
  AOI22D1BWP30P140LVT U11093 ( .A1(i_data_bus[297]), .A2(n10980), .B1(
        i_data_bus[361]), .B2(n10978), .ZN(n10527) );
  AOI22D1BWP30P140LVT U11094 ( .A1(i_data_bus[553]), .A2(n10958), .B1(
        i_data_bus[169]), .B2(n10976), .ZN(n10526) );
  AOI22D1BWP30P140LVT U11095 ( .A1(i_data_bus[73]), .A2(n10959), .B1(
        i_data_bus[873]), .B2(n10982), .ZN(n10525) );
  AOI22D1BWP30P140LVT U11096 ( .A1(i_data_bus[521]), .A2(n10957), .B1(
        i_data_bus[681]), .B2(n10977), .ZN(n10524) );
  ND4D1BWP30P140LVT U11097 ( .A1(n10527), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(n10528) );
  OR4D1BWP30P140LVT U11098 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .Z(o_data_bus[201]) );
  AOI22D1BWP30P140LVT U11099 ( .A1(i_data_bus[970]), .A2(n10953), .B1(
        i_data_bus[906]), .B2(n10952), .ZN(n10535) );
  AOI22D1BWP30P140LVT U11100 ( .A1(i_data_bus[1002]), .A2(n10955), .B1(
        i_data_bus[938]), .B2(n10954), .ZN(n10534) );
  AOI22D1BWP30P140LVT U11101 ( .A1(i_data_bus[522]), .A2(n10957), .B1(
        i_data_bus[202]), .B2(n10983), .ZN(n10533) );
  AOI22D1BWP30P140LVT U11102 ( .A1(i_data_bus[490]), .A2(n10989), .B1(
        i_data_bus[682]), .B2(n10977), .ZN(n10532) );
  ND4D1BWP30P140LVT U11103 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(n10551) );
  AOI22D1BWP30P140LVT U11104 ( .A1(i_data_bus[42]), .A2(n10979), .B1(
        i_data_bus[650]), .B2(n10965), .ZN(n10539) );
  AOI22D1BWP30P140LVT U11105 ( .A1(i_data_bus[170]), .A2(n10976), .B1(
        i_data_bus[266]), .B2(n10968), .ZN(n10538) );
  AOI22D1BWP30P140LVT U11106 ( .A1(i_data_bus[554]), .A2(n10958), .B1(
        i_data_bus[74]), .B2(n10959), .ZN(n10537) );
  AOI22D1BWP30P140LVT U11107 ( .A1(i_data_bus[842]), .A2(n10993), .B1(
        i_data_bus[298]), .B2(n10980), .ZN(n10536) );
  ND4D1BWP30P140LVT U11108 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(n10550) );
  AOI22D1BWP30P140LVT U11109 ( .A1(i_data_bus[778]), .A2(n10956), .B1(
        i_data_bus[362]), .B2(n10978), .ZN(n10543) );
  AOI22D1BWP30P140LVT U11110 ( .A1(i_data_bus[458]), .A2(n10992), .B1(
        i_data_bus[138]), .B2(n10966), .ZN(n10542) );
  AOI22D1BWP30P140LVT U11111 ( .A1(i_data_bus[234]), .A2(n10990), .B1(
        i_data_bus[394]), .B2(n10994), .ZN(n10541) );
  AOI22D1BWP30P140LVT U11112 ( .A1(i_data_bus[586]), .A2(n10981), .B1(
        i_data_bus[330]), .B2(n10964), .ZN(n10540) );
  ND4D1BWP30P140LVT U11113 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(n10549) );
  AOI22D1BWP30P140LVT U11114 ( .A1(i_data_bus[10]), .A2(n10967), .B1(
        i_data_bus[426]), .B2(n10969), .ZN(n10547) );
  AOI22D1BWP30P140LVT U11115 ( .A1(i_data_bus[714]), .A2(n10995), .B1(
        i_data_bus[746]), .B2(n10988), .ZN(n10546) );
  AOI22D1BWP30P140LVT U11116 ( .A1(i_data_bus[618]), .A2(n10971), .B1(
        i_data_bus[874]), .B2(n10982), .ZN(n10545) );
  AOI22D1BWP30P140LVT U11117 ( .A1(i_data_bus[106]), .A2(n10991), .B1(
        i_data_bus[810]), .B2(n10970), .ZN(n10544) );
  ND4D1BWP30P140LVT U11118 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(n10548) );
  OR4D1BWP30P140LVT U11119 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .Z(o_data_bus[202]) );
  AOI22D1BWP30P140LVT U11120 ( .A1(i_data_bus[907]), .A2(n10952), .B1(
        i_data_bus[1003]), .B2(n10955), .ZN(n10555) );
  AOI22D1BWP30P140LVT U11121 ( .A1(i_data_bus[939]), .A2(n10954), .B1(
        i_data_bus[971]), .B2(n10953), .ZN(n10554) );
  AOI22D1BWP30P140LVT U11122 ( .A1(i_data_bus[811]), .A2(n10970), .B1(
        i_data_bus[331]), .B2(n10964), .ZN(n10553) );
  AOI22D1BWP30P140LVT U11123 ( .A1(i_data_bus[139]), .A2(n10966), .B1(
        i_data_bus[715]), .B2(n10995), .ZN(n10552) );
  ND4D1BWP30P140LVT U11124 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(n10571) );
  AOI22D1BWP30P140LVT U11125 ( .A1(i_data_bus[875]), .A2(n10982), .B1(
        i_data_bus[747]), .B2(n10988), .ZN(n10559) );
  AOI22D1BWP30P140LVT U11126 ( .A1(i_data_bus[75]), .A2(n10959), .B1(
        i_data_bus[235]), .B2(n10990), .ZN(n10558) );
  AOI22D1BWP30P140LVT U11127 ( .A1(i_data_bus[43]), .A2(n10979), .B1(
        i_data_bus[843]), .B2(n10993), .ZN(n10557) );
  AOI22D1BWP30P140LVT U11128 ( .A1(i_data_bus[587]), .A2(n10981), .B1(
        i_data_bus[427]), .B2(n10969), .ZN(n10556) );
  ND4D1BWP30P140LVT U11129 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(n10570) );
  AOI22D1BWP30P140LVT U11130 ( .A1(i_data_bus[619]), .A2(n10971), .B1(
        i_data_bus[555]), .B2(n10958), .ZN(n10563) );
  AOI22D1BWP30P140LVT U11131 ( .A1(i_data_bus[11]), .A2(n10967), .B1(
        i_data_bus[203]), .B2(n10983), .ZN(n10562) );
  AOI22D1BWP30P140LVT U11132 ( .A1(i_data_bus[107]), .A2(n10991), .B1(
        i_data_bus[299]), .B2(n10980), .ZN(n10561) );
  AOI22D1BWP30P140LVT U11133 ( .A1(i_data_bus[523]), .A2(n10957), .B1(
        i_data_bus[491]), .B2(n10989), .ZN(n10560) );
  ND4D1BWP30P140LVT U11134 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(n10569) );
  AOI22D1BWP30P140LVT U11135 ( .A1(i_data_bus[171]), .A2(n10976), .B1(
        i_data_bus[651]), .B2(n10965), .ZN(n10567) );
  AOI22D1BWP30P140LVT U11136 ( .A1(i_data_bus[363]), .A2(n10978), .B1(
        i_data_bus[459]), .B2(n10992), .ZN(n10566) );
  AOI22D1BWP30P140LVT U11137 ( .A1(i_data_bus[779]), .A2(n10956), .B1(
        i_data_bus[267]), .B2(n10968), .ZN(n10565) );
  AOI22D1BWP30P140LVT U11138 ( .A1(i_data_bus[395]), .A2(n10994), .B1(
        i_data_bus[683]), .B2(n10977), .ZN(n10564) );
  ND4D1BWP30P140LVT U11139 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(n10568) );
  OR4D1BWP30P140LVT U11140 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .Z(o_data_bus[203]) );
  AOI22D1BWP30P140LVT U11141 ( .A1(i_data_bus[908]), .A2(n10952), .B1(
        i_data_bus[1004]), .B2(n10955), .ZN(n10575) );
  AOI22D1BWP30P140LVT U11142 ( .A1(i_data_bus[940]), .A2(n10954), .B1(
        i_data_bus[972]), .B2(n10953), .ZN(n10574) );
  AOI22D1BWP30P140LVT U11143 ( .A1(i_data_bus[524]), .A2(n10957), .B1(
        i_data_bus[652]), .B2(n10965), .ZN(n10573) );
  AOI22D1BWP30P140LVT U11144 ( .A1(i_data_bus[716]), .A2(n10995), .B1(
        i_data_bus[268]), .B2(n10968), .ZN(n10572) );
  ND4D1BWP30P140LVT U11145 ( .A1(n10575), .A2(n10574), .A3(n10573), .A4(n10572), .ZN(n10591) );
  AOI22D1BWP30P140LVT U11146 ( .A1(i_data_bus[140]), .A2(n10966), .B1(
        i_data_bus[236]), .B2(n10990), .ZN(n10579) );
  AOI22D1BWP30P140LVT U11147 ( .A1(i_data_bus[556]), .A2(n10958), .B1(
        i_data_bus[460]), .B2(n10992), .ZN(n10578) );
  AOI22D1BWP30P140LVT U11148 ( .A1(i_data_bus[108]), .A2(n10991), .B1(
        i_data_bus[300]), .B2(n10980), .ZN(n10577) );
  AOI22D1BWP30P140LVT U11149 ( .A1(i_data_bus[428]), .A2(n10969), .B1(
        i_data_bus[844]), .B2(n10993), .ZN(n10576) );
  ND4D1BWP30P140LVT U11150 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(n10590) );
  AOI22D1BWP30P140LVT U11151 ( .A1(i_data_bus[780]), .A2(n10956), .B1(
        i_data_bus[332]), .B2(n10964), .ZN(n10583) );
  AOI22D1BWP30P140LVT U11152 ( .A1(i_data_bus[588]), .A2(n10981), .B1(
        i_data_bus[684]), .B2(n10977), .ZN(n10582) );
  AOI22D1BWP30P140LVT U11153 ( .A1(i_data_bus[620]), .A2(n10971), .B1(
        i_data_bus[876]), .B2(n10982), .ZN(n10581) );
  AOI22D1BWP30P140LVT U11154 ( .A1(i_data_bus[44]), .A2(n10979), .B1(
        i_data_bus[172]), .B2(n10976), .ZN(n10580) );
  ND4D1BWP30P140LVT U11155 ( .A1(n10583), .A2(n10582), .A3(n10581), .A4(n10580), .ZN(n10589) );
  AOI22D1BWP30P140LVT U11156 ( .A1(i_data_bus[204]), .A2(n10983), .B1(
        i_data_bus[492]), .B2(n10989), .ZN(n10587) );
  AOI22D1BWP30P140LVT U11157 ( .A1(i_data_bus[364]), .A2(n10978), .B1(
        i_data_bus[396]), .B2(n10994), .ZN(n10586) );
  AOI22D1BWP30P140LVT U11158 ( .A1(i_data_bus[76]), .A2(n10959), .B1(
        i_data_bus[812]), .B2(n10970), .ZN(n10585) );
  AOI22D1BWP30P140LVT U11159 ( .A1(i_data_bus[12]), .A2(n10967), .B1(
        i_data_bus[748]), .B2(n10988), .ZN(n10584) );
  ND4D1BWP30P140LVT U11160 ( .A1(n10587), .A2(n10586), .A3(n10585), .A4(n10584), .ZN(n10588) );
  OR4D1BWP30P140LVT U11161 ( .A1(n10591), .A2(n10590), .A3(n10589), .A4(n10588), .Z(o_data_bus[204]) );
  AOI22D1BWP30P140LVT U11162 ( .A1(i_data_bus[973]), .A2(n10953), .B1(
        i_data_bus[941]), .B2(n10954), .ZN(n10595) );
  AOI22D1BWP30P140LVT U11163 ( .A1(i_data_bus[909]), .A2(n10952), .B1(
        i_data_bus[1005]), .B2(n10955), .ZN(n10594) );
  AOI22D1BWP30P140LVT U11164 ( .A1(i_data_bus[77]), .A2(n10959), .B1(
        i_data_bus[749]), .B2(n10988), .ZN(n10593) );
  AOI22D1BWP30P140LVT U11165 ( .A1(i_data_bus[109]), .A2(n10991), .B1(
        i_data_bus[877]), .B2(n10982), .ZN(n10592) );
  ND4D1BWP30P140LVT U11166 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(n10611) );
  AOI22D1BWP30P140LVT U11167 ( .A1(i_data_bus[589]), .A2(n10981), .B1(
        i_data_bus[685]), .B2(n10977), .ZN(n10599) );
  AOI22D1BWP30P140LVT U11168 ( .A1(i_data_bus[365]), .A2(n10978), .B1(
        i_data_bus[781]), .B2(n10956), .ZN(n10598) );
  AOI22D1BWP30P140LVT U11169 ( .A1(i_data_bus[621]), .A2(n10971), .B1(
        i_data_bus[301]), .B2(n10980), .ZN(n10597) );
  AOI22D1BWP30P140LVT U11170 ( .A1(i_data_bus[237]), .A2(n10990), .B1(
        i_data_bus[653]), .B2(n10965), .ZN(n10596) );
  ND4D1BWP30P140LVT U11171 ( .A1(n10599), .A2(n10598), .A3(n10597), .A4(n10596), .ZN(n10610) );
  AOI22D1BWP30P140LVT U11172 ( .A1(i_data_bus[397]), .A2(n10994), .B1(
        i_data_bus[429]), .B2(n10969), .ZN(n10603) );
  AOI22D1BWP30P140LVT U11173 ( .A1(i_data_bus[845]), .A2(n10993), .B1(
        i_data_bus[813]), .B2(n10970), .ZN(n10602) );
  AOI22D1BWP30P140LVT U11174 ( .A1(i_data_bus[45]), .A2(n10979), .B1(
        i_data_bus[173]), .B2(n10976), .ZN(n10601) );
  AOI22D1BWP30P140LVT U11175 ( .A1(i_data_bus[525]), .A2(n10957), .B1(
        i_data_bus[269]), .B2(n10968), .ZN(n10600) );
  ND4D1BWP30P140LVT U11176 ( .A1(n10603), .A2(n10602), .A3(n10601), .A4(n10600), .ZN(n10609) );
  AOI22D1BWP30P140LVT U11177 ( .A1(i_data_bus[333]), .A2(n10964), .B1(
        i_data_bus[717]), .B2(n10995), .ZN(n10607) );
  AOI22D1BWP30P140LVT U11178 ( .A1(i_data_bus[13]), .A2(n10967), .B1(
        i_data_bus[461]), .B2(n10992), .ZN(n10606) );
  AOI22D1BWP30P140LVT U11179 ( .A1(i_data_bus[557]), .A2(n10958), .B1(
        i_data_bus[205]), .B2(n10983), .ZN(n10605) );
  AOI22D1BWP30P140LVT U11180 ( .A1(i_data_bus[493]), .A2(n10989), .B1(
        i_data_bus[141]), .B2(n10966), .ZN(n10604) );
  ND4D1BWP30P140LVT U11181 ( .A1(n10607), .A2(n10606), .A3(n10605), .A4(n10604), .ZN(n10608) );
  OR4D1BWP30P140LVT U11182 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .Z(o_data_bus[205]) );
  AOI22D1BWP30P140LVT U11183 ( .A1(i_data_bus[1006]), .A2(n10955), .B1(
        i_data_bus[974]), .B2(n10953), .ZN(n10615) );
  AOI22D1BWP30P140LVT U11184 ( .A1(i_data_bus[910]), .A2(n10952), .B1(
        i_data_bus[942]), .B2(n10954), .ZN(n10614) );
  AOI22D1BWP30P140LVT U11185 ( .A1(i_data_bus[46]), .A2(n10979), .B1(
        i_data_bus[206]), .B2(n10983), .ZN(n10613) );
  AOI22D1BWP30P140LVT U11186 ( .A1(i_data_bus[430]), .A2(n10969), .B1(
        i_data_bus[750]), .B2(n10988), .ZN(n10612) );
  ND4D1BWP30P140LVT U11187 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(n10631) );
  AOI22D1BWP30P140LVT U11188 ( .A1(i_data_bus[302]), .A2(n10980), .B1(
        i_data_bus[782]), .B2(n10956), .ZN(n10619) );
  AOI22D1BWP30P140LVT U11189 ( .A1(i_data_bus[590]), .A2(n10981), .B1(
        i_data_bus[558]), .B2(n10958), .ZN(n10618) );
  AOI22D1BWP30P140LVT U11190 ( .A1(i_data_bus[174]), .A2(n10976), .B1(
        i_data_bus[686]), .B2(n10977), .ZN(n10617) );
  AOI22D1BWP30P140LVT U11191 ( .A1(i_data_bus[622]), .A2(n10971), .B1(
        i_data_bus[238]), .B2(n10990), .ZN(n10616) );
  ND4D1BWP30P140LVT U11192 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(n10630) );
  AOI22D1BWP30P140LVT U11193 ( .A1(i_data_bus[78]), .A2(n10959), .B1(
        i_data_bus[366]), .B2(n10978), .ZN(n10623) );
  AOI22D1BWP30P140LVT U11194 ( .A1(i_data_bus[526]), .A2(n10957), .B1(
        i_data_bus[334]), .B2(n10964), .ZN(n10622) );
  AOI22D1BWP30P140LVT U11195 ( .A1(i_data_bus[14]), .A2(n10967), .B1(
        i_data_bus[270]), .B2(n10968), .ZN(n10621) );
  AOI22D1BWP30P140LVT U11196 ( .A1(i_data_bus[462]), .A2(n10992), .B1(
        i_data_bus[846]), .B2(n10993), .ZN(n10620) );
  ND4D1BWP30P140LVT U11197 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(n10629) );
  AOI22D1BWP30P140LVT U11198 ( .A1(i_data_bus[110]), .A2(n10991), .B1(
        i_data_bus[398]), .B2(n10994), .ZN(n10627) );
  AOI22D1BWP30P140LVT U11199 ( .A1(i_data_bus[814]), .A2(n10970), .B1(
        i_data_bus[878]), .B2(n10982), .ZN(n10626) );
  AOI22D1BWP30P140LVT U11200 ( .A1(i_data_bus[494]), .A2(n10989), .B1(
        i_data_bus[654]), .B2(n10965), .ZN(n10625) );
  AOI22D1BWP30P140LVT U11201 ( .A1(i_data_bus[142]), .A2(n10966), .B1(
        i_data_bus[718]), .B2(n10995), .ZN(n10624) );
  ND4D1BWP30P140LVT U11202 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(n10628) );
  OR4D1BWP30P140LVT U11203 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .Z(o_data_bus[206]) );
  AOI22D1BWP30P140LVT U11204 ( .A1(i_data_bus[1007]), .A2(n10955), .B1(
        i_data_bus[943]), .B2(n10954), .ZN(n10635) );
  AOI22D1BWP30P140LVT U11205 ( .A1(i_data_bus[975]), .A2(n10953), .B1(
        i_data_bus[911]), .B2(n10952), .ZN(n10634) );
  AOI22D1BWP30P140LVT U11206 ( .A1(i_data_bus[111]), .A2(n10991), .B1(
        i_data_bus[335]), .B2(n10964), .ZN(n10633) );
  AOI22D1BWP30P140LVT U11207 ( .A1(i_data_bus[271]), .A2(n10968), .B1(
        i_data_bus[815]), .B2(n10970), .ZN(n10632) );
  ND4D1BWP30P140LVT U11208 ( .A1(n10635), .A2(n10634), .A3(n10633), .A4(n10632), .ZN(n10651) );
  AOI22D1BWP30P140LVT U11209 ( .A1(i_data_bus[47]), .A2(n10979), .B1(
        i_data_bus[207]), .B2(n10983), .ZN(n10639) );
  AOI22D1BWP30P140LVT U11210 ( .A1(i_data_bus[79]), .A2(n10959), .B1(
        i_data_bus[431]), .B2(n10969), .ZN(n10638) );
  AOI22D1BWP30P140LVT U11211 ( .A1(i_data_bus[847]), .A2(n10993), .B1(
        i_data_bus[143]), .B2(n10966), .ZN(n10637) );
  AOI22D1BWP30P140LVT U11212 ( .A1(i_data_bus[15]), .A2(n10967), .B1(
        i_data_bus[175]), .B2(n10976), .ZN(n10636) );
  ND4D1BWP30P140LVT U11213 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(n10650) );
  AOI22D1BWP30P140LVT U11214 ( .A1(i_data_bus[463]), .A2(n10992), .B1(
        i_data_bus[399]), .B2(n10994), .ZN(n10643) );
  AOI22D1BWP30P140LVT U11215 ( .A1(i_data_bus[527]), .A2(n10957), .B1(
        i_data_bus[623]), .B2(n10971), .ZN(n10642) );
  AOI22D1BWP30P140LVT U11216 ( .A1(i_data_bus[559]), .A2(n10958), .B1(
        i_data_bus[303]), .B2(n10980), .ZN(n10641) );
  AOI22D1BWP30P140LVT U11217 ( .A1(i_data_bus[719]), .A2(n10995), .B1(
        i_data_bus[239]), .B2(n10990), .ZN(n10640) );
  ND4D1BWP30P140LVT U11218 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(n10649) );
  AOI22D1BWP30P140LVT U11219 ( .A1(i_data_bus[655]), .A2(n10965), .B1(
        i_data_bus[783]), .B2(n10956), .ZN(n10647) );
  AOI22D1BWP30P140LVT U11220 ( .A1(i_data_bus[495]), .A2(n10989), .B1(
        i_data_bus[879]), .B2(n10982), .ZN(n10646) );
  AOI22D1BWP30P140LVT U11221 ( .A1(i_data_bus[751]), .A2(n10988), .B1(
        i_data_bus[687]), .B2(n10977), .ZN(n10645) );
  AOI22D1BWP30P140LVT U11222 ( .A1(i_data_bus[591]), .A2(n10981), .B1(
        i_data_bus[367]), .B2(n10978), .ZN(n10644) );
  ND4D1BWP30P140LVT U11223 ( .A1(n10647), .A2(n10646), .A3(n10645), .A4(n10644), .ZN(n10648) );
  OR4D1BWP30P140LVT U11224 ( .A1(n10651), .A2(n10650), .A3(n10649), .A4(n10648), .Z(o_data_bus[207]) );
  AOI22D1BWP30P140LVT U11225 ( .A1(i_data_bus[944]), .A2(n10954), .B1(
        i_data_bus[976]), .B2(n10953), .ZN(n10655) );
  AOI22D1BWP30P140LVT U11226 ( .A1(i_data_bus[912]), .A2(n10952), .B1(
        i_data_bus[1008]), .B2(n10955), .ZN(n10654) );
  AOI22D1BWP30P140LVT U11227 ( .A1(i_data_bus[496]), .A2(n10989), .B1(
        i_data_bus[720]), .B2(n10995), .ZN(n10653) );
  AOI22D1BWP30P140LVT U11228 ( .A1(i_data_bus[528]), .A2(n10957), .B1(
        i_data_bus[144]), .B2(n10966), .ZN(n10652) );
  ND4D1BWP30P140LVT U11229 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(n10671) );
  AOI22D1BWP30P140LVT U11230 ( .A1(i_data_bus[80]), .A2(n10959), .B1(
        i_data_bus[112]), .B2(n10991), .ZN(n10659) );
  AOI22D1BWP30P140LVT U11231 ( .A1(i_data_bus[304]), .A2(n10980), .B1(
        i_data_bus[208]), .B2(n10983), .ZN(n10658) );
  AOI22D1BWP30P140LVT U11232 ( .A1(i_data_bus[784]), .A2(n10956), .B1(
        i_data_bus[400]), .B2(n10994), .ZN(n10657) );
  AOI22D1BWP30P140LVT U11233 ( .A1(i_data_bus[560]), .A2(n10958), .B1(
        i_data_bus[880]), .B2(n10982), .ZN(n10656) );
  ND4D1BWP30P140LVT U11234 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(n10670) );
  AOI22D1BWP30P140LVT U11235 ( .A1(i_data_bus[432]), .A2(n10969), .B1(
        i_data_bus[752]), .B2(n10988), .ZN(n10663) );
  AOI22D1BWP30P140LVT U11236 ( .A1(i_data_bus[656]), .A2(n10965), .B1(
        i_data_bus[176]), .B2(n10976), .ZN(n10662) );
  AOI22D1BWP30P140LVT U11237 ( .A1(i_data_bus[624]), .A2(n10971), .B1(
        i_data_bus[816]), .B2(n10970), .ZN(n10661) );
  AOI22D1BWP30P140LVT U11238 ( .A1(i_data_bus[336]), .A2(n10964), .B1(
        i_data_bus[848]), .B2(n10993), .ZN(n10660) );
  ND4D1BWP30P140LVT U11239 ( .A1(n10663), .A2(n10662), .A3(n10661), .A4(n10660), .ZN(n10669) );
  AOI22D1BWP30P140LVT U11240 ( .A1(i_data_bus[592]), .A2(n10981), .B1(
        i_data_bus[688]), .B2(n10977), .ZN(n10667) );
  AOI22D1BWP30P140LVT U11241 ( .A1(i_data_bus[16]), .A2(n10967), .B1(
        i_data_bus[464]), .B2(n10992), .ZN(n10666) );
  AOI22D1BWP30P140LVT U11242 ( .A1(i_data_bus[48]), .A2(n10979), .B1(
        i_data_bus[368]), .B2(n10978), .ZN(n10665) );
  AOI22D1BWP30P140LVT U11243 ( .A1(i_data_bus[272]), .A2(n10968), .B1(
        i_data_bus[240]), .B2(n10990), .ZN(n10664) );
  ND4D1BWP30P140LVT U11244 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(n10668) );
  OR4D1BWP30P140LVT U11245 ( .A1(n10671), .A2(n10670), .A3(n10669), .A4(n10668), .Z(o_data_bus[208]) );
  AOI22D1BWP30P140LVT U11246 ( .A1(i_data_bus[1009]), .A2(n10955), .B1(
        i_data_bus[913]), .B2(n10952), .ZN(n10675) );
  AOI22D1BWP30P140LVT U11247 ( .A1(i_data_bus[945]), .A2(n10954), .B1(
        i_data_bus[977]), .B2(n10953), .ZN(n10674) );
  AOI22D1BWP30P140LVT U11248 ( .A1(i_data_bus[49]), .A2(n10979), .B1(
        i_data_bus[145]), .B2(n10966), .ZN(n10673) );
  AOI22D1BWP30P140LVT U11249 ( .A1(i_data_bus[401]), .A2(n10994), .B1(
        i_data_bus[209]), .B2(n10983), .ZN(n10672) );
  ND4D1BWP30P140LVT U11250 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10672), .ZN(n10691) );
  AOI22D1BWP30P140LVT U11251 ( .A1(i_data_bus[721]), .A2(n10995), .B1(
        i_data_bus[657]), .B2(n10965), .ZN(n10679) );
  AOI22D1BWP30P140LVT U11252 ( .A1(i_data_bus[753]), .A2(n10988), .B1(
        i_data_bus[465]), .B2(n10992), .ZN(n10678) );
  AOI22D1BWP30P140LVT U11253 ( .A1(i_data_bus[273]), .A2(n10968), .B1(
        i_data_bus[369]), .B2(n10978), .ZN(n10677) );
  AOI22D1BWP30P140LVT U11254 ( .A1(i_data_bus[529]), .A2(n10957), .B1(
        i_data_bus[433]), .B2(n10969), .ZN(n10676) );
  ND4D1BWP30P140LVT U11255 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(n10690) );
  AOI22D1BWP30P140LVT U11256 ( .A1(i_data_bus[881]), .A2(n10982), .B1(
        i_data_bus[305]), .B2(n10980), .ZN(n10683) );
  AOI22D1BWP30P140LVT U11257 ( .A1(i_data_bus[241]), .A2(n10990), .B1(
        i_data_bus[817]), .B2(n10970), .ZN(n10682) );
  AOI22D1BWP30P140LVT U11258 ( .A1(i_data_bus[625]), .A2(n10971), .B1(
        i_data_bus[81]), .B2(n10959), .ZN(n10681) );
  AOI22D1BWP30P140LVT U11259 ( .A1(i_data_bus[113]), .A2(n10991), .B1(
        i_data_bus[177]), .B2(n10976), .ZN(n10680) );
  ND4D1BWP30P140LVT U11260 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(n10689) );
  AOI22D1BWP30P140LVT U11261 ( .A1(i_data_bus[689]), .A2(n10977), .B1(
        i_data_bus[785]), .B2(n10956), .ZN(n10687) );
  AOI22D1BWP30P140LVT U11262 ( .A1(i_data_bus[17]), .A2(n10967), .B1(
        i_data_bus[497]), .B2(n10989), .ZN(n10686) );
  AOI22D1BWP30P140LVT U11263 ( .A1(i_data_bus[593]), .A2(n10981), .B1(
        i_data_bus[849]), .B2(n10993), .ZN(n10685) );
  AOI22D1BWP30P140LVT U11264 ( .A1(i_data_bus[561]), .A2(n10958), .B1(
        i_data_bus[337]), .B2(n10964), .ZN(n10684) );
  ND4D1BWP30P140LVT U11265 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(n10688) );
  OR4D1BWP30P140LVT U11266 ( .A1(n10691), .A2(n10690), .A3(n10689), .A4(n10688), .Z(o_data_bus[209]) );
  AOI22D1BWP30P140LVT U11267 ( .A1(i_data_bus[978]), .A2(n10953), .B1(
        i_data_bus[914]), .B2(n10952), .ZN(n10695) );
  AOI22D1BWP30P140LVT U11268 ( .A1(i_data_bus[1010]), .A2(n10955), .B1(
        i_data_bus[946]), .B2(n10954), .ZN(n10694) );
  AOI22D1BWP30P140LVT U11269 ( .A1(i_data_bus[370]), .A2(n10978), .B1(
        i_data_bus[434]), .B2(n10969), .ZN(n10693) );
  AOI22D1BWP30P140LVT U11270 ( .A1(i_data_bus[626]), .A2(n10971), .B1(
        i_data_bus[146]), .B2(n10966), .ZN(n10692) );
  ND4D1BWP30P140LVT U11271 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(n10711) );
  AOI22D1BWP30P140LVT U11272 ( .A1(i_data_bus[882]), .A2(n10982), .B1(
        i_data_bus[690]), .B2(n10977), .ZN(n10699) );
  AOI22D1BWP30P140LVT U11273 ( .A1(i_data_bus[594]), .A2(n10981), .B1(
        i_data_bus[18]), .B2(n10967), .ZN(n10698) );
  AOI22D1BWP30P140LVT U11274 ( .A1(i_data_bus[402]), .A2(n10994), .B1(
        i_data_bus[498]), .B2(n10989), .ZN(n10697) );
  AOI22D1BWP30P140LVT U11275 ( .A1(i_data_bus[850]), .A2(n10993), .B1(
        i_data_bus[274]), .B2(n10968), .ZN(n10696) );
  ND4D1BWP30P140LVT U11276 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(n10710) );
  AOI22D1BWP30P140LVT U11277 ( .A1(i_data_bus[50]), .A2(n10979), .B1(
        i_data_bus[114]), .B2(n10991), .ZN(n10703) );
  AOI22D1BWP30P140LVT U11278 ( .A1(i_data_bus[82]), .A2(n10959), .B1(
        i_data_bus[658]), .B2(n10965), .ZN(n10702) );
  AOI22D1BWP30P140LVT U11279 ( .A1(i_data_bus[562]), .A2(n10958), .B1(
        i_data_bus[210]), .B2(n10983), .ZN(n10701) );
  AOI22D1BWP30P140LVT U11280 ( .A1(i_data_bus[178]), .A2(n10976), .B1(
        i_data_bus[754]), .B2(n10988), .ZN(n10700) );
  ND4D1BWP30P140LVT U11281 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(n10709) );
  AOI22D1BWP30P140LVT U11282 ( .A1(i_data_bus[242]), .A2(n10990), .B1(
        i_data_bus[306]), .B2(n10980), .ZN(n10707) );
  AOI22D1BWP30P140LVT U11283 ( .A1(i_data_bus[818]), .A2(n10970), .B1(
        i_data_bus[338]), .B2(n10964), .ZN(n10706) );
  AOI22D1BWP30P140LVT U11284 ( .A1(i_data_bus[530]), .A2(n10957), .B1(
        i_data_bus[722]), .B2(n10995), .ZN(n10705) );
  AOI22D1BWP30P140LVT U11285 ( .A1(i_data_bus[466]), .A2(n10992), .B1(
        i_data_bus[786]), .B2(n10956), .ZN(n10704) );
  ND4D1BWP30P140LVT U11286 ( .A1(n10707), .A2(n10706), .A3(n10705), .A4(n10704), .ZN(n10708) );
  OR4D1BWP30P140LVT U11287 ( .A1(n10711), .A2(n10710), .A3(n10709), .A4(n10708), .Z(o_data_bus[210]) );
  AOI22D1BWP30P140LVT U11288 ( .A1(i_data_bus[979]), .A2(n10953), .B1(
        i_data_bus[915]), .B2(n10952), .ZN(n10715) );
  AOI22D1BWP30P140LVT U11289 ( .A1(i_data_bus[1011]), .A2(n10955), .B1(
        i_data_bus[947]), .B2(n10954), .ZN(n10714) );
  AOI22D1BWP30P140LVT U11290 ( .A1(i_data_bus[211]), .A2(n10983), .B1(
        i_data_bus[307]), .B2(n10980), .ZN(n10713) );
  AOI22D1BWP30P140LVT U11291 ( .A1(i_data_bus[755]), .A2(n10988), .B1(
        i_data_bus[659]), .B2(n10965), .ZN(n10712) );
  ND4D1BWP30P140LVT U11292 ( .A1(n10715), .A2(n10714), .A3(n10713), .A4(n10712), .ZN(n10731) );
  AOI22D1BWP30P140LVT U11293 ( .A1(i_data_bus[531]), .A2(n10957), .B1(
        i_data_bus[19]), .B2(n10967), .ZN(n10719) );
  AOI22D1BWP30P140LVT U11294 ( .A1(i_data_bus[51]), .A2(n10979), .B1(
        i_data_bus[595]), .B2(n10981), .ZN(n10718) );
  AOI22D1BWP30P140LVT U11295 ( .A1(i_data_bus[563]), .A2(n10958), .B1(
        i_data_bus[787]), .B2(n10956), .ZN(n10717) );
  AOI22D1BWP30P140LVT U11296 ( .A1(i_data_bus[627]), .A2(n10971), .B1(
        i_data_bus[723]), .B2(n10995), .ZN(n10716) );
  ND4D1BWP30P140LVT U11297 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(n10730) );
  AOI22D1BWP30P140LVT U11298 ( .A1(i_data_bus[115]), .A2(n10991), .B1(
        i_data_bus[275]), .B2(n10968), .ZN(n10723) );
  AOI22D1BWP30P140LVT U11299 ( .A1(i_data_bus[371]), .A2(n10978), .B1(
        i_data_bus[467]), .B2(n10992), .ZN(n10722) );
  AOI22D1BWP30P140LVT U11300 ( .A1(i_data_bus[243]), .A2(n10990), .B1(
        i_data_bus[819]), .B2(n10970), .ZN(n10721) );
  AOI22D1BWP30P140LVT U11301 ( .A1(i_data_bus[339]), .A2(n10964), .B1(
        i_data_bus[435]), .B2(n10969), .ZN(n10720) );
  ND4D1BWP30P140LVT U11302 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(n10729) );
  AOI22D1BWP30P140LVT U11303 ( .A1(i_data_bus[883]), .A2(n10982), .B1(
        i_data_bus[691]), .B2(n10977), .ZN(n10727) );
  AOI22D1BWP30P140LVT U11304 ( .A1(i_data_bus[403]), .A2(n10994), .B1(
        i_data_bus[851]), .B2(n10993), .ZN(n10726) );
  AOI22D1BWP30P140LVT U11305 ( .A1(i_data_bus[83]), .A2(n10959), .B1(
        i_data_bus[147]), .B2(n10966), .ZN(n10725) );
  AOI22D1BWP30P140LVT U11306 ( .A1(i_data_bus[179]), .A2(n10976), .B1(
        i_data_bus[499]), .B2(n10989), .ZN(n10724) );
  ND4D1BWP30P140LVT U11307 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(n10728) );
  OR4D1BWP30P140LVT U11308 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .Z(o_data_bus[211]) );
  AOI22D1BWP30P140LVT U11309 ( .A1(i_data_bus[980]), .A2(n10953), .B1(
        i_data_bus[916]), .B2(n10952), .ZN(n10735) );
  AOI22D1BWP30P140LVT U11310 ( .A1(i_data_bus[1012]), .A2(n10955), .B1(
        i_data_bus[948]), .B2(n10954), .ZN(n10734) );
  AOI22D1BWP30P140LVT U11311 ( .A1(i_data_bus[788]), .A2(n10956), .B1(
        i_data_bus[372]), .B2(n10978), .ZN(n10733) );
  AOI22D1BWP30P140LVT U11312 ( .A1(i_data_bus[212]), .A2(n10983), .B1(
        i_data_bus[660]), .B2(n10965), .ZN(n10732) );
  ND4D1BWP30P140LVT U11313 ( .A1(n10735), .A2(n10734), .A3(n10733), .A4(n10732), .ZN(n10751) );
  AOI22D1BWP30P140LVT U11314 ( .A1(i_data_bus[628]), .A2(n10971), .B1(
        i_data_bus[436]), .B2(n10969), .ZN(n10739) );
  AOI22D1BWP30P140LVT U11315 ( .A1(i_data_bus[596]), .A2(n10981), .B1(
        i_data_bus[852]), .B2(n10993), .ZN(n10738) );
  AOI22D1BWP30P140LVT U11316 ( .A1(i_data_bus[532]), .A2(n10957), .B1(
        i_data_bus[884]), .B2(n10982), .ZN(n10737) );
  AOI22D1BWP30P140LVT U11317 ( .A1(i_data_bus[52]), .A2(n10979), .B1(
        i_data_bus[276]), .B2(n10968), .ZN(n10736) );
  ND4D1BWP30P140LVT U11318 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(n10750) );
  AOI22D1BWP30P140LVT U11319 ( .A1(i_data_bus[756]), .A2(n10988), .B1(
        i_data_bus[692]), .B2(n10977), .ZN(n10743) );
  AOI22D1BWP30P140LVT U11320 ( .A1(i_data_bus[20]), .A2(n10967), .B1(
        i_data_bus[820]), .B2(n10970), .ZN(n10742) );
  AOI22D1BWP30P140LVT U11321 ( .A1(i_data_bus[84]), .A2(n10959), .B1(
        i_data_bus[468]), .B2(n10992), .ZN(n10741) );
  AOI22D1BWP30P140LVT U11322 ( .A1(i_data_bus[244]), .A2(n10990), .B1(
        i_data_bus[308]), .B2(n10980), .ZN(n10740) );
  ND4D1BWP30P140LVT U11323 ( .A1(n10743), .A2(n10742), .A3(n10741), .A4(n10740), .ZN(n10749) );
  AOI22D1BWP30P140LVT U11324 ( .A1(i_data_bus[116]), .A2(n10991), .B1(
        i_data_bus[180]), .B2(n10976), .ZN(n10747) );
  AOI22D1BWP30P140LVT U11325 ( .A1(i_data_bus[724]), .A2(n10995), .B1(
        i_data_bus[500]), .B2(n10989), .ZN(n10746) );
  AOI22D1BWP30P140LVT U11326 ( .A1(i_data_bus[404]), .A2(n10994), .B1(
        i_data_bus[148]), .B2(n10966), .ZN(n10745) );
  AOI22D1BWP30P140LVT U11327 ( .A1(i_data_bus[564]), .A2(n10958), .B1(
        i_data_bus[340]), .B2(n10964), .ZN(n10744) );
  ND4D1BWP30P140LVT U11328 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(n10748) );
  OR4D1BWP30P140LVT U11329 ( .A1(n10751), .A2(n10750), .A3(n10749), .A4(n10748), .Z(o_data_bus[212]) );
  AOI22D1BWP30P140LVT U11330 ( .A1(i_data_bus[917]), .A2(n10952), .B1(
        i_data_bus[1013]), .B2(n10955), .ZN(n10755) );
  AOI22D1BWP30P140LVT U11331 ( .A1(i_data_bus[949]), .A2(n10954), .B1(
        i_data_bus[981]), .B2(n10953), .ZN(n10754) );
  AOI22D1BWP30P140LVT U11332 ( .A1(i_data_bus[501]), .A2(n10989), .B1(
        i_data_bus[373]), .B2(n10978), .ZN(n10753) );
  AOI22D1BWP30P140LVT U11333 ( .A1(i_data_bus[565]), .A2(n10958), .B1(
        i_data_bus[853]), .B2(n10993), .ZN(n10752) );
  ND4D1BWP30P140LVT U11334 ( .A1(n10755), .A2(n10754), .A3(n10753), .A4(n10752), .ZN(n10771) );
  AOI22D1BWP30P140LVT U11335 ( .A1(i_data_bus[53]), .A2(n10979), .B1(
        i_data_bus[885]), .B2(n10982), .ZN(n10759) );
  AOI22D1BWP30P140LVT U11336 ( .A1(i_data_bus[629]), .A2(n10971), .B1(
        i_data_bus[533]), .B2(n10957), .ZN(n10758) );
  AOI22D1BWP30P140LVT U11337 ( .A1(i_data_bus[597]), .A2(n10981), .B1(
        i_data_bus[277]), .B2(n10968), .ZN(n10757) );
  AOI22D1BWP30P140LVT U11338 ( .A1(i_data_bus[341]), .A2(n10964), .B1(
        i_data_bus[309]), .B2(n10980), .ZN(n10756) );
  ND4D1BWP30P140LVT U11339 ( .A1(n10759), .A2(n10758), .A3(n10757), .A4(n10756), .ZN(n10770) );
  AOI22D1BWP30P140LVT U11340 ( .A1(i_data_bus[213]), .A2(n10983), .B1(
        i_data_bus[469]), .B2(n10992), .ZN(n10763) );
  AOI22D1BWP30P140LVT U11341 ( .A1(i_data_bus[789]), .A2(n10956), .B1(
        i_data_bus[149]), .B2(n10966), .ZN(n10762) );
  AOI22D1BWP30P140LVT U11342 ( .A1(i_data_bus[85]), .A2(n10959), .B1(
        i_data_bus[661]), .B2(n10965), .ZN(n10761) );
  AOI22D1BWP30P140LVT U11343 ( .A1(i_data_bus[21]), .A2(n10967), .B1(
        i_data_bus[725]), .B2(n10995), .ZN(n10760) );
  ND4D1BWP30P140LVT U11344 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10760), .ZN(n10769) );
  AOI22D1BWP30P140LVT U11345 ( .A1(i_data_bus[757]), .A2(n10988), .B1(
        i_data_bus[821]), .B2(n10970), .ZN(n10767) );
  AOI22D1BWP30P140LVT U11346 ( .A1(i_data_bus[245]), .A2(n10990), .B1(
        i_data_bus[405]), .B2(n10994), .ZN(n10766) );
  AOI22D1BWP30P140LVT U11347 ( .A1(i_data_bus[117]), .A2(n10991), .B1(
        i_data_bus[437]), .B2(n10969), .ZN(n10765) );
  AOI22D1BWP30P140LVT U11348 ( .A1(i_data_bus[181]), .A2(n10976), .B1(
        i_data_bus[693]), .B2(n10977), .ZN(n10764) );
  ND4D1BWP30P140LVT U11349 ( .A1(n10767), .A2(n10766), .A3(n10765), .A4(n10764), .ZN(n10768) );
  OR4D1BWP30P140LVT U11350 ( .A1(n10771), .A2(n10770), .A3(n10769), .A4(n10768), .Z(o_data_bus[213]) );
  AOI22D1BWP30P140LVT U11351 ( .A1(i_data_bus[1014]), .A2(n10955), .B1(
        i_data_bus[918]), .B2(n10952), .ZN(n10775) );
  AOI22D1BWP30P140LVT U11352 ( .A1(i_data_bus[950]), .A2(n10954), .B1(
        i_data_bus[982]), .B2(n10953), .ZN(n10774) );
  AOI22D1BWP30P140LVT U11353 ( .A1(i_data_bus[822]), .A2(n10970), .B1(
        i_data_bus[246]), .B2(n10990), .ZN(n10773) );
  AOI22D1BWP30P140LVT U11354 ( .A1(i_data_bus[374]), .A2(n10978), .B1(
        i_data_bus[150]), .B2(n10966), .ZN(n10772) );
  ND4D1BWP30P140LVT U11355 ( .A1(n10775), .A2(n10774), .A3(n10773), .A4(n10772), .ZN(n10791) );
  AOI22D1BWP30P140LVT U11356 ( .A1(i_data_bus[406]), .A2(n10994), .B1(
        i_data_bus[662]), .B2(n10965), .ZN(n10779) );
  AOI22D1BWP30P140LVT U11357 ( .A1(i_data_bus[630]), .A2(n10971), .B1(
        i_data_bus[214]), .B2(n10983), .ZN(n10778) );
  AOI22D1BWP30P140LVT U11358 ( .A1(i_data_bus[118]), .A2(n10991), .B1(
        i_data_bus[310]), .B2(n10980), .ZN(n10777) );
  AOI22D1BWP30P140LVT U11359 ( .A1(i_data_bus[598]), .A2(n10981), .B1(
        i_data_bus[854]), .B2(n10993), .ZN(n10776) );
  ND4D1BWP30P140LVT U11360 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(n10790) );
  AOI22D1BWP30P140LVT U11361 ( .A1(i_data_bus[54]), .A2(n10979), .B1(
        i_data_bus[566]), .B2(n10958), .ZN(n10783) );
  AOI22D1BWP30P140LVT U11362 ( .A1(i_data_bus[502]), .A2(n10989), .B1(
        i_data_bus[470]), .B2(n10992), .ZN(n10782) );
  AOI22D1BWP30P140LVT U11363 ( .A1(i_data_bus[726]), .A2(n10995), .B1(
        i_data_bus[278]), .B2(n10968), .ZN(n10781) );
  AOI22D1BWP30P140LVT U11364 ( .A1(i_data_bus[22]), .A2(n10967), .B1(
        i_data_bus[342]), .B2(n10964), .ZN(n10780) );
  ND4D1BWP30P140LVT U11365 ( .A1(n10783), .A2(n10782), .A3(n10781), .A4(n10780), .ZN(n10789) );
  AOI22D1BWP30P140LVT U11366 ( .A1(i_data_bus[86]), .A2(n10959), .B1(
        i_data_bus[886]), .B2(n10982), .ZN(n10787) );
  AOI22D1BWP30P140LVT U11367 ( .A1(i_data_bus[534]), .A2(n10957), .B1(
        i_data_bus[438]), .B2(n10969), .ZN(n10786) );
  AOI22D1BWP30P140LVT U11368 ( .A1(i_data_bus[790]), .A2(n10956), .B1(
        i_data_bus[182]), .B2(n10976), .ZN(n10785) );
  AOI22D1BWP30P140LVT U11369 ( .A1(i_data_bus[694]), .A2(n10977), .B1(
        i_data_bus[758]), .B2(n10988), .ZN(n10784) );
  ND4D1BWP30P140LVT U11370 ( .A1(n10787), .A2(n10786), .A3(n10785), .A4(n10784), .ZN(n10788) );
  OR4D1BWP30P140LVT U11371 ( .A1(n10791), .A2(n10790), .A3(n10789), .A4(n10788), .Z(o_data_bus[214]) );
  AOI22D1BWP30P140LVT U11372 ( .A1(i_data_bus[951]), .A2(n10954), .B1(
        i_data_bus[919]), .B2(n10952), .ZN(n10795) );
  AOI22D1BWP30P140LVT U11373 ( .A1(i_data_bus[1015]), .A2(n10955), .B1(
        i_data_bus[983]), .B2(n10953), .ZN(n10794) );
  AOI22D1BWP30P140LVT U11374 ( .A1(i_data_bus[727]), .A2(n10995), .B1(
        i_data_bus[823]), .B2(n10970), .ZN(n10793) );
  AOI22D1BWP30P140LVT U11375 ( .A1(i_data_bus[535]), .A2(n10957), .B1(
        i_data_bus[151]), .B2(n10966), .ZN(n10792) );
  ND4D1BWP30P140LVT U11376 ( .A1(n10795), .A2(n10794), .A3(n10793), .A4(n10792), .ZN(n10811) );
  AOI22D1BWP30P140LVT U11377 ( .A1(i_data_bus[503]), .A2(n10989), .B1(
        i_data_bus[407]), .B2(n10994), .ZN(n10799) );
  AOI22D1BWP30P140LVT U11378 ( .A1(i_data_bus[119]), .A2(n10991), .B1(
        i_data_bus[759]), .B2(n10988), .ZN(n10798) );
  AOI22D1BWP30P140LVT U11379 ( .A1(i_data_bus[695]), .A2(n10977), .B1(
        i_data_bus[663]), .B2(n10965), .ZN(n10797) );
  AOI22D1BWP30P140LVT U11380 ( .A1(i_data_bus[471]), .A2(n10992), .B1(
        i_data_bus[855]), .B2(n10993), .ZN(n10796) );
  ND4D1BWP30P140LVT U11381 ( .A1(n10799), .A2(n10798), .A3(n10797), .A4(n10796), .ZN(n10810) );
  AOI22D1BWP30P140LVT U11382 ( .A1(i_data_bus[599]), .A2(n10981), .B1(
        i_data_bus[887]), .B2(n10982), .ZN(n10803) );
  AOI22D1BWP30P140LVT U11383 ( .A1(i_data_bus[311]), .A2(n10980), .B1(
        i_data_bus[343]), .B2(n10964), .ZN(n10802) );
  AOI22D1BWP30P140LVT U11384 ( .A1(i_data_bus[247]), .A2(n10990), .B1(
        i_data_bus[791]), .B2(n10956), .ZN(n10801) );
  AOI22D1BWP30P140LVT U11385 ( .A1(i_data_bus[23]), .A2(n10967), .B1(
        i_data_bus[567]), .B2(n10958), .ZN(n10800) );
  ND4D1BWP30P140LVT U11386 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(n10809) );
  AOI22D1BWP30P140LVT U11387 ( .A1(i_data_bus[87]), .A2(n10959), .B1(
        i_data_bus[183]), .B2(n10976), .ZN(n10807) );
  AOI22D1BWP30P140LVT U11388 ( .A1(i_data_bus[55]), .A2(n10979), .B1(
        i_data_bus[375]), .B2(n10978), .ZN(n10806) );
  AOI22D1BWP30P140LVT U11389 ( .A1(i_data_bus[279]), .A2(n10968), .B1(
        i_data_bus[215]), .B2(n10983), .ZN(n10805) );
  AOI22D1BWP30P140LVT U11390 ( .A1(i_data_bus[631]), .A2(n10971), .B1(
        i_data_bus[439]), .B2(n10969), .ZN(n10804) );
  ND4D1BWP30P140LVT U11391 ( .A1(n10807), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(n10808) );
  OR4D1BWP30P140LVT U11392 ( .A1(n10811), .A2(n10810), .A3(n10809), .A4(n10808), .Z(o_data_bus[215]) );
  AOI22D1BWP30P140LVT U11393 ( .A1(i_data_bus[952]), .A2(n10954), .B1(
        i_data_bus[920]), .B2(n10952), .ZN(n10815) );
  AOI22D1BWP30P140LVT U11394 ( .A1(i_data_bus[984]), .A2(n10953), .B1(
        i_data_bus[1016]), .B2(n10955), .ZN(n10814) );
  AOI22D1BWP30P140LVT U11395 ( .A1(i_data_bus[600]), .A2(n10981), .B1(
        i_data_bus[472]), .B2(n10992), .ZN(n10813) );
  AOI22D1BWP30P140LVT U11396 ( .A1(i_data_bus[568]), .A2(n10958), .B1(
        i_data_bus[504]), .B2(n10989), .ZN(n10812) );
  ND4D1BWP30P140LVT U11397 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(n10831) );
  AOI22D1BWP30P140LVT U11398 ( .A1(i_data_bus[440]), .A2(n10969), .B1(
        i_data_bus[728]), .B2(n10995), .ZN(n10819) );
  AOI22D1BWP30P140LVT U11399 ( .A1(i_data_bus[632]), .A2(n10971), .B1(
        i_data_bus[88]), .B2(n10959), .ZN(n10818) );
  AOI22D1BWP30P140LVT U11400 ( .A1(i_data_bus[408]), .A2(n10994), .B1(
        i_data_bus[184]), .B2(n10976), .ZN(n10817) );
  AOI22D1BWP30P140LVT U11401 ( .A1(i_data_bus[856]), .A2(n10993), .B1(
        i_data_bus[824]), .B2(n10970), .ZN(n10816) );
  ND4D1BWP30P140LVT U11402 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(n10830) );
  AOI22D1BWP30P140LVT U11403 ( .A1(i_data_bus[120]), .A2(n10991), .B1(
        i_data_bus[280]), .B2(n10968), .ZN(n10823) );
  AOI22D1BWP30P140LVT U11404 ( .A1(i_data_bus[24]), .A2(n10967), .B1(
        i_data_bus[376]), .B2(n10978), .ZN(n10822) );
  AOI22D1BWP30P140LVT U11405 ( .A1(i_data_bus[536]), .A2(n10957), .B1(
        i_data_bus[792]), .B2(n10956), .ZN(n10821) );
  AOI22D1BWP30P140LVT U11406 ( .A1(i_data_bus[248]), .A2(n10990), .B1(
        i_data_bus[152]), .B2(n10966), .ZN(n10820) );
  ND4D1BWP30P140LVT U11407 ( .A1(n10823), .A2(n10822), .A3(n10821), .A4(n10820), .ZN(n10829) );
  AOI22D1BWP30P140LVT U11408 ( .A1(i_data_bus[344]), .A2(n10964), .B1(
        i_data_bus[312]), .B2(n10980), .ZN(n10827) );
  AOI22D1BWP30P140LVT U11409 ( .A1(i_data_bus[56]), .A2(n10979), .B1(
        i_data_bus[696]), .B2(n10977), .ZN(n10826) );
  AOI22D1BWP30P140LVT U11410 ( .A1(i_data_bus[888]), .A2(n10982), .B1(
        i_data_bus[760]), .B2(n10988), .ZN(n10825) );
  AOI22D1BWP30P140LVT U11411 ( .A1(i_data_bus[664]), .A2(n10965), .B1(
        i_data_bus[216]), .B2(n10983), .ZN(n10824) );
  ND4D1BWP30P140LVT U11412 ( .A1(n10827), .A2(n10826), .A3(n10825), .A4(n10824), .ZN(n10828) );
  OR4D1BWP30P140LVT U11413 ( .A1(n10831), .A2(n10830), .A3(n10829), .A4(n10828), .Z(o_data_bus[216]) );
  AOI22D1BWP30P140LVT U11414 ( .A1(i_data_bus[1017]), .A2(n10955), .B1(
        i_data_bus[921]), .B2(n10952), .ZN(n10835) );
  AOI22D1BWP30P140LVT U11415 ( .A1(i_data_bus[985]), .A2(n10953), .B1(
        i_data_bus[953]), .B2(n10954), .ZN(n10834) );
  AOI22D1BWP30P140LVT U11416 ( .A1(i_data_bus[665]), .A2(n10965), .B1(
        i_data_bus[153]), .B2(n10966), .ZN(n10833) );
  AOI22D1BWP30P140LVT U11417 ( .A1(i_data_bus[601]), .A2(n10981), .B1(
        i_data_bus[281]), .B2(n10968), .ZN(n10832) );
  ND4D1BWP30P140LVT U11418 ( .A1(n10835), .A2(n10834), .A3(n10833), .A4(n10832), .ZN(n10851) );
  AOI22D1BWP30P140LVT U11419 ( .A1(i_data_bus[761]), .A2(n10988), .B1(
        i_data_bus[505]), .B2(n10989), .ZN(n10839) );
  AOI22D1BWP30P140LVT U11420 ( .A1(i_data_bus[633]), .A2(n10971), .B1(
        i_data_bus[345]), .B2(n10964), .ZN(n10838) );
  AOI22D1BWP30P140LVT U11421 ( .A1(i_data_bus[729]), .A2(n10995), .B1(
        i_data_bus[441]), .B2(n10969), .ZN(n10837) );
  AOI22D1BWP30P140LVT U11422 ( .A1(i_data_bus[537]), .A2(n10957), .B1(
        i_data_bus[857]), .B2(n10993), .ZN(n10836) );
  ND4D1BWP30P140LVT U11423 ( .A1(n10839), .A2(n10838), .A3(n10837), .A4(n10836), .ZN(n10850) );
  AOI22D1BWP30P140LVT U11424 ( .A1(i_data_bus[89]), .A2(n10959), .B1(
        i_data_bus[409]), .B2(n10994), .ZN(n10843) );
  AOI22D1BWP30P140LVT U11425 ( .A1(i_data_bus[25]), .A2(n10967), .B1(
        i_data_bus[313]), .B2(n10980), .ZN(n10842) );
  AOI22D1BWP30P140LVT U11426 ( .A1(i_data_bus[473]), .A2(n10992), .B1(
        i_data_bus[249]), .B2(n10990), .ZN(n10841) );
  AOI22D1BWP30P140LVT U11427 ( .A1(i_data_bus[793]), .A2(n10956), .B1(
        i_data_bus[377]), .B2(n10978), .ZN(n10840) );
  ND4D1BWP30P140LVT U11428 ( .A1(n10843), .A2(n10842), .A3(n10841), .A4(n10840), .ZN(n10849) );
  AOI22D1BWP30P140LVT U11429 ( .A1(i_data_bus[57]), .A2(n10979), .B1(
        i_data_bus[185]), .B2(n10976), .ZN(n10847) );
  AOI22D1BWP30P140LVT U11430 ( .A1(i_data_bus[697]), .A2(n10977), .B1(
        i_data_bus[217]), .B2(n10983), .ZN(n10846) );
  AOI22D1BWP30P140LVT U11431 ( .A1(i_data_bus[825]), .A2(n10970), .B1(
        i_data_bus[889]), .B2(n10982), .ZN(n10845) );
  AOI22D1BWP30P140LVT U11432 ( .A1(i_data_bus[569]), .A2(n10958), .B1(
        i_data_bus[121]), .B2(n10991), .ZN(n10844) );
  ND4D1BWP30P140LVT U11433 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(n10848) );
  OR4D1BWP30P140LVT U11434 ( .A1(n10851), .A2(n10850), .A3(n10849), .A4(n10848), .Z(o_data_bus[217]) );
  AOI22D1BWP30P140LVT U11435 ( .A1(i_data_bus[954]), .A2(n10954), .B1(
        i_data_bus[986]), .B2(n10953), .ZN(n10855) );
  AOI22D1BWP30P140LVT U11436 ( .A1(i_data_bus[1018]), .A2(n10955), .B1(
        i_data_bus[922]), .B2(n10952), .ZN(n10854) );
  AOI22D1BWP30P140LVT U11437 ( .A1(i_data_bus[538]), .A2(n10957), .B1(
        i_data_bus[666]), .B2(n10965), .ZN(n10853) );
  AOI22D1BWP30P140LVT U11438 ( .A1(i_data_bus[698]), .A2(n10977), .B1(
        i_data_bus[378]), .B2(n10978), .ZN(n10852) );
  ND4D1BWP30P140LVT U11439 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(n10871) );
  AOI22D1BWP30P140LVT U11440 ( .A1(i_data_bus[602]), .A2(n10981), .B1(
        i_data_bus[730]), .B2(n10995), .ZN(n10859) );
  AOI22D1BWP30P140LVT U11441 ( .A1(i_data_bus[570]), .A2(n10958), .B1(
        i_data_bus[506]), .B2(n10989), .ZN(n10858) );
  AOI22D1BWP30P140LVT U11442 ( .A1(i_data_bus[218]), .A2(n10983), .B1(
        i_data_bus[346]), .B2(n10964), .ZN(n10857) );
  AOI22D1BWP30P140LVT U11443 ( .A1(i_data_bus[442]), .A2(n10969), .B1(
        i_data_bus[762]), .B2(n10988), .ZN(n10856) );
  ND4D1BWP30P140LVT U11444 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(n10870) );
  AOI22D1BWP30P140LVT U11445 ( .A1(i_data_bus[634]), .A2(n10971), .B1(
        i_data_bus[282]), .B2(n10968), .ZN(n10863) );
  AOI22D1BWP30P140LVT U11446 ( .A1(i_data_bus[58]), .A2(n10979), .B1(
        i_data_bus[314]), .B2(n10980), .ZN(n10862) );
  AOI22D1BWP30P140LVT U11447 ( .A1(i_data_bus[26]), .A2(n10967), .B1(
        i_data_bus[794]), .B2(n10956), .ZN(n10861) );
  AOI22D1BWP30P140LVT U11448 ( .A1(i_data_bus[826]), .A2(n10970), .B1(
        i_data_bus[474]), .B2(n10992), .ZN(n10860) );
  ND4D1BWP30P140LVT U11449 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(n10869) );
  AOI22D1BWP30P140LVT U11450 ( .A1(i_data_bus[858]), .A2(n10993), .B1(
        i_data_bus[250]), .B2(n10990), .ZN(n10867) );
  AOI22D1BWP30P140LVT U11451 ( .A1(i_data_bus[90]), .A2(n10959), .B1(
        i_data_bus[186]), .B2(n10976), .ZN(n10866) );
  AOI22D1BWP30P140LVT U11452 ( .A1(i_data_bus[890]), .A2(n10982), .B1(
        i_data_bus[154]), .B2(n10966), .ZN(n10865) );
  AOI22D1BWP30P140LVT U11453 ( .A1(i_data_bus[122]), .A2(n10991), .B1(
        i_data_bus[410]), .B2(n10994), .ZN(n10864) );
  ND4D1BWP30P140LVT U11454 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(n10868) );
  OR4D1BWP30P140LVT U11455 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .Z(o_data_bus[218]) );
  AOI22D1BWP30P140LVT U11456 ( .A1(i_data_bus[987]), .A2(n10953), .B1(
        i_data_bus[923]), .B2(n10952), .ZN(n10875) );
  AOI22D1BWP30P140LVT U11457 ( .A1(i_data_bus[1019]), .A2(n10955), .B1(
        i_data_bus[955]), .B2(n10954), .ZN(n10874) );
  AOI22D1BWP30P140LVT U11458 ( .A1(i_data_bus[91]), .A2(n10959), .B1(
        i_data_bus[891]), .B2(n10982), .ZN(n10873) );
  AOI22D1BWP30P140LVT U11459 ( .A1(i_data_bus[539]), .A2(n10957), .B1(
        i_data_bus[27]), .B2(n10967), .ZN(n10872) );
  ND4D1BWP30P140LVT U11460 ( .A1(n10875), .A2(n10874), .A3(n10873), .A4(n10872), .ZN(n10891) );
  AOI22D1BWP30P140LVT U11461 ( .A1(i_data_bus[123]), .A2(n10991), .B1(
        i_data_bus[251]), .B2(n10990), .ZN(n10879) );
  AOI22D1BWP30P140LVT U11462 ( .A1(i_data_bus[603]), .A2(n10981), .B1(
        i_data_bus[219]), .B2(n10983), .ZN(n10878) );
  AOI22D1BWP30P140LVT U11463 ( .A1(i_data_bus[763]), .A2(n10988), .B1(
        i_data_bus[187]), .B2(n10976), .ZN(n10877) );
  AOI22D1BWP30P140LVT U11464 ( .A1(i_data_bus[571]), .A2(n10958), .B1(
        i_data_bus[635]), .B2(n10971), .ZN(n10876) );
  ND4D1BWP30P140LVT U11465 ( .A1(n10879), .A2(n10878), .A3(n10877), .A4(n10876), .ZN(n10890) );
  AOI22D1BWP30P140LVT U11466 ( .A1(i_data_bus[443]), .A2(n10969), .B1(
        i_data_bus[315]), .B2(n10980), .ZN(n10883) );
  AOI22D1BWP30P140LVT U11467 ( .A1(i_data_bus[59]), .A2(n10979), .B1(
        i_data_bus[379]), .B2(n10978), .ZN(n10882) );
  AOI22D1BWP30P140LVT U11468 ( .A1(i_data_bus[411]), .A2(n10994), .B1(
        i_data_bus[795]), .B2(n10956), .ZN(n10881) );
  AOI22D1BWP30P140LVT U11469 ( .A1(i_data_bus[155]), .A2(n10966), .B1(
        i_data_bus[667]), .B2(n10965), .ZN(n10880) );
  ND4D1BWP30P140LVT U11470 ( .A1(n10883), .A2(n10882), .A3(n10881), .A4(n10880), .ZN(n10889) );
  AOI22D1BWP30P140LVT U11471 ( .A1(i_data_bus[731]), .A2(n10995), .B1(
        i_data_bus[859]), .B2(n10993), .ZN(n10887) );
  AOI22D1BWP30P140LVT U11472 ( .A1(i_data_bus[283]), .A2(n10968), .B1(
        i_data_bus[475]), .B2(n10992), .ZN(n10886) );
  AOI22D1BWP30P140LVT U11473 ( .A1(i_data_bus[827]), .A2(n10970), .B1(
        i_data_bus[699]), .B2(n10977), .ZN(n10885) );
  AOI22D1BWP30P140LVT U11474 ( .A1(i_data_bus[507]), .A2(n10989), .B1(
        i_data_bus[347]), .B2(n10964), .ZN(n10884) );
  ND4D1BWP30P140LVT U11475 ( .A1(n10887), .A2(n10886), .A3(n10885), .A4(n10884), .ZN(n10888) );
  OR4D1BWP30P140LVT U11476 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .Z(o_data_bus[219]) );
  AOI22D1BWP30P140LVT U11477 ( .A1(i_data_bus[988]), .A2(n10953), .B1(
        i_data_bus[956]), .B2(n10954), .ZN(n10895) );
  AOI22D1BWP30P140LVT U11478 ( .A1(i_data_bus[924]), .A2(n10952), .B1(
        i_data_bus[1020]), .B2(n10955), .ZN(n10894) );
  AOI22D1BWP30P140LVT U11479 ( .A1(i_data_bus[764]), .A2(n10988), .B1(
        i_data_bus[316]), .B2(n10980), .ZN(n10893) );
  AOI22D1BWP30P140LVT U11480 ( .A1(i_data_bus[188]), .A2(n10976), .B1(
        i_data_bus[860]), .B2(n10993), .ZN(n10892) );
  ND4D1BWP30P140LVT U11481 ( .A1(n10895), .A2(n10894), .A3(n10893), .A4(n10892), .ZN(n10911) );
  AOI22D1BWP30P140LVT U11482 ( .A1(i_data_bus[348]), .A2(n10964), .B1(
        i_data_bus[796]), .B2(n10956), .ZN(n10899) );
  AOI22D1BWP30P140LVT U11483 ( .A1(i_data_bus[28]), .A2(n10967), .B1(
        i_data_bus[444]), .B2(n10969), .ZN(n10898) );
  AOI22D1BWP30P140LVT U11484 ( .A1(i_data_bus[636]), .A2(n10971), .B1(
        i_data_bus[572]), .B2(n10958), .ZN(n10897) );
  AOI22D1BWP30P140LVT U11485 ( .A1(i_data_bus[604]), .A2(n10981), .B1(
        i_data_bus[380]), .B2(n10978), .ZN(n10896) );
  ND4D1BWP30P140LVT U11486 ( .A1(n10899), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(n10910) );
  AOI22D1BWP30P140LVT U11487 ( .A1(i_data_bus[732]), .A2(n10995), .B1(
        i_data_bus[412]), .B2(n10994), .ZN(n10903) );
  AOI22D1BWP30P140LVT U11488 ( .A1(i_data_bus[124]), .A2(n10991), .B1(
        i_data_bus[284]), .B2(n10968), .ZN(n10902) );
  AOI22D1BWP30P140LVT U11489 ( .A1(i_data_bus[252]), .A2(n10990), .B1(
        i_data_bus[700]), .B2(n10977), .ZN(n10901) );
  AOI22D1BWP30P140LVT U11490 ( .A1(i_data_bus[60]), .A2(n10979), .B1(
        i_data_bus[892]), .B2(n10982), .ZN(n10900) );
  ND4D1BWP30P140LVT U11491 ( .A1(n10903), .A2(n10902), .A3(n10901), .A4(n10900), .ZN(n10909) );
  AOI22D1BWP30P140LVT U11492 ( .A1(i_data_bus[828]), .A2(n10970), .B1(
        i_data_bus[156]), .B2(n10966), .ZN(n10907) );
  AOI22D1BWP30P140LVT U11493 ( .A1(i_data_bus[540]), .A2(n10957), .B1(
        i_data_bus[92]), .B2(n10959), .ZN(n10906) );
  AOI22D1BWP30P140LVT U11494 ( .A1(i_data_bus[220]), .A2(n10983), .B1(
        i_data_bus[476]), .B2(n10992), .ZN(n10905) );
  AOI22D1BWP30P140LVT U11495 ( .A1(i_data_bus[508]), .A2(n10989), .B1(
        i_data_bus[668]), .B2(n10965), .ZN(n10904) );
  ND4D1BWP30P140LVT U11496 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(n10908) );
  OR4D1BWP30P140LVT U11497 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .Z(o_data_bus[220]) );
  AOI22D1BWP30P140LVT U11498 ( .A1(i_data_bus[957]), .A2(n10954), .B1(
        i_data_bus[989]), .B2(n10953), .ZN(n10915) );
  AOI22D1BWP30P140LVT U11499 ( .A1(i_data_bus[925]), .A2(n10952), .B1(
        i_data_bus[1021]), .B2(n10955), .ZN(n10914) );
  AOI22D1BWP30P140LVT U11500 ( .A1(i_data_bus[93]), .A2(n10959), .B1(
        i_data_bus[893]), .B2(n10982), .ZN(n10913) );
  AOI22D1BWP30P140LVT U11501 ( .A1(i_data_bus[797]), .A2(n10956), .B1(
        i_data_bus[381]), .B2(n10978), .ZN(n10912) );
  ND4D1BWP30P140LVT U11502 ( .A1(n10915), .A2(n10914), .A3(n10913), .A4(n10912), .ZN(n10931) );
  AOI22D1BWP30P140LVT U11503 ( .A1(i_data_bus[445]), .A2(n10969), .B1(
        i_data_bus[189]), .B2(n10976), .ZN(n10919) );
  AOI22D1BWP30P140LVT U11504 ( .A1(i_data_bus[637]), .A2(n10971), .B1(
        i_data_bus[669]), .B2(n10965), .ZN(n10918) );
  AOI22D1BWP30P140LVT U11505 ( .A1(i_data_bus[701]), .A2(n10977), .B1(
        i_data_bus[509]), .B2(n10989), .ZN(n10917) );
  AOI22D1BWP30P140LVT U11506 ( .A1(i_data_bus[573]), .A2(n10958), .B1(
        i_data_bus[829]), .B2(n10970), .ZN(n10916) );
  ND4D1BWP30P140LVT U11507 ( .A1(n10919), .A2(n10918), .A3(n10917), .A4(n10916), .ZN(n10930) );
  AOI22D1BWP30P140LVT U11508 ( .A1(i_data_bus[157]), .A2(n10966), .B1(
        i_data_bus[349]), .B2(n10964), .ZN(n10923) );
  AOI22D1BWP30P140LVT U11509 ( .A1(i_data_bus[61]), .A2(n10979), .B1(
        i_data_bus[317]), .B2(n10980), .ZN(n10922) );
  AOI22D1BWP30P140LVT U11510 ( .A1(i_data_bus[765]), .A2(n10988), .B1(
        i_data_bus[733]), .B2(n10995), .ZN(n10921) );
  AOI22D1BWP30P140LVT U11511 ( .A1(i_data_bus[29]), .A2(n10967), .B1(
        i_data_bus[477]), .B2(n10992), .ZN(n10920) );
  ND4D1BWP30P140LVT U11512 ( .A1(n10923), .A2(n10922), .A3(n10921), .A4(n10920), .ZN(n10929) );
  AOI22D1BWP30P140LVT U11513 ( .A1(i_data_bus[413]), .A2(n10994), .B1(
        i_data_bus[253]), .B2(n10990), .ZN(n10927) );
  AOI22D1BWP30P140LVT U11514 ( .A1(i_data_bus[605]), .A2(n10981), .B1(
        i_data_bus[221]), .B2(n10983), .ZN(n10926) );
  AOI22D1BWP30P140LVT U11515 ( .A1(i_data_bus[541]), .A2(n10957), .B1(
        i_data_bus[285]), .B2(n10968), .ZN(n10925) );
  AOI22D1BWP30P140LVT U11516 ( .A1(i_data_bus[125]), .A2(n10991), .B1(
        i_data_bus[861]), .B2(n10993), .ZN(n10924) );
  ND4D1BWP30P140LVT U11517 ( .A1(n10927), .A2(n10926), .A3(n10925), .A4(n10924), .ZN(n10928) );
  OR4D1BWP30P140LVT U11518 ( .A1(n10931), .A2(n10930), .A3(n10929), .A4(n10928), .Z(o_data_bus[221]) );
  AOI22D1BWP30P140LVT U11519 ( .A1(i_data_bus[958]), .A2(n10954), .B1(
        i_data_bus[990]), .B2(n10953), .ZN(n10935) );
  AOI22D1BWP30P140LVT U11520 ( .A1(i_data_bus[926]), .A2(n10952), .B1(
        i_data_bus[1022]), .B2(n10955), .ZN(n10934) );
  AOI22D1BWP30P140LVT U11521 ( .A1(i_data_bus[574]), .A2(n10958), .B1(
        i_data_bus[222]), .B2(n10983), .ZN(n10933) );
  AOI22D1BWP30P140LVT U11522 ( .A1(i_data_bus[542]), .A2(n10957), .B1(
        i_data_bus[318]), .B2(n10980), .ZN(n10932) );
  ND4D1BWP30P140LVT U11523 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10932), .ZN(n10951) );
  AOI22D1BWP30P140LVT U11524 ( .A1(i_data_bus[62]), .A2(n10979), .B1(
        i_data_bus[350]), .B2(n10964), .ZN(n10939) );
  AOI22D1BWP30P140LVT U11525 ( .A1(i_data_bus[446]), .A2(n10969), .B1(
        i_data_bus[510]), .B2(n10989), .ZN(n10938) );
  AOI22D1BWP30P140LVT U11526 ( .A1(i_data_bus[830]), .A2(n10970), .B1(
        i_data_bus[414]), .B2(n10994), .ZN(n10937) );
  AOI22D1BWP30P140LVT U11527 ( .A1(i_data_bus[286]), .A2(n10968), .B1(
        i_data_bus[702]), .B2(n10977), .ZN(n10936) );
  ND4D1BWP30P140LVT U11528 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(n10950) );
  AOI22D1BWP30P140LVT U11529 ( .A1(i_data_bus[126]), .A2(n10991), .B1(
        i_data_bus[158]), .B2(n10966), .ZN(n10943) );
  AOI22D1BWP30P140LVT U11530 ( .A1(i_data_bus[254]), .A2(n10990), .B1(
        i_data_bus[478]), .B2(n10992), .ZN(n10942) );
  AOI22D1BWP30P140LVT U11531 ( .A1(i_data_bus[670]), .A2(n10965), .B1(
        i_data_bus[734]), .B2(n10995), .ZN(n10941) );
  AOI22D1BWP30P140LVT U11532 ( .A1(i_data_bus[94]), .A2(n10959), .B1(
        i_data_bus[862]), .B2(n10993), .ZN(n10940) );
  ND4D1BWP30P140LVT U11533 ( .A1(n10943), .A2(n10942), .A3(n10941), .A4(n10940), .ZN(n10949) );
  AOI22D1BWP30P140LVT U11534 ( .A1(i_data_bus[798]), .A2(n10956), .B1(
        i_data_bus[382]), .B2(n10978), .ZN(n10947) );
  AOI22D1BWP30P140LVT U11535 ( .A1(i_data_bus[190]), .A2(n10976), .B1(
        i_data_bus[766]), .B2(n10988), .ZN(n10946) );
  AOI22D1BWP30P140LVT U11536 ( .A1(i_data_bus[30]), .A2(n10967), .B1(
        i_data_bus[606]), .B2(n10981), .ZN(n10945) );
  AOI22D1BWP30P140LVT U11537 ( .A1(i_data_bus[638]), .A2(n10971), .B1(
        i_data_bus[894]), .B2(n10982), .ZN(n10944) );
  ND4D1BWP30P140LVT U11538 ( .A1(n10947), .A2(n10946), .A3(n10945), .A4(n10944), .ZN(n10948) );
  OR4D1BWP30P140LVT U11539 ( .A1(n10951), .A2(n10950), .A3(n10949), .A4(n10948), .Z(o_data_bus[222]) );
  AOI22D1BWP30P140LVT U11540 ( .A1(i_data_bus[991]), .A2(n10953), .B1(
        i_data_bus[927]), .B2(n10952), .ZN(n10963) );
  AOI22D1BWP30P140LVT U11541 ( .A1(i_data_bus[1023]), .A2(n10955), .B1(
        i_data_bus[959]), .B2(n10954), .ZN(n10962) );
  AOI22D1BWP30P140LVT U11542 ( .A1(i_data_bus[543]), .A2(n10957), .B1(
        i_data_bus[799]), .B2(n10956), .ZN(n10961) );
  AOI22D1BWP30P140LVT U11543 ( .A1(i_data_bus[95]), .A2(n10959), .B1(
        i_data_bus[575]), .B2(n10958), .ZN(n10960) );
  ND4D1BWP30P140LVT U11544 ( .A1(n10963), .A2(n10962), .A3(n10961), .A4(n10960), .ZN(n11003) );
  AOI22D1BWP30P140LVT U11545 ( .A1(i_data_bus[671]), .A2(n10965), .B1(
        i_data_bus[351]), .B2(n10964), .ZN(n10975) );
  AOI22D1BWP30P140LVT U11546 ( .A1(i_data_bus[31]), .A2(n10967), .B1(
        i_data_bus[159]), .B2(n10966), .ZN(n10974) );
  AOI22D1BWP30P140LVT U11547 ( .A1(i_data_bus[447]), .A2(n10969), .B1(
        i_data_bus[287]), .B2(n10968), .ZN(n10973) );
  AOI22D1BWP30P140LVT U11548 ( .A1(i_data_bus[639]), .A2(n10971), .B1(
        i_data_bus[831]), .B2(n10970), .ZN(n10972) );
  ND4D1BWP30P140LVT U11549 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(n11002) );
  AOI22D1BWP30P140LVT U11550 ( .A1(i_data_bus[703]), .A2(n10977), .B1(
        i_data_bus[191]), .B2(n10976), .ZN(n10987) );
  AOI22D1BWP30P140LVT U11551 ( .A1(i_data_bus[63]), .A2(n10979), .B1(
        i_data_bus[383]), .B2(n10978), .ZN(n10986) );
  AOI22D1BWP30P140LVT U11552 ( .A1(i_data_bus[607]), .A2(n10981), .B1(
        i_data_bus[319]), .B2(n10980), .ZN(n10985) );
  AOI22D1BWP30P140LVT U11553 ( .A1(i_data_bus[223]), .A2(n10983), .B1(
        i_data_bus[895]), .B2(n10982), .ZN(n10984) );
  ND4D1BWP30P140LVT U11554 ( .A1(n10987), .A2(n10986), .A3(n10985), .A4(n10984), .ZN(n11001) );
  AOI22D1BWP30P140LVT U11555 ( .A1(i_data_bus[511]), .A2(n10989), .B1(
        i_data_bus[767]), .B2(n10988), .ZN(n10999) );
  AOI22D1BWP30P140LVT U11556 ( .A1(i_data_bus[127]), .A2(n10991), .B1(
        i_data_bus[255]), .B2(n10990), .ZN(n10998) );
  AOI22D1BWP30P140LVT U11557 ( .A1(i_data_bus[863]), .A2(n10993), .B1(
        i_data_bus[479]), .B2(n10992), .ZN(n10997) );
  AOI22D1BWP30P140LVT U11558 ( .A1(i_data_bus[735]), .A2(n10995), .B1(
        i_data_bus[415]), .B2(n10994), .ZN(n10996) );
  ND4D1BWP30P140LVT U11559 ( .A1(n10999), .A2(n10998), .A3(n10997), .A4(n10996), .ZN(n11000) );
  OR4D1BWP30P140LVT U11560 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .Z(o_data_bus[223]) );
  NR3D0P7BWP30P140LVT U11561 ( .A1(n11717), .A2(n11004), .A3(n11013), .ZN(
        n11646) );
  INR3D0BWP30P140LVT U11562 ( .A1(i_cmd[9]), .B1(n11737), .B2(n11011), .ZN(
        n11648) );
  AOI22D1BWP30P140LVT U11563 ( .A1(i_data_bus[992]), .A2(n11646), .B1(
        i_data_bus[32]), .B2(n11648), .ZN(n11010) );
  INR3D0BWP30P140LVT U11564 ( .A1(i_cmd[137]), .B1(n11701), .B2(n11015), .ZN(
        n11650) );
  INR3D0BWP30P140LVT U11565 ( .A1(i_cmd[25]), .B1(n11011), .B2(n11726), .ZN(
        n11660) );
  AOI22D1BWP30P140LVT U11566 ( .A1(i_data_bus[544]), .A2(n11650), .B1(
        i_data_bus[96]), .B2(n11660), .ZN(n11009) );
  NR3D0P7BWP30P140LVT U11567 ( .A1(n6721), .A2(n11015), .A3(n11713), .ZN(
        n11658) );
  NR3D0P7BWP30P140LVT U11568 ( .A1(n11005), .A2(n11013), .A3(n11740), .ZN(
        n11659) );
  AOI22D1BWP30P140LVT U11569 ( .A1(i_data_bus[512]), .A2(n11658), .B1(
        i_data_bus[928]), .B2(n11659), .ZN(n11008) );
  INVD1BWP30P140LVT U11570 ( .I(i_cmd[1]), .ZN(n11006) );
  NR3D0P7BWP30P140LVT U11571 ( .A1(n11006), .A2(n11011), .A3(n11703), .ZN(
        n11652) );
  INR3D0BWP30P140LVT U11572 ( .A1(i_cmd[145]), .B1(n11015), .B2(n11733), .ZN(
        n11651) );
  AOI22D1BWP30P140LVT U11573 ( .A1(i_data_bus[0]), .A2(n11652), .B1(
        i_data_bus[576]), .B2(n11651), .ZN(n11007) );
  ND4D1BWP30P140LVT U11574 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(n11044) );
  INR3D0BWP30P140LVT U11575 ( .A1(i_cmd[17]), .B1(n11011), .B2(n11699), .ZN(
        n11645) );
  NR3D0P7BWP30P140LVT U11576 ( .A1(n11012), .A2(n11013), .A3(n11715), .ZN(
        n11647) );
  AOI22D1BWP30P140LVT U11577 ( .A1(i_data_bus[64]), .A2(n11645), .B1(
        i_data_bus[960]), .B2(n11647), .ZN(n11020) );
  NR3D0P7BWP30P140LVT U11578 ( .A1(n11014), .A2(n11013), .A3(n11735), .ZN(
        n11649) );
  INR3D0BWP30P140LVT U11579 ( .A1(i_cmd[153]), .B1(n11015), .B2(n11697), .ZN(
        n11657) );
  AOI22D1BWP30P140LVT U11580 ( .A1(i_data_bus[896]), .A2(n11649), .B1(
        i_data_bus[608]), .B2(n11657), .ZN(n11019) );
  NR3D0P7BWP30P140LVT U11581 ( .A1(n11016), .A2(n11705), .A3(n11024), .ZN(
        n11674) );
  INR3D0BWP30P140LVT U11582 ( .A1(i_cmd[121]), .B1(n11024), .B2(n11719), .ZN(
        n11664) );
  AOI22D1BWP30P140LVT U11583 ( .A1(i_data_bus[384]), .A2(n11674), .B1(
        i_data_bus[480]), .B2(n11664), .ZN(n11018) );
  INR3D0BWP30P140LVT U11584 ( .A1(i_cmd[105]), .B1(n11024), .B2(n11698), .ZN(
        n11662) );
  INR3D0BWP30P140LVT U11585 ( .A1(i_cmd[209]), .B1(n11745), .B2(n11034), .ZN(
        n11676) );
  AOI22D1BWP30P140LVT U11586 ( .A1(i_data_bus[416]), .A2(n11662), .B1(
        i_data_bus[832]), .B2(n11676), .ZN(n11017) );
  ND4D1BWP30P140LVT U11587 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(n11043) );
  NR3D0P7BWP30P140LVT U11588 ( .A1(n11021), .A2(n11747), .A3(n11031), .ZN(
        n11672) );
  INR3D0BWP30P140LVT U11589 ( .A1(i_cmd[185]), .B1(n11031), .B2(n11750), .ZN(
        n11671) );
  AOI22D1BWP30P140LVT U11590 ( .A1(i_data_bus[640]), .A2(n11672), .B1(
        i_data_bus[736]), .B2(n11671), .ZN(n11029) );
  NR3D0P7BWP30P140LVT U11591 ( .A1(n11022), .A2(n11034), .A3(n11754), .ZN(
        n11670) );
  INR3D0BWP30P140LVT U11592 ( .A1(i_cmd[41]), .B1(n11023), .B2(n11033), .ZN(
        n11684) );
  AOI22D1BWP30P140LVT U11593 ( .A1(i_data_bus[768]), .A2(n11670), .B1(
        i_data_bus[160]), .B2(n11684), .ZN(n11028) );
  INR3D0BWP30P140LVT U11594 ( .A1(i_cmd[113]), .B1(n11024), .B2(n11706), .ZN(
        n11686) );
  INVD1BWP30P140LVT U11595 ( .I(i_cmd[33]), .ZN(n11025) );
  NR3D0P7BWP30P140LVT U11596 ( .A1(n11025), .A2(n11033), .A3(n11721), .ZN(
        n11682) );
  AOI22D1BWP30P140LVT U11597 ( .A1(i_data_bus[448]), .A2(n11686), .B1(
        i_data_bus[128]), .B2(n11682), .ZN(n11027) );
  INR3D0BWP30P140LVT U11598 ( .A1(i_cmd[89]), .B1(n11731), .B2(n11035), .ZN(
        n11685) );
  INR3D0BWP30P140LVT U11599 ( .A1(i_cmd[177]), .B1(n11031), .B2(n11748), .ZN(
        n11669) );
  AOI22D1BWP30P140LVT U11600 ( .A1(i_data_bus[352]), .A2(n11685), .B1(
        i_data_bus[704]), .B2(n11669), .ZN(n11026) );
  ND4D1BWP30P140LVT U11601 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(n11042) );
  INR3D0BWP30P140LVT U11602 ( .A1(i_cmd[49]), .B1(n11033), .B2(n11030), .ZN(
        n11675) );
  INR3D0BWP30P140LVT U11603 ( .A1(i_cmd[169]), .B1(n11031), .B2(n11756), .ZN(
        n11683) );
  AOI22D1BWP30P140LVT U11604 ( .A1(i_data_bus[192]), .A2(n11675), .B1(
        i_data_bus[672]), .B2(n11683), .ZN(n11040) );
  INR3D0BWP30P140LVT U11605 ( .A1(i_cmd[57]), .B1(n11033), .B2(n11032), .ZN(
        n11688) );
  INR3D0BWP30P140LVT U11606 ( .A1(i_cmd[217]), .B1(n11034), .B2(n11749), .ZN(
        n11681) );
  AOI22D1BWP30P140LVT U11607 ( .A1(i_data_bus[224]), .A2(n11688), .B1(
        i_data_bus[864]), .B2(n11681), .ZN(n11039) );
  INR3D0BWP30P140LVT U11608 ( .A1(i_cmd[73]), .B1(n11035), .B2(n11711), .ZN(
        n11661) );
  INR3D0BWP30P140LVT U11609 ( .A1(i_cmd[201]), .B1(n11034), .B2(n11751), .ZN(
        n11673) );
  AOI22D1BWP30P140LVT U11610 ( .A1(i_data_bus[288]), .A2(n11661), .B1(
        i_data_bus[800]), .B2(n11673), .ZN(n11038) );
  INR3D0BWP30P140LVT U11611 ( .A1(i_cmd[81]), .B1(n11035), .B2(n11700), .ZN(
        n11687) );
  INVD1BWP30P140LVT U11612 ( .I(i_cmd[65]), .ZN(n11036) );
  NR3D0P7BWP30P140LVT U11613 ( .A1(n11036), .A2(n11035), .A3(n11728), .ZN(
        n11663) );
  AOI22D1BWP30P140LVT U11614 ( .A1(i_data_bus[320]), .A2(n11687), .B1(
        i_data_bus[256]), .B2(n11663), .ZN(n11037) );
  ND4D1BWP30P140LVT U11615 ( .A1(n11040), .A2(n11039), .A3(n11038), .A4(n11037), .ZN(n11041) );
  OR4D1BWP30P140LVT U11616 ( .A1(n11044), .A2(n11043), .A3(n11042), .A4(n11041), .Z(o_data_bus[32]) );
  AOI22D1BWP30P140LVT U11617 ( .A1(n11660), .A2(i_data_bus[97]), .B1(n11651), 
        .B2(i_data_bus[577]), .ZN(n11048) );
  AOI22D1BWP30P140LVT U11618 ( .A1(n11650), .A2(i_data_bus[545]), .B1(n11649), 
        .B2(i_data_bus[897]), .ZN(n11047) );
  AOI22D1BWP30P140LVT U11619 ( .A1(n11646), .A2(i_data_bus[993]), .B1(n11647), 
        .B2(i_data_bus[961]), .ZN(n11046) );
  AOI22D1BWP30P140LVT U11620 ( .A1(n11648), .A2(i_data_bus[33]), .B1(n11659), 
        .B2(i_data_bus[929]), .ZN(n11045) );
  ND4D1BWP30P140LVT U11621 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(n11064) );
  AOI22D1BWP30P140LVT U11622 ( .A1(n11645), .A2(i_data_bus[65]), .B1(n11657), 
        .B2(i_data_bus[609]), .ZN(n11052) );
  AOI22D1BWP30P140LVT U11623 ( .A1(n11658), .A2(i_data_bus[513]), .B1(n11652), 
        .B2(i_data_bus[1]), .ZN(n11051) );
  AOI22D1BWP30P140LVT U11624 ( .A1(n11670), .A2(i_data_bus[769]), .B1(n11669), 
        .B2(i_data_bus[705]), .ZN(n11050) );
  AOI22D1BWP30P140LVT U11625 ( .A1(n11674), .A2(i_data_bus[385]), .B1(n11683), 
        .B2(i_data_bus[673]), .ZN(n11049) );
  ND4D1BWP30P140LVT U11626 ( .A1(n11052), .A2(n11051), .A3(n11050), .A4(n11049), .ZN(n11063) );
  AOI22D1BWP30P140LVT U11627 ( .A1(n11672), .A2(i_data_bus[641]), .B1(n11681), 
        .B2(i_data_bus[865]), .ZN(n11056) );
  AOI22D1BWP30P140LVT U11628 ( .A1(n11664), .A2(i_data_bus[481]), .B1(n11673), 
        .B2(i_data_bus[801]), .ZN(n11055) );
  AOI22D1BWP30P140LVT U11629 ( .A1(n11684), .A2(i_data_bus[161]), .B1(n11685), 
        .B2(i_data_bus[353]), .ZN(n11054) );
  AOI22D1BWP30P140LVT U11630 ( .A1(n11688), .A2(i_data_bus[225]), .B1(n11663), 
        .B2(i_data_bus[257]), .ZN(n11053) );
  ND4D1BWP30P140LVT U11631 ( .A1(n11056), .A2(n11055), .A3(n11054), .A4(n11053), .ZN(n11062) );
  AOI22D1BWP30P140LVT U11632 ( .A1(n11686), .A2(i_data_bus[449]), .B1(n11661), 
        .B2(i_data_bus[289]), .ZN(n11060) );
  AOI22D1BWP30P140LVT U11633 ( .A1(n11671), .A2(i_data_bus[737]), .B1(n11675), 
        .B2(i_data_bus[193]), .ZN(n11059) );
  AOI22D1BWP30P140LVT U11634 ( .A1(n11662), .A2(i_data_bus[417]), .B1(n11682), 
        .B2(i_data_bus[129]), .ZN(n11058) );
  AOI22D1BWP30P140LVT U11635 ( .A1(n11676), .A2(i_data_bus[833]), .B1(n11687), 
        .B2(i_data_bus[321]), .ZN(n11057) );
  ND4D1BWP30P140LVT U11636 ( .A1(n11060), .A2(n11059), .A3(n11058), .A4(n11057), .ZN(n11061) );
  OR4D1BWP30P140LVT U11637 ( .A1(n11064), .A2(n11063), .A3(n11062), .A4(n11061), .Z(o_data_bus[33]) );
  AOI22D1BWP30P140LVT U11638 ( .A1(n11650), .A2(i_data_bus[546]), .B1(n11651), 
        .B2(i_data_bus[578]), .ZN(n11068) );
  AOI22D1BWP30P140LVT U11639 ( .A1(n11645), .A2(i_data_bus[66]), .B1(n11647), 
        .B2(i_data_bus[962]), .ZN(n11067) );
  AOI22D1BWP30P140LVT U11640 ( .A1(n11648), .A2(i_data_bus[34]), .B1(n11649), 
        .B2(i_data_bus[898]), .ZN(n11066) );
  AOI22D1BWP30P140LVT U11641 ( .A1(n11658), .A2(i_data_bus[514]), .B1(n11652), 
        .B2(i_data_bus[2]), .ZN(n11065) );
  ND4D1BWP30P140LVT U11642 ( .A1(n11068), .A2(n11067), .A3(n11066), .A4(n11065), .ZN(n11084) );
  AOI22D1BWP30P140LVT U11643 ( .A1(n11646), .A2(i_data_bus[994]), .B1(n11660), 
        .B2(i_data_bus[98]), .ZN(n11072) );
  AOI22D1BWP30P140LVT U11644 ( .A1(n11659), .A2(i_data_bus[930]), .B1(n11657), 
        .B2(i_data_bus[610]), .ZN(n11071) );
  AOI22D1BWP30P140LVT U11645 ( .A1(n11684), .A2(i_data_bus[162]), .B1(n11681), 
        .B2(i_data_bus[866]), .ZN(n11070) );
  AOI22D1BWP30P140LVT U11646 ( .A1(n11675), .A2(i_data_bus[194]), .B1(n11683), 
        .B2(i_data_bus[674]), .ZN(n11069) );
  ND4D1BWP30P140LVT U11647 ( .A1(n11072), .A2(n11071), .A3(n11070), .A4(n11069), .ZN(n11083) );
  AOI22D1BWP30P140LVT U11648 ( .A1(n11664), .A2(i_data_bus[482]), .B1(n11661), 
        .B2(i_data_bus[290]), .ZN(n11076) );
  AOI22D1BWP30P140LVT U11649 ( .A1(n11674), .A2(i_data_bus[386]), .B1(n11662), 
        .B2(i_data_bus[418]), .ZN(n11075) );
  AOI22D1BWP30P140LVT U11650 ( .A1(n11686), .A2(i_data_bus[450]), .B1(n11673), 
        .B2(i_data_bus[802]), .ZN(n11074) );
  AOI22D1BWP30P140LVT U11651 ( .A1(n11670), .A2(i_data_bus[770]), .B1(n11688), 
        .B2(i_data_bus[226]), .ZN(n11073) );
  ND4D1BWP30P140LVT U11652 ( .A1(n11076), .A2(n11075), .A3(n11074), .A4(n11073), .ZN(n11082) );
  AOI22D1BWP30P140LVT U11653 ( .A1(n11676), .A2(i_data_bus[834]), .B1(n11671), 
        .B2(i_data_bus[738]), .ZN(n11080) );
  AOI22D1BWP30P140LVT U11654 ( .A1(n11685), .A2(i_data_bus[354]), .B1(n11669), 
        .B2(i_data_bus[706]), .ZN(n11079) );
  AOI22D1BWP30P140LVT U11655 ( .A1(n11672), .A2(i_data_bus[642]), .B1(n11682), 
        .B2(i_data_bus[130]), .ZN(n11078) );
  AOI22D1BWP30P140LVT U11656 ( .A1(n11687), .A2(i_data_bus[322]), .B1(n11663), 
        .B2(i_data_bus[258]), .ZN(n11077) );
  ND4D1BWP30P140LVT U11657 ( .A1(n11080), .A2(n11079), .A3(n11078), .A4(n11077), .ZN(n11081) );
  OR4D1BWP30P140LVT U11658 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .Z(o_data_bus[34]) );
  AOI22D1BWP30P140LVT U11659 ( .A1(n11658), .A2(i_data_bus[515]), .B1(n11645), 
        .B2(i_data_bus[67]), .ZN(n11088) );
  AOI22D1BWP30P140LVT U11660 ( .A1(n11651), .A2(i_data_bus[579]), .B1(n11649), 
        .B2(i_data_bus[899]), .ZN(n11087) );
  AOI22D1BWP30P140LVT U11661 ( .A1(n11648), .A2(i_data_bus[35]), .B1(n11652), 
        .B2(i_data_bus[3]), .ZN(n11086) );
  AOI22D1BWP30P140LVT U11662 ( .A1(n11660), .A2(i_data_bus[99]), .B1(n11647), 
        .B2(i_data_bus[963]), .ZN(n11085) );
  ND4D1BWP30P140LVT U11663 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(n11104) );
  AOI22D1BWP30P140LVT U11664 ( .A1(n11650), .A2(i_data_bus[547]), .B1(n11657), 
        .B2(i_data_bus[611]), .ZN(n11092) );
  AOI22D1BWP30P140LVT U11665 ( .A1(n11646), .A2(i_data_bus[995]), .B1(n11659), 
        .B2(i_data_bus[931]), .ZN(n11091) );
  AOI22D1BWP30P140LVT U11666 ( .A1(n11685), .A2(i_data_bus[355]), .B1(n11663), 
        .B2(i_data_bus[259]), .ZN(n11090) );
  AOI22D1BWP30P140LVT U11667 ( .A1(n11674), .A2(i_data_bus[387]), .B1(n11676), 
        .B2(i_data_bus[835]), .ZN(n11089) );
  ND4D1BWP30P140LVT U11668 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(n11103) );
  AOI22D1BWP30P140LVT U11669 ( .A1(n11664), .A2(i_data_bus[483]), .B1(n11662), 
        .B2(i_data_bus[419]), .ZN(n11096) );
  AOI22D1BWP30P140LVT U11670 ( .A1(n11682), .A2(i_data_bus[131]), .B1(n11687), 
        .B2(i_data_bus[323]), .ZN(n11095) );
  AOI22D1BWP30P140LVT U11671 ( .A1(n11671), .A2(i_data_bus[739]), .B1(n11670), 
        .B2(i_data_bus[771]), .ZN(n11094) );
  AOI22D1BWP30P140LVT U11672 ( .A1(n11684), .A2(i_data_bus[163]), .B1(n11683), 
        .B2(i_data_bus[675]), .ZN(n11093) );
  ND4D1BWP30P140LVT U11673 ( .A1(n11096), .A2(n11095), .A3(n11094), .A4(n11093), .ZN(n11102) );
  AOI22D1BWP30P140LVT U11674 ( .A1(n11672), .A2(i_data_bus[643]), .B1(n11688), 
        .B2(i_data_bus[227]), .ZN(n11100) );
  AOI22D1BWP30P140LVT U11675 ( .A1(n11681), .A2(i_data_bus[867]), .B1(n11661), 
        .B2(i_data_bus[291]), .ZN(n11099) );
  AOI22D1BWP30P140LVT U11676 ( .A1(n11669), .A2(i_data_bus[707]), .B1(n11673), 
        .B2(i_data_bus[803]), .ZN(n11098) );
  AOI22D1BWP30P140LVT U11677 ( .A1(n11686), .A2(i_data_bus[451]), .B1(n11675), 
        .B2(i_data_bus[195]), .ZN(n11097) );
  ND4D1BWP30P140LVT U11678 ( .A1(n11100), .A2(n11099), .A3(n11098), .A4(n11097), .ZN(n11101) );
  OR4D1BWP30P140LVT U11679 ( .A1(n11104), .A2(n11103), .A3(n11102), .A4(n11101), .Z(o_data_bus[35]) );
  AOI22D1BWP30P140LVT U11680 ( .A1(n11650), .A2(i_data_bus[548]), .B1(n11660), 
        .B2(i_data_bus[100]), .ZN(n11108) );
  AOI22D1BWP30P140LVT U11681 ( .A1(n11647), .A2(i_data_bus[964]), .B1(n11657), 
        .B2(i_data_bus[612]), .ZN(n11107) );
  AOI22D1BWP30P140LVT U11682 ( .A1(n11659), .A2(i_data_bus[932]), .B1(n11649), 
        .B2(i_data_bus[900]), .ZN(n11106) );
  AOI22D1BWP30P140LVT U11683 ( .A1(n11658), .A2(i_data_bus[516]), .B1(n11645), 
        .B2(i_data_bus[68]), .ZN(n11105) );
  ND4D1BWP30P140LVT U11684 ( .A1(n11108), .A2(n11107), .A3(n11106), .A4(n11105), .ZN(n11124) );
  AOI22D1BWP30P140LVT U11685 ( .A1(n11646), .A2(i_data_bus[996]), .B1(n11648), 
        .B2(i_data_bus[36]), .ZN(n11112) );
  AOI22D1BWP30P140LVT U11686 ( .A1(n11652), .A2(i_data_bus[4]), .B1(n11651), 
        .B2(i_data_bus[580]), .ZN(n11111) );
  AOI22D1BWP30P140LVT U11687 ( .A1(n11671), .A2(i_data_bus[740]), .B1(n11675), 
        .B2(i_data_bus[196]), .ZN(n11110) );
  AOI22D1BWP30P140LVT U11688 ( .A1(n11670), .A2(i_data_bus[772]), .B1(n11669), 
        .B2(i_data_bus[708]), .ZN(n11109) );
  ND4D1BWP30P140LVT U11689 ( .A1(n11112), .A2(n11111), .A3(n11110), .A4(n11109), .ZN(n11123) );
  AOI22D1BWP30P140LVT U11690 ( .A1(n11682), .A2(i_data_bus[132]), .B1(n11688), 
        .B2(i_data_bus[228]), .ZN(n11116) );
  AOI22D1BWP30P140LVT U11691 ( .A1(n11662), .A2(i_data_bus[420]), .B1(n11686), 
        .B2(i_data_bus[452]), .ZN(n11115) );
  AOI22D1BWP30P140LVT U11692 ( .A1(n11664), .A2(i_data_bus[484]), .B1(n11681), 
        .B2(i_data_bus[868]), .ZN(n11114) );
  AOI22D1BWP30P140LVT U11693 ( .A1(n11684), .A2(i_data_bus[164]), .B1(n11683), 
        .B2(i_data_bus[676]), .ZN(n11113) );
  ND4D1BWP30P140LVT U11694 ( .A1(n11116), .A2(n11115), .A3(n11114), .A4(n11113), .ZN(n11122) );
  AOI22D1BWP30P140LVT U11695 ( .A1(n11661), .A2(i_data_bus[292]), .B1(n11687), 
        .B2(i_data_bus[324]), .ZN(n11120) );
  AOI22D1BWP30P140LVT U11696 ( .A1(n11672), .A2(i_data_bus[644]), .B1(n11685), 
        .B2(i_data_bus[356]), .ZN(n11119) );
  AOI22D1BWP30P140LVT U11697 ( .A1(n11676), .A2(i_data_bus[836]), .B1(n11663), 
        .B2(i_data_bus[260]), .ZN(n11118) );
  AOI22D1BWP30P140LVT U11698 ( .A1(n11674), .A2(i_data_bus[388]), .B1(n11673), 
        .B2(i_data_bus[804]), .ZN(n11117) );
  ND4D1BWP30P140LVT U11699 ( .A1(n11120), .A2(n11119), .A3(n11118), .A4(n11117), .ZN(n11121) );
  OR4D1BWP30P140LVT U11700 ( .A1(n11124), .A2(n11123), .A3(n11122), .A4(n11121), .Z(o_data_bus[36]) );
  AOI22D1BWP30P140LVT U11701 ( .A1(n11658), .A2(i_data_bus[517]), .B1(n11649), 
        .B2(i_data_bus[901]), .ZN(n11128) );
  AOI22D1BWP30P140LVT U11702 ( .A1(n11648), .A2(i_data_bus[37]), .B1(n11650), 
        .B2(i_data_bus[549]), .ZN(n11127) );
  AOI22D1BWP30P140LVT U11703 ( .A1(n11652), .A2(i_data_bus[5]), .B1(n11651), 
        .B2(i_data_bus[581]), .ZN(n11126) );
  AOI22D1BWP30P140LVT U11704 ( .A1(n11660), .A2(i_data_bus[101]), .B1(n11659), 
        .B2(i_data_bus[933]), .ZN(n11125) );
  ND4D1BWP30P140LVT U11705 ( .A1(n11128), .A2(n11127), .A3(n11126), .A4(n11125), .ZN(n11144) );
  AOI22D1BWP30P140LVT U11706 ( .A1(n11647), .A2(i_data_bus[965]), .B1(n11657), 
        .B2(i_data_bus[613]), .ZN(n11132) );
  AOI22D1BWP30P140LVT U11707 ( .A1(n11646), .A2(i_data_bus[997]), .B1(n11645), 
        .B2(i_data_bus[69]), .ZN(n11131) );
  AOI22D1BWP30P140LVT U11708 ( .A1(n11670), .A2(i_data_bus[773]), .B1(n11675), 
        .B2(i_data_bus[197]), .ZN(n11130) );
  AOI22D1BWP30P140LVT U11709 ( .A1(n11672), .A2(i_data_bus[645]), .B1(n11683), 
        .B2(i_data_bus[677]), .ZN(n11129) );
  ND4D1BWP30P140LVT U11710 ( .A1(n11132), .A2(n11131), .A3(n11130), .A4(n11129), .ZN(n11143) );
  AOI22D1BWP30P140LVT U11711 ( .A1(n11676), .A2(i_data_bus[837]), .B1(n11673), 
        .B2(i_data_bus[805]), .ZN(n11136) );
  AOI22D1BWP30P140LVT U11712 ( .A1(n11684), .A2(i_data_bus[165]), .B1(n11681), 
        .B2(i_data_bus[869]), .ZN(n11135) );
  AOI22D1BWP30P140LVT U11713 ( .A1(n11686), .A2(i_data_bus[453]), .B1(n11669), 
        .B2(i_data_bus[709]), .ZN(n11134) );
  AOI22D1BWP30P140LVT U11714 ( .A1(n11664), .A2(i_data_bus[485]), .B1(n11685), 
        .B2(i_data_bus[357]), .ZN(n11133) );
  ND4D1BWP30P140LVT U11715 ( .A1(n11136), .A2(n11135), .A3(n11134), .A4(n11133), .ZN(n11142) );
  AOI22D1BWP30P140LVT U11716 ( .A1(n11662), .A2(i_data_bus[421]), .B1(n11661), 
        .B2(i_data_bus[293]), .ZN(n11140) );
  AOI22D1BWP30P140LVT U11717 ( .A1(n11671), .A2(i_data_bus[741]), .B1(n11682), 
        .B2(i_data_bus[133]), .ZN(n11139) );
  AOI22D1BWP30P140LVT U11718 ( .A1(n11687), .A2(i_data_bus[325]), .B1(n11663), 
        .B2(i_data_bus[261]), .ZN(n11138) );
  AOI22D1BWP30P140LVT U11719 ( .A1(n11674), .A2(i_data_bus[389]), .B1(n11688), 
        .B2(i_data_bus[229]), .ZN(n11137) );
  ND4D1BWP30P140LVT U11720 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(n11141) );
  OR4D1BWP30P140LVT U11721 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .Z(o_data_bus[37]) );
  AOI22D1BWP30P140LVT U11722 ( .A1(n11651), .A2(i_data_bus[582]), .B1(n11647), 
        .B2(i_data_bus[966]), .ZN(n11148) );
  AOI22D1BWP30P140LVT U11723 ( .A1(n11650), .A2(i_data_bus[550]), .B1(n11657), 
        .B2(i_data_bus[614]), .ZN(n11147) );
  AOI22D1BWP30P140LVT U11724 ( .A1(n11648), .A2(i_data_bus[38]), .B1(n11659), 
        .B2(i_data_bus[934]), .ZN(n11146) );
  AOI22D1BWP30P140LVT U11725 ( .A1(n11652), .A2(i_data_bus[6]), .B1(n11645), 
        .B2(i_data_bus[70]), .ZN(n11145) );
  ND4D1BWP30P140LVT U11726 ( .A1(n11148), .A2(n11147), .A3(n11146), .A4(n11145), .ZN(n11164) );
  AOI22D1BWP30P140LVT U11727 ( .A1(n11660), .A2(i_data_bus[102]), .B1(n11658), 
        .B2(i_data_bus[518]), .ZN(n11152) );
  AOI22D1BWP30P140LVT U11728 ( .A1(n11646), .A2(i_data_bus[998]), .B1(n11649), 
        .B2(i_data_bus[902]), .ZN(n11151) );
  AOI22D1BWP30P140LVT U11729 ( .A1(n11681), .A2(i_data_bus[870]), .B1(n11673), 
        .B2(i_data_bus[806]), .ZN(n11150) );
  AOI22D1BWP30P140LVT U11730 ( .A1(n11664), .A2(i_data_bus[486]), .B1(n11676), 
        .B2(i_data_bus[838]), .ZN(n11149) );
  ND4D1BWP30P140LVT U11731 ( .A1(n11152), .A2(n11151), .A3(n11150), .A4(n11149), .ZN(n11163) );
  AOI22D1BWP30P140LVT U11732 ( .A1(n11671), .A2(i_data_bus[742]), .B1(n11688), 
        .B2(i_data_bus[230]), .ZN(n11156) );
  AOI22D1BWP30P140LVT U11733 ( .A1(n11672), .A2(i_data_bus[646]), .B1(n11684), 
        .B2(i_data_bus[166]), .ZN(n11155) );
  AOI22D1BWP30P140LVT U11734 ( .A1(n11674), .A2(i_data_bus[390]), .B1(n11686), 
        .B2(i_data_bus[454]), .ZN(n11154) );
  AOI22D1BWP30P140LVT U11735 ( .A1(n11685), .A2(i_data_bus[358]), .B1(n11669), 
        .B2(i_data_bus[710]), .ZN(n11153) );
  ND4D1BWP30P140LVT U11736 ( .A1(n11156), .A2(n11155), .A3(n11154), .A4(n11153), .ZN(n11162) );
  AOI22D1BWP30P140LVT U11737 ( .A1(n11670), .A2(i_data_bus[774]), .B1(n11675), 
        .B2(i_data_bus[198]), .ZN(n11160) );
  AOI22D1BWP30P140LVT U11738 ( .A1(n11662), .A2(i_data_bus[422]), .B1(n11661), 
        .B2(i_data_bus[294]), .ZN(n11159) );
  AOI22D1BWP30P140LVT U11739 ( .A1(n11682), .A2(i_data_bus[134]), .B1(n11683), 
        .B2(i_data_bus[678]), .ZN(n11158) );
  AOI22D1BWP30P140LVT U11740 ( .A1(n11687), .A2(i_data_bus[326]), .B1(n11663), 
        .B2(i_data_bus[262]), .ZN(n11157) );
  ND4D1BWP30P140LVT U11741 ( .A1(n11160), .A2(n11159), .A3(n11158), .A4(n11157), .ZN(n11161) );
  OR4D1BWP30P140LVT U11742 ( .A1(n11164), .A2(n11163), .A3(n11162), .A4(n11161), .Z(o_data_bus[38]) );
  AOI22D1BWP30P140LVT U11743 ( .A1(n11648), .A2(i_data_bus[39]), .B1(n11657), 
        .B2(i_data_bus[615]), .ZN(n11168) );
  AOI22D1BWP30P140LVT U11744 ( .A1(n11658), .A2(i_data_bus[519]), .B1(n11649), 
        .B2(i_data_bus[903]), .ZN(n11167) );
  AOI22D1BWP30P140LVT U11745 ( .A1(n11650), .A2(i_data_bus[551]), .B1(n11651), 
        .B2(i_data_bus[583]), .ZN(n11166) );
  AOI22D1BWP30P140LVT U11746 ( .A1(n11660), .A2(i_data_bus[103]), .B1(n11647), 
        .B2(i_data_bus[967]), .ZN(n11165) );
  ND4D1BWP30P140LVT U11747 ( .A1(n11168), .A2(n11167), .A3(n11166), .A4(n11165), .ZN(n11184) );
  AOI22D1BWP30P140LVT U11748 ( .A1(n11646), .A2(i_data_bus[999]), .B1(n11659), 
        .B2(i_data_bus[935]), .ZN(n11172) );
  AOI22D1BWP30P140LVT U11749 ( .A1(n11652), .A2(i_data_bus[7]), .B1(n11645), 
        .B2(i_data_bus[71]), .ZN(n11171) );
  AOI22D1BWP30P140LVT U11750 ( .A1(n11686), .A2(i_data_bus[455]), .B1(n11685), 
        .B2(i_data_bus[359]), .ZN(n11170) );
  AOI22D1BWP30P140LVT U11751 ( .A1(n11681), .A2(i_data_bus[871]), .B1(n11663), 
        .B2(i_data_bus[263]), .ZN(n11169) );
  ND4D1BWP30P140LVT U11752 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(n11183) );
  AOI22D1BWP30P140LVT U11753 ( .A1(n11674), .A2(i_data_bus[391]), .B1(n11683), 
        .B2(i_data_bus[679]), .ZN(n11176) );
  AOI22D1BWP30P140LVT U11754 ( .A1(n11664), .A2(i_data_bus[487]), .B1(n11673), 
        .B2(i_data_bus[807]), .ZN(n11175) );
  AOI22D1BWP30P140LVT U11755 ( .A1(n11676), .A2(i_data_bus[839]), .B1(n11671), 
        .B2(i_data_bus[743]), .ZN(n11174) );
  AOI22D1BWP30P140LVT U11756 ( .A1(n11670), .A2(i_data_bus[775]), .B1(n11669), 
        .B2(i_data_bus[711]), .ZN(n11173) );
  ND4D1BWP30P140LVT U11757 ( .A1(n11176), .A2(n11175), .A3(n11174), .A4(n11173), .ZN(n11182) );
  AOI22D1BWP30P140LVT U11758 ( .A1(n11684), .A2(i_data_bus[167]), .B1(n11682), 
        .B2(i_data_bus[135]), .ZN(n11180) );
  AOI22D1BWP30P140LVT U11759 ( .A1(n11672), .A2(i_data_bus[647]), .B1(n11661), 
        .B2(i_data_bus[295]), .ZN(n11179) );
  AOI22D1BWP30P140LVT U11760 ( .A1(n11662), .A2(i_data_bus[423]), .B1(n11687), 
        .B2(i_data_bus[327]), .ZN(n11178) );
  AOI22D1BWP30P140LVT U11761 ( .A1(n11675), .A2(i_data_bus[199]), .B1(n11688), 
        .B2(i_data_bus[231]), .ZN(n11177) );
  ND4D1BWP30P140LVT U11762 ( .A1(n11180), .A2(n11179), .A3(n11178), .A4(n11177), .ZN(n11181) );
  OR4D1BWP30P140LVT U11763 ( .A1(n11184), .A2(n11183), .A3(n11182), .A4(n11181), .Z(o_data_bus[39]) );
  AOI22D1BWP30P140LVT U11764 ( .A1(n11652), .A2(i_data_bus[8]), .B1(n11647), 
        .B2(i_data_bus[968]), .ZN(n11188) );
  AOI22D1BWP30P140LVT U11765 ( .A1(n11659), .A2(i_data_bus[936]), .B1(n11657), 
        .B2(i_data_bus[616]), .ZN(n11187) );
  AOI22D1BWP30P140LVT U11766 ( .A1(n11650), .A2(i_data_bus[552]), .B1(n11660), 
        .B2(i_data_bus[104]), .ZN(n11186) );
  AOI22D1BWP30P140LVT U11767 ( .A1(n11646), .A2(i_data_bus[1000]), .B1(n11649), 
        .B2(i_data_bus[904]), .ZN(n11185) );
  ND4D1BWP30P140LVT U11768 ( .A1(n11188), .A2(n11187), .A3(n11186), .A4(n11185), .ZN(n11204) );
  AOI22D1BWP30P140LVT U11769 ( .A1(n11658), .A2(i_data_bus[520]), .B1(n11651), 
        .B2(i_data_bus[584]), .ZN(n11192) );
  AOI22D1BWP30P140LVT U11770 ( .A1(n11648), .A2(i_data_bus[40]), .B1(n11645), 
        .B2(i_data_bus[72]), .ZN(n11191) );
  AOI22D1BWP30P140LVT U11771 ( .A1(n11686), .A2(i_data_bus[456]), .B1(n11663), 
        .B2(i_data_bus[264]), .ZN(n11190) );
  AOI22D1BWP30P140LVT U11772 ( .A1(n11662), .A2(i_data_bus[424]), .B1(n11684), 
        .B2(i_data_bus[168]), .ZN(n11189) );
  ND4D1BWP30P140LVT U11773 ( .A1(n11192), .A2(n11191), .A3(n11190), .A4(n11189), .ZN(n11203) );
  AOI22D1BWP30P140LVT U11774 ( .A1(n11676), .A2(i_data_bus[840]), .B1(n11671), 
        .B2(i_data_bus[744]), .ZN(n11196) );
  AOI22D1BWP30P140LVT U11775 ( .A1(n11683), .A2(i_data_bus[680]), .B1(n11687), 
        .B2(i_data_bus[328]), .ZN(n11195) );
  AOI22D1BWP30P140LVT U11776 ( .A1(n11675), .A2(i_data_bus[200]), .B1(n11673), 
        .B2(i_data_bus[808]), .ZN(n11194) );
  AOI22D1BWP30P140LVT U11777 ( .A1(n11664), .A2(i_data_bus[488]), .B1(n11661), 
        .B2(i_data_bus[296]), .ZN(n11193) );
  ND4D1BWP30P140LVT U11778 ( .A1(n11196), .A2(n11195), .A3(n11194), .A4(n11193), .ZN(n11202) );
  AOI22D1BWP30P140LVT U11779 ( .A1(n11669), .A2(i_data_bus[712]), .B1(n11681), 
        .B2(i_data_bus[872]), .ZN(n11200) );
  AOI22D1BWP30P140LVT U11780 ( .A1(n11674), .A2(i_data_bus[392]), .B1(n11685), 
        .B2(i_data_bus[360]), .ZN(n11199) );
  AOI22D1BWP30P140LVT U11781 ( .A1(n11682), .A2(i_data_bus[136]), .B1(n11688), 
        .B2(i_data_bus[232]), .ZN(n11198) );
  AOI22D1BWP30P140LVT U11782 ( .A1(n11672), .A2(i_data_bus[648]), .B1(n11670), 
        .B2(i_data_bus[776]), .ZN(n11197) );
  ND4D1BWP30P140LVT U11783 ( .A1(n11200), .A2(n11199), .A3(n11198), .A4(n11197), .ZN(n11201) );
  OR4D1BWP30P140LVT U11784 ( .A1(n11204), .A2(n11203), .A3(n11202), .A4(n11201), .Z(o_data_bus[40]) );
  AOI22D1BWP30P140LVT U11785 ( .A1(n11658), .A2(i_data_bus[521]), .B1(n11652), 
        .B2(i_data_bus[9]), .ZN(n11208) );
  AOI22D1BWP30P140LVT U11786 ( .A1(n11645), .A2(i_data_bus[73]), .B1(n11649), 
        .B2(i_data_bus[905]), .ZN(n11207) );
  AOI22D1BWP30P140LVT U11787 ( .A1(n11651), .A2(i_data_bus[585]), .B1(n11657), 
        .B2(i_data_bus[617]), .ZN(n11206) );
  AOI22D1BWP30P140LVT U11788 ( .A1(n11650), .A2(i_data_bus[553]), .B1(n11660), 
        .B2(i_data_bus[105]), .ZN(n11205) );
  ND4D1BWP30P140LVT U11789 ( .A1(n11208), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(n11224) );
  AOI22D1BWP30P140LVT U11790 ( .A1(n11646), .A2(i_data_bus[1001]), .B1(n11647), 
        .B2(i_data_bus[969]), .ZN(n11212) );
  AOI22D1BWP30P140LVT U11791 ( .A1(n11648), .A2(i_data_bus[41]), .B1(n11659), 
        .B2(i_data_bus[937]), .ZN(n11211) );
  AOI22D1BWP30P140LVT U11792 ( .A1(n11664), .A2(i_data_bus[489]), .B1(n11675), 
        .B2(i_data_bus[201]), .ZN(n11210) );
  AOI22D1BWP30P140LVT U11793 ( .A1(n11671), .A2(i_data_bus[745]), .B1(n11688), 
        .B2(i_data_bus[233]), .ZN(n11209) );
  ND4D1BWP30P140LVT U11794 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(n11223) );
  AOI22D1BWP30P140LVT U11795 ( .A1(n11683), .A2(i_data_bus[681]), .B1(n11661), 
        .B2(i_data_bus[297]), .ZN(n11216) );
  AOI22D1BWP30P140LVT U11796 ( .A1(n11684), .A2(i_data_bus[169]), .B1(n11681), 
        .B2(i_data_bus[873]), .ZN(n11215) );
  AOI22D1BWP30P140LVT U11797 ( .A1(n11682), .A2(i_data_bus[137]), .B1(n11687), 
        .B2(i_data_bus[329]), .ZN(n11214) );
  AOI22D1BWP30P140LVT U11798 ( .A1(n11662), .A2(i_data_bus[425]), .B1(n11669), 
        .B2(i_data_bus[713]), .ZN(n11213) );
  ND4D1BWP30P140LVT U11799 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(n11222) );
  AOI22D1BWP30P140LVT U11800 ( .A1(n11673), .A2(i_data_bus[809]), .B1(n11663), 
        .B2(i_data_bus[265]), .ZN(n11220) );
  AOI22D1BWP30P140LVT U11801 ( .A1(n11670), .A2(i_data_bus[777]), .B1(n11685), 
        .B2(i_data_bus[361]), .ZN(n11219) );
  AOI22D1BWP30P140LVT U11802 ( .A1(n11674), .A2(i_data_bus[393]), .B1(n11686), 
        .B2(i_data_bus[457]), .ZN(n11218) );
  AOI22D1BWP30P140LVT U11803 ( .A1(n11676), .A2(i_data_bus[841]), .B1(n11672), 
        .B2(i_data_bus[649]), .ZN(n11217) );
  ND4D1BWP30P140LVT U11804 ( .A1(n11220), .A2(n11219), .A3(n11218), .A4(n11217), .ZN(n11221) );
  OR4D1BWP30P140LVT U11805 ( .A1(n11224), .A2(n11223), .A3(n11222), .A4(n11221), .Z(o_data_bus[41]) );
  AOI22D1BWP30P140LVT U11806 ( .A1(n11646), .A2(i_data_bus[1002]), .B1(n11650), 
        .B2(i_data_bus[554]), .ZN(n11228) );
  AOI22D1BWP30P140LVT U11807 ( .A1(n11648), .A2(i_data_bus[42]), .B1(n11652), 
        .B2(i_data_bus[10]), .ZN(n11227) );
  AOI22D1BWP30P140LVT U11808 ( .A1(n11647), .A2(i_data_bus[970]), .B1(n11657), 
        .B2(i_data_bus[618]), .ZN(n11226) );
  AOI22D1BWP30P140LVT U11809 ( .A1(n11660), .A2(i_data_bus[106]), .B1(n11645), 
        .B2(i_data_bus[74]), .ZN(n11225) );
  ND4D1BWP30P140LVT U11810 ( .A1(n11228), .A2(n11227), .A3(n11226), .A4(n11225), .ZN(n11244) );
  AOI22D1BWP30P140LVT U11811 ( .A1(n11651), .A2(i_data_bus[586]), .B1(n11649), 
        .B2(i_data_bus[906]), .ZN(n11232) );
  AOI22D1BWP30P140LVT U11812 ( .A1(n11658), .A2(i_data_bus[522]), .B1(n11659), 
        .B2(i_data_bus[938]), .ZN(n11231) );
  AOI22D1BWP30P140LVT U11813 ( .A1(n11675), .A2(i_data_bus[202]), .B1(n11687), 
        .B2(i_data_bus[330]), .ZN(n11230) );
  AOI22D1BWP30P140LVT U11814 ( .A1(n11664), .A2(i_data_bus[490]), .B1(n11688), 
        .B2(i_data_bus[234]), .ZN(n11229) );
  ND4D1BWP30P140LVT U11815 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(n11243) );
  AOI22D1BWP30P140LVT U11816 ( .A1(n11672), .A2(i_data_bus[650]), .B1(n11670), 
        .B2(i_data_bus[778]), .ZN(n11236) );
  AOI22D1BWP30P140LVT U11817 ( .A1(n11676), .A2(i_data_bus[842]), .B1(n11684), 
        .B2(i_data_bus[170]), .ZN(n11235) );
  AOI22D1BWP30P140LVT U11818 ( .A1(n11685), .A2(i_data_bus[362]), .B1(n11661), 
        .B2(i_data_bus[298]), .ZN(n11234) );
  AOI22D1BWP30P140LVT U11819 ( .A1(n11674), .A2(i_data_bus[394]), .B1(n11681), 
        .B2(i_data_bus[874]), .ZN(n11233) );
  ND4D1BWP30P140LVT U11820 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(n11242) );
  AOI22D1BWP30P140LVT U11821 ( .A1(n11662), .A2(i_data_bus[426]), .B1(n11686), 
        .B2(i_data_bus[458]), .ZN(n11240) );
  AOI22D1BWP30P140LVT U11822 ( .A1(n11669), .A2(i_data_bus[714]), .B1(n11673), 
        .B2(i_data_bus[810]), .ZN(n11239) );
  AOI22D1BWP30P140LVT U11823 ( .A1(n11671), .A2(i_data_bus[746]), .B1(n11683), 
        .B2(i_data_bus[682]), .ZN(n11238) );
  AOI22D1BWP30P140LVT U11824 ( .A1(n11682), .A2(i_data_bus[138]), .B1(n11663), 
        .B2(i_data_bus[266]), .ZN(n11237) );
  ND4D1BWP30P140LVT U11825 ( .A1(n11240), .A2(n11239), .A3(n11238), .A4(n11237), .ZN(n11241) );
  OR4D1BWP30P140LVT U11826 ( .A1(n11244), .A2(n11243), .A3(n11242), .A4(n11241), .Z(o_data_bus[42]) );
  AOI22D1BWP30P140LVT U11827 ( .A1(n11658), .A2(i_data_bus[523]), .B1(n11659), 
        .B2(i_data_bus[939]), .ZN(n11248) );
  AOI22D1BWP30P140LVT U11828 ( .A1(n11649), .A2(i_data_bus[907]), .B1(n11657), 
        .B2(i_data_bus[619]), .ZN(n11247) );
  AOI22D1BWP30P140LVT U11829 ( .A1(n11646), .A2(i_data_bus[1003]), .B1(n11652), 
        .B2(i_data_bus[11]), .ZN(n11246) );
  AOI22D1BWP30P140LVT U11830 ( .A1(n11660), .A2(i_data_bus[107]), .B1(n11647), 
        .B2(i_data_bus[971]), .ZN(n11245) );
  ND4D1BWP30P140LVT U11831 ( .A1(n11248), .A2(n11247), .A3(n11246), .A4(n11245), .ZN(n11264) );
  AOI22D1BWP30P140LVT U11832 ( .A1(n11648), .A2(i_data_bus[43]), .B1(n11645), 
        .B2(i_data_bus[75]), .ZN(n11252) );
  AOI22D1BWP30P140LVT U11833 ( .A1(n11650), .A2(i_data_bus[555]), .B1(n11651), 
        .B2(i_data_bus[587]), .ZN(n11251) );
  AOI22D1BWP30P140LVT U11834 ( .A1(n11685), .A2(i_data_bus[363]), .B1(n11675), 
        .B2(i_data_bus[203]), .ZN(n11250) );
  AOI22D1BWP30P140LVT U11835 ( .A1(n11664), .A2(i_data_bus[491]), .B1(n11662), 
        .B2(i_data_bus[427]), .ZN(n11249) );
  ND4D1BWP30P140LVT U11836 ( .A1(n11252), .A2(n11251), .A3(n11250), .A4(n11249), .ZN(n11263) );
  AOI22D1BWP30P140LVT U11837 ( .A1(n11674), .A2(i_data_bus[395]), .B1(n11684), 
        .B2(i_data_bus[171]), .ZN(n11256) );
  AOI22D1BWP30P140LVT U11838 ( .A1(n11686), .A2(i_data_bus[459]), .B1(n11681), 
        .B2(i_data_bus[875]), .ZN(n11255) );
  AOI22D1BWP30P140LVT U11839 ( .A1(n11671), .A2(i_data_bus[747]), .B1(n11682), 
        .B2(i_data_bus[139]), .ZN(n11254) );
  AOI22D1BWP30P140LVT U11840 ( .A1(n11676), .A2(i_data_bus[843]), .B1(n11673), 
        .B2(i_data_bus[811]), .ZN(n11253) );
  ND4D1BWP30P140LVT U11841 ( .A1(n11256), .A2(n11255), .A3(n11254), .A4(n11253), .ZN(n11262) );
  AOI22D1BWP30P140LVT U11842 ( .A1(n11670), .A2(i_data_bus[779]), .B1(n11688), 
        .B2(i_data_bus[235]), .ZN(n11260) );
  AOI22D1BWP30P140LVT U11843 ( .A1(n11661), .A2(i_data_bus[299]), .B1(n11687), 
        .B2(i_data_bus[331]), .ZN(n11259) );
  AOI22D1BWP30P140LVT U11844 ( .A1(n11672), .A2(i_data_bus[651]), .B1(n11683), 
        .B2(i_data_bus[683]), .ZN(n11258) );
  AOI22D1BWP30P140LVT U11845 ( .A1(n11669), .A2(i_data_bus[715]), .B1(n11663), 
        .B2(i_data_bus[267]), .ZN(n11257) );
  ND4D1BWP30P140LVT U11846 ( .A1(n11260), .A2(n11259), .A3(n11258), .A4(n11257), .ZN(n11261) );
  OR4D1BWP30P140LVT U11847 ( .A1(n11264), .A2(n11263), .A3(n11262), .A4(n11261), .Z(o_data_bus[43]) );
  AOI22D1BWP30P140LVT U11848 ( .A1(n11659), .A2(i_data_bus[940]), .B1(n11652), 
        .B2(i_data_bus[12]), .ZN(n11268) );
  AOI22D1BWP30P140LVT U11849 ( .A1(n11650), .A2(i_data_bus[556]), .B1(n11657), 
        .B2(i_data_bus[620]), .ZN(n11267) );
  AOI22D1BWP30P140LVT U11850 ( .A1(n11648), .A2(i_data_bus[44]), .B1(n11645), 
        .B2(i_data_bus[76]), .ZN(n11266) );
  AOI22D1BWP30P140LVT U11851 ( .A1(n11658), .A2(i_data_bus[524]), .B1(n11649), 
        .B2(i_data_bus[908]), .ZN(n11265) );
  ND4D1BWP30P140LVT U11852 ( .A1(n11268), .A2(n11267), .A3(n11266), .A4(n11265), .ZN(n11284) );
  AOI22D1BWP30P140LVT U11853 ( .A1(n11646), .A2(i_data_bus[1004]), .B1(n11651), 
        .B2(i_data_bus[588]), .ZN(n11272) );
  AOI22D1BWP30P140LVT U11854 ( .A1(n11660), .A2(i_data_bus[108]), .B1(n11647), 
        .B2(i_data_bus[972]), .ZN(n11271) );
  AOI22D1BWP30P140LVT U11855 ( .A1(n11670), .A2(i_data_bus[780]), .B1(n11686), 
        .B2(i_data_bus[460]), .ZN(n11270) );
  AOI22D1BWP30P140LVT U11856 ( .A1(n11669), .A2(i_data_bus[716]), .B1(n11661), 
        .B2(i_data_bus[300]), .ZN(n11269) );
  ND4D1BWP30P140LVT U11857 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(n11283) );
  AOI22D1BWP30P140LVT U11858 ( .A1(n11685), .A2(i_data_bus[364]), .B1(n11683), 
        .B2(i_data_bus[684]), .ZN(n11276) );
  AOI22D1BWP30P140LVT U11859 ( .A1(n11662), .A2(i_data_bus[428]), .B1(n11663), 
        .B2(i_data_bus[268]), .ZN(n11275) );
  AOI22D1BWP30P140LVT U11860 ( .A1(n11671), .A2(i_data_bus[748]), .B1(n11682), 
        .B2(i_data_bus[140]), .ZN(n11274) );
  AOI22D1BWP30P140LVT U11861 ( .A1(n11675), .A2(i_data_bus[204]), .B1(n11673), 
        .B2(i_data_bus[812]), .ZN(n11273) );
  ND4D1BWP30P140LVT U11862 ( .A1(n11276), .A2(n11275), .A3(n11274), .A4(n11273), .ZN(n11282) );
  AOI22D1BWP30P140LVT U11863 ( .A1(n11674), .A2(i_data_bus[396]), .B1(n11688), 
        .B2(i_data_bus[236]), .ZN(n11280) );
  AOI22D1BWP30P140LVT U11864 ( .A1(n11664), .A2(i_data_bus[492]), .B1(n11676), 
        .B2(i_data_bus[844]), .ZN(n11279) );
  AOI22D1BWP30P140LVT U11865 ( .A1(n11672), .A2(i_data_bus[652]), .B1(n11681), 
        .B2(i_data_bus[876]), .ZN(n11278) );
  AOI22D1BWP30P140LVT U11866 ( .A1(n11684), .A2(i_data_bus[172]), .B1(n11687), 
        .B2(i_data_bus[332]), .ZN(n11277) );
  ND4D1BWP30P140LVT U11867 ( .A1(n11280), .A2(n11279), .A3(n11278), .A4(n11277), .ZN(n11281) );
  OR4D1BWP30P140LVT U11868 ( .A1(n11284), .A2(n11283), .A3(n11282), .A4(n11281), .Z(o_data_bus[44]) );
  AOI22D1BWP30P140LVT U11869 ( .A1(n11648), .A2(i_data_bus[45]), .B1(n11658), 
        .B2(i_data_bus[525]), .ZN(n11288) );
  AOI22D1BWP30P140LVT U11870 ( .A1(n11649), .A2(i_data_bus[909]), .B1(n11657), 
        .B2(i_data_bus[621]), .ZN(n11287) );
  AOI22D1BWP30P140LVT U11871 ( .A1(n11650), .A2(i_data_bus[557]), .B1(n11647), 
        .B2(i_data_bus[973]), .ZN(n11286) );
  AOI22D1BWP30P140LVT U11872 ( .A1(n11646), .A2(i_data_bus[1005]), .B1(n11651), 
        .B2(i_data_bus[589]), .ZN(n11285) );
  ND4D1BWP30P140LVT U11873 ( .A1(n11288), .A2(n11287), .A3(n11286), .A4(n11285), .ZN(n11304) );
  AOI22D1BWP30P140LVT U11874 ( .A1(n11660), .A2(i_data_bus[109]), .B1(n11645), 
        .B2(i_data_bus[77]), .ZN(n11292) );
  AOI22D1BWP30P140LVT U11875 ( .A1(n11659), .A2(i_data_bus[941]), .B1(n11652), 
        .B2(i_data_bus[13]), .ZN(n11291) );
  AOI22D1BWP30P140LVT U11876 ( .A1(n11674), .A2(i_data_bus[397]), .B1(n11688), 
        .B2(i_data_bus[237]), .ZN(n11290) );
  AOI22D1BWP30P140LVT U11877 ( .A1(n11685), .A2(i_data_bus[365]), .B1(n11663), 
        .B2(i_data_bus[269]), .ZN(n11289) );
  ND4D1BWP30P140LVT U11878 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(n11303) );
  AOI22D1BWP30P140LVT U11879 ( .A1(n11664), .A2(i_data_bus[493]), .B1(n11662), 
        .B2(i_data_bus[429]), .ZN(n11296) );
  AOI22D1BWP30P140LVT U11880 ( .A1(n11682), .A2(i_data_bus[141]), .B1(n11681), 
        .B2(i_data_bus[877]), .ZN(n11295) );
  AOI22D1BWP30P140LVT U11881 ( .A1(n11671), .A2(i_data_bus[749]), .B1(n11670), 
        .B2(i_data_bus[781]), .ZN(n11294) );
  AOI22D1BWP30P140LVT U11882 ( .A1(n11675), .A2(i_data_bus[205]), .B1(n11661), 
        .B2(i_data_bus[301]), .ZN(n11293) );
  ND4D1BWP30P140LVT U11883 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(n11302) );
  AOI22D1BWP30P140LVT U11884 ( .A1(n11676), .A2(i_data_bus[845]), .B1(n11683), 
        .B2(i_data_bus[685]), .ZN(n11300) );
  AOI22D1BWP30P140LVT U11885 ( .A1(n11672), .A2(i_data_bus[653]), .B1(n11687), 
        .B2(i_data_bus[333]), .ZN(n11299) );
  AOI22D1BWP30P140LVT U11886 ( .A1(n11684), .A2(i_data_bus[173]), .B1(n11673), 
        .B2(i_data_bus[813]), .ZN(n11298) );
  AOI22D1BWP30P140LVT U11887 ( .A1(n11686), .A2(i_data_bus[461]), .B1(n11669), 
        .B2(i_data_bus[717]), .ZN(n11297) );
  ND4D1BWP30P140LVT U11888 ( .A1(n11300), .A2(n11299), .A3(n11298), .A4(n11297), .ZN(n11301) );
  OR4D1BWP30P140LVT U11889 ( .A1(n11304), .A2(n11303), .A3(n11302), .A4(n11301), .Z(o_data_bus[45]) );
  AOI22D1BWP30P140LVT U11890 ( .A1(n11660), .A2(i_data_bus[110]), .B1(n11649), 
        .B2(i_data_bus[910]), .ZN(n11308) );
  AOI22D1BWP30P140LVT U11891 ( .A1(n11646), .A2(i_data_bus[1006]), .B1(n11645), 
        .B2(i_data_bus[78]), .ZN(n11307) );
  AOI22D1BWP30P140LVT U11892 ( .A1(n11652), .A2(i_data_bus[14]), .B1(n11651), 
        .B2(i_data_bus[590]), .ZN(n11306) );
  AOI22D1BWP30P140LVT U11893 ( .A1(n11648), .A2(i_data_bus[46]), .B1(n11650), 
        .B2(i_data_bus[558]), .ZN(n11305) );
  ND4D1BWP30P140LVT U11894 ( .A1(n11308), .A2(n11307), .A3(n11306), .A4(n11305), .ZN(n11324) );
  AOI22D1BWP30P140LVT U11895 ( .A1(n11659), .A2(i_data_bus[942]), .B1(n11647), 
        .B2(i_data_bus[974]), .ZN(n11312) );
  AOI22D1BWP30P140LVT U11896 ( .A1(n11658), .A2(i_data_bus[526]), .B1(n11657), 
        .B2(i_data_bus[622]), .ZN(n11311) );
  AOI22D1BWP30P140LVT U11897 ( .A1(n11684), .A2(i_data_bus[174]), .B1(n11663), 
        .B2(i_data_bus[270]), .ZN(n11310) );
  AOI22D1BWP30P140LVT U11898 ( .A1(n11685), .A2(i_data_bus[366]), .B1(n11675), 
        .B2(i_data_bus[206]), .ZN(n11309) );
  ND4D1BWP30P140LVT U11899 ( .A1(n11312), .A2(n11311), .A3(n11310), .A4(n11309), .ZN(n11323) );
  AOI22D1BWP30P140LVT U11900 ( .A1(n11686), .A2(i_data_bus[462]), .B1(n11688), 
        .B2(i_data_bus[238]), .ZN(n11316) );
  AOI22D1BWP30P140LVT U11901 ( .A1(n11682), .A2(i_data_bus[142]), .B1(n11673), 
        .B2(i_data_bus[814]), .ZN(n11315) );
  AOI22D1BWP30P140LVT U11902 ( .A1(n11676), .A2(i_data_bus[846]), .B1(n11661), 
        .B2(i_data_bus[302]), .ZN(n11314) );
  AOI22D1BWP30P140LVT U11903 ( .A1(n11670), .A2(i_data_bus[782]), .B1(n11687), 
        .B2(i_data_bus[334]), .ZN(n11313) );
  ND4D1BWP30P140LVT U11904 ( .A1(n11316), .A2(n11315), .A3(n11314), .A4(n11313), .ZN(n11322) );
  AOI22D1BWP30P140LVT U11905 ( .A1(n11683), .A2(i_data_bus[686]), .B1(n11681), 
        .B2(i_data_bus[878]), .ZN(n11320) );
  AOI22D1BWP30P140LVT U11906 ( .A1(n11674), .A2(i_data_bus[398]), .B1(n11662), 
        .B2(i_data_bus[430]), .ZN(n11319) );
  AOI22D1BWP30P140LVT U11907 ( .A1(n11664), .A2(i_data_bus[494]), .B1(n11671), 
        .B2(i_data_bus[750]), .ZN(n11318) );
  AOI22D1BWP30P140LVT U11908 ( .A1(n11672), .A2(i_data_bus[654]), .B1(n11669), 
        .B2(i_data_bus[718]), .ZN(n11317) );
  ND4D1BWP30P140LVT U11909 ( .A1(n11320), .A2(n11319), .A3(n11318), .A4(n11317), .ZN(n11321) );
  OR4D1BWP30P140LVT U11910 ( .A1(n11324), .A2(n11323), .A3(n11322), .A4(n11321), .Z(o_data_bus[46]) );
  AOI22D1BWP30P140LVT U11911 ( .A1(n11645), .A2(i_data_bus[79]), .B1(n11647), 
        .B2(i_data_bus[975]), .ZN(n11328) );
  AOI22D1BWP30P140LVT U11912 ( .A1(n11651), .A2(i_data_bus[591]), .B1(n11649), 
        .B2(i_data_bus[911]), .ZN(n11327) );
  AOI22D1BWP30P140LVT U11913 ( .A1(n11650), .A2(i_data_bus[559]), .B1(n11660), 
        .B2(i_data_bus[111]), .ZN(n11326) );
  AOI22D1BWP30P140LVT U11914 ( .A1(n11648), .A2(i_data_bus[47]), .B1(n11658), 
        .B2(i_data_bus[527]), .ZN(n11325) );
  ND4D1BWP30P140LVT U11915 ( .A1(n11328), .A2(n11327), .A3(n11326), .A4(n11325), .ZN(n11344) );
  AOI22D1BWP30P140LVT U11916 ( .A1(n11652), .A2(i_data_bus[15]), .B1(n11657), 
        .B2(i_data_bus[623]), .ZN(n11332) );
  AOI22D1BWP30P140LVT U11917 ( .A1(n11646), .A2(i_data_bus[1007]), .B1(n11659), 
        .B2(i_data_bus[943]), .ZN(n11331) );
  AOI22D1BWP30P140LVT U11918 ( .A1(n11671), .A2(i_data_bus[751]), .B1(n11669), 
        .B2(i_data_bus[719]), .ZN(n11330) );
  AOI22D1BWP30P140LVT U11919 ( .A1(n11676), .A2(i_data_bus[847]), .B1(n11663), 
        .B2(i_data_bus[271]), .ZN(n11329) );
  ND4D1BWP30P140LVT U11920 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(n11343) );
  AOI22D1BWP30P140LVT U11921 ( .A1(n11662), .A2(i_data_bus[431]), .B1(n11675), 
        .B2(i_data_bus[207]), .ZN(n11336) );
  AOI22D1BWP30P140LVT U11922 ( .A1(n11684), .A2(i_data_bus[175]), .B1(n11688), 
        .B2(i_data_bus[239]), .ZN(n11335) );
  AOI22D1BWP30P140LVT U11923 ( .A1(n11664), .A2(i_data_bus[495]), .B1(n11682), 
        .B2(i_data_bus[143]), .ZN(n11334) );
  AOI22D1BWP30P140LVT U11924 ( .A1(n11672), .A2(i_data_bus[655]), .B1(n11686), 
        .B2(i_data_bus[463]), .ZN(n11333) );
  ND4D1BWP30P140LVT U11925 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(n11342) );
  AOI22D1BWP30P140LVT U11926 ( .A1(n11670), .A2(i_data_bus[783]), .B1(n11681), 
        .B2(i_data_bus[879]), .ZN(n11340) );
  AOI22D1BWP30P140LVT U11927 ( .A1(n11674), .A2(i_data_bus[399]), .B1(n11673), 
        .B2(i_data_bus[815]), .ZN(n11339) );
  AOI22D1BWP30P140LVT U11928 ( .A1(n11683), .A2(i_data_bus[687]), .B1(n11687), 
        .B2(i_data_bus[335]), .ZN(n11338) );
  AOI22D1BWP30P140LVT U11929 ( .A1(n11685), .A2(i_data_bus[367]), .B1(n11661), 
        .B2(i_data_bus[303]), .ZN(n11337) );
  ND4D1BWP30P140LVT U11930 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(n11341) );
  OR4D1BWP30P140LVT U11931 ( .A1(n11344), .A2(n11343), .A3(n11342), .A4(n11341), .Z(o_data_bus[47]) );
  AOI22D1BWP30P140LVT U11932 ( .A1(n11650), .A2(i_data_bus[560]), .B1(n11659), 
        .B2(i_data_bus[944]), .ZN(n11348) );
  AOI22D1BWP30P140LVT U11933 ( .A1(n11648), .A2(i_data_bus[48]), .B1(n11645), 
        .B2(i_data_bus[80]), .ZN(n11347) );
  AOI22D1BWP30P140LVT U11934 ( .A1(n11658), .A2(i_data_bus[528]), .B1(n11657), 
        .B2(i_data_bus[624]), .ZN(n11346) );
  AOI22D1BWP30P140LVT U11935 ( .A1(n11647), .A2(i_data_bus[976]), .B1(n11649), 
        .B2(i_data_bus[912]), .ZN(n11345) );
  ND4D1BWP30P140LVT U11936 ( .A1(n11348), .A2(n11347), .A3(n11346), .A4(n11345), .ZN(n11364) );
  AOI22D1BWP30P140LVT U11937 ( .A1(n11660), .A2(i_data_bus[112]), .B1(n11651), 
        .B2(i_data_bus[592]), .ZN(n11352) );
  AOI22D1BWP30P140LVT U11938 ( .A1(n11646), .A2(i_data_bus[1008]), .B1(n11652), 
        .B2(i_data_bus[16]), .ZN(n11351) );
  AOI22D1BWP30P140LVT U11939 ( .A1(n11662), .A2(i_data_bus[432]), .B1(n11661), 
        .B2(i_data_bus[304]), .ZN(n11350) );
  AOI22D1BWP30P140LVT U11940 ( .A1(n11664), .A2(i_data_bus[496]), .B1(n11687), 
        .B2(i_data_bus[336]), .ZN(n11349) );
  ND4D1BWP30P140LVT U11941 ( .A1(n11352), .A2(n11351), .A3(n11350), .A4(n11349), .ZN(n11363) );
  AOI22D1BWP30P140LVT U11942 ( .A1(n11682), .A2(i_data_bus[144]), .B1(n11681), 
        .B2(i_data_bus[880]), .ZN(n11356) );
  AOI22D1BWP30P140LVT U11943 ( .A1(n11672), .A2(i_data_bus[656]), .B1(n11670), 
        .B2(i_data_bus[784]), .ZN(n11355) );
  AOI22D1BWP30P140LVT U11944 ( .A1(n11671), .A2(i_data_bus[752]), .B1(n11669), 
        .B2(i_data_bus[720]), .ZN(n11354) );
  AOI22D1BWP30P140LVT U11945 ( .A1(n11675), .A2(i_data_bus[208]), .B1(n11673), 
        .B2(i_data_bus[816]), .ZN(n11353) );
  ND4D1BWP30P140LVT U11946 ( .A1(n11356), .A2(n11355), .A3(n11354), .A4(n11353), .ZN(n11362) );
  AOI22D1BWP30P140LVT U11947 ( .A1(n11686), .A2(i_data_bus[464]), .B1(n11663), 
        .B2(i_data_bus[272]), .ZN(n11360) );
  AOI22D1BWP30P140LVT U11948 ( .A1(n11684), .A2(i_data_bus[176]), .B1(n11685), 
        .B2(i_data_bus[368]), .ZN(n11359) );
  AOI22D1BWP30P140LVT U11949 ( .A1(n11674), .A2(i_data_bus[400]), .B1(n11688), 
        .B2(i_data_bus[240]), .ZN(n11358) );
  AOI22D1BWP30P140LVT U11950 ( .A1(n11676), .A2(i_data_bus[848]), .B1(n11683), 
        .B2(i_data_bus[688]), .ZN(n11357) );
  ND4D1BWP30P140LVT U11951 ( .A1(n11360), .A2(n11359), .A3(n11358), .A4(n11357), .ZN(n11361) );
  OR4D1BWP30P140LVT U11952 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .Z(o_data_bus[48]) );
  AOI22D1BWP30P140LVT U11953 ( .A1(n11652), .A2(i_data_bus[17]), .B1(n11657), 
        .B2(i_data_bus[625]), .ZN(n11368) );
  AOI22D1BWP30P140LVT U11954 ( .A1(n11646), .A2(i_data_bus[1009]), .B1(n11648), 
        .B2(i_data_bus[49]), .ZN(n11367) );
  AOI22D1BWP30P140LVT U11955 ( .A1(n11645), .A2(i_data_bus[81]), .B1(n11649), 
        .B2(i_data_bus[913]), .ZN(n11366) );
  AOI22D1BWP30P140LVT U11956 ( .A1(n11659), .A2(i_data_bus[945]), .B1(n11651), 
        .B2(i_data_bus[593]), .ZN(n11365) );
  ND4D1BWP30P140LVT U11957 ( .A1(n11368), .A2(n11367), .A3(n11366), .A4(n11365), .ZN(n11384) );
  AOI22D1BWP30P140LVT U11958 ( .A1(n11660), .A2(i_data_bus[113]), .B1(n11647), 
        .B2(i_data_bus[977]), .ZN(n11372) );
  AOI22D1BWP30P140LVT U11959 ( .A1(n11650), .A2(i_data_bus[561]), .B1(n11658), 
        .B2(i_data_bus[529]), .ZN(n11371) );
  AOI22D1BWP30P140LVT U11960 ( .A1(n11683), .A2(i_data_bus[689]), .B1(n11681), 
        .B2(i_data_bus[881]), .ZN(n11370) );
  AOI22D1BWP30P140LVT U11961 ( .A1(n11662), .A2(i_data_bus[433]), .B1(n11676), 
        .B2(i_data_bus[849]), .ZN(n11369) );
  ND4D1BWP30P140LVT U11962 ( .A1(n11372), .A2(n11371), .A3(n11370), .A4(n11369), .ZN(n11383) );
  AOI22D1BWP30P140LVT U11963 ( .A1(n11682), .A2(i_data_bus[145]), .B1(n11687), 
        .B2(i_data_bus[337]), .ZN(n11376) );
  AOI22D1BWP30P140LVT U11964 ( .A1(n11674), .A2(i_data_bus[401]), .B1(n11688), 
        .B2(i_data_bus[241]), .ZN(n11375) );
  AOI22D1BWP30P140LVT U11965 ( .A1(n11670), .A2(i_data_bus[785]), .B1(n11675), 
        .B2(i_data_bus[209]), .ZN(n11374) );
  AOI22D1BWP30P140LVT U11966 ( .A1(n11669), .A2(i_data_bus[721]), .B1(n11663), 
        .B2(i_data_bus[273]), .ZN(n11373) );
  ND4D1BWP30P140LVT U11967 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(n11382) );
  AOI22D1BWP30P140LVT U11968 ( .A1(n11684), .A2(i_data_bus[177]), .B1(n11661), 
        .B2(i_data_bus[305]), .ZN(n11380) );
  AOI22D1BWP30P140LVT U11969 ( .A1(n11672), .A2(i_data_bus[657]), .B1(n11671), 
        .B2(i_data_bus[753]), .ZN(n11379) );
  AOI22D1BWP30P140LVT U11970 ( .A1(n11664), .A2(i_data_bus[497]), .B1(n11686), 
        .B2(i_data_bus[465]), .ZN(n11378) );
  AOI22D1BWP30P140LVT U11971 ( .A1(n11685), .A2(i_data_bus[369]), .B1(n11673), 
        .B2(i_data_bus[817]), .ZN(n11377) );
  ND4D1BWP30P140LVT U11972 ( .A1(n11380), .A2(n11379), .A3(n11378), .A4(n11377), .ZN(n11381) );
  OR4D1BWP30P140LVT U11973 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .Z(o_data_bus[49]) );
  AOI22D1BWP30P140LVT U11974 ( .A1(n11651), .A2(i_data_bus[594]), .B1(n11657), 
        .B2(i_data_bus[626]), .ZN(n11388) );
  AOI22D1BWP30P140LVT U11975 ( .A1(n11648), .A2(i_data_bus[50]), .B1(n11647), 
        .B2(i_data_bus[978]), .ZN(n11387) );
  AOI22D1BWP30P140LVT U11976 ( .A1(n11660), .A2(i_data_bus[114]), .B1(n11658), 
        .B2(i_data_bus[530]), .ZN(n11386) );
  AOI22D1BWP30P140LVT U11977 ( .A1(n11646), .A2(i_data_bus[1010]), .B1(n11650), 
        .B2(i_data_bus[562]), .ZN(n11385) );
  ND4D1BWP30P140LVT U11978 ( .A1(n11388), .A2(n11387), .A3(n11386), .A4(n11385), .ZN(n11404) );
  AOI22D1BWP30P140LVT U11979 ( .A1(n11645), .A2(i_data_bus[82]), .B1(n11649), 
        .B2(i_data_bus[914]), .ZN(n11392) );
  AOI22D1BWP30P140LVT U11980 ( .A1(n11659), .A2(i_data_bus[946]), .B1(n11652), 
        .B2(i_data_bus[18]), .ZN(n11391) );
  AOI22D1BWP30P140LVT U11981 ( .A1(n11669), .A2(i_data_bus[722]), .B1(n11681), 
        .B2(i_data_bus[882]), .ZN(n11390) );
  AOI22D1BWP30P140LVT U11982 ( .A1(n11674), .A2(i_data_bus[402]), .B1(n11688), 
        .B2(i_data_bus[242]), .ZN(n11389) );
  ND4D1BWP30P140LVT U11983 ( .A1(n11392), .A2(n11391), .A3(n11390), .A4(n11389), .ZN(n11403) );
  AOI22D1BWP30P140LVT U11984 ( .A1(n11675), .A2(i_data_bus[210]), .B1(n11673), 
        .B2(i_data_bus[818]), .ZN(n11396) );
  AOI22D1BWP30P140LVT U11985 ( .A1(n11685), .A2(i_data_bus[370]), .B1(n11683), 
        .B2(i_data_bus[690]), .ZN(n11395) );
  AOI22D1BWP30P140LVT U11986 ( .A1(n11664), .A2(i_data_bus[498]), .B1(n11684), 
        .B2(i_data_bus[178]), .ZN(n11394) );
  AOI22D1BWP30P140LVT U11987 ( .A1(n11676), .A2(i_data_bus[850]), .B1(n11661), 
        .B2(i_data_bus[306]), .ZN(n11393) );
  ND4D1BWP30P140LVT U11988 ( .A1(n11396), .A2(n11395), .A3(n11394), .A4(n11393), .ZN(n11402) );
  AOI22D1BWP30P140LVT U11989 ( .A1(n11672), .A2(i_data_bus[658]), .B1(n11686), 
        .B2(i_data_bus[466]), .ZN(n11400) );
  AOI22D1BWP30P140LVT U11990 ( .A1(n11682), .A2(i_data_bus[146]), .B1(n11663), 
        .B2(i_data_bus[274]), .ZN(n11399) );
  AOI22D1BWP30P140LVT U11991 ( .A1(n11671), .A2(i_data_bus[754]), .B1(n11670), 
        .B2(i_data_bus[786]), .ZN(n11398) );
  AOI22D1BWP30P140LVT U11992 ( .A1(n11662), .A2(i_data_bus[434]), .B1(n11687), 
        .B2(i_data_bus[338]), .ZN(n11397) );
  ND4D1BWP30P140LVT U11993 ( .A1(n11400), .A2(n11399), .A3(n11398), .A4(n11397), .ZN(n11401) );
  OR4D1BWP30P140LVT U11994 ( .A1(n11404), .A2(n11403), .A3(n11402), .A4(n11401), .Z(o_data_bus[50]) );
  AOI22D1BWP30P140LVT U11995 ( .A1(n11650), .A2(i_data_bus[563]), .B1(n11647), 
        .B2(i_data_bus[979]), .ZN(n11408) );
  AOI22D1BWP30P140LVT U11996 ( .A1(n11648), .A2(i_data_bus[51]), .B1(n11658), 
        .B2(i_data_bus[531]), .ZN(n11407) );
  AOI22D1BWP30P140LVT U11997 ( .A1(n11646), .A2(i_data_bus[1011]), .B1(n11660), 
        .B2(i_data_bus[115]), .ZN(n11406) );
  AOI22D1BWP30P140LVT U11998 ( .A1(n11659), .A2(i_data_bus[947]), .B1(n11645), 
        .B2(i_data_bus[83]), .ZN(n11405) );
  ND4D1BWP30P140LVT U11999 ( .A1(n11408), .A2(n11407), .A3(n11406), .A4(n11405), .ZN(n11424) );
  AOI22D1BWP30P140LVT U12000 ( .A1(n11652), .A2(i_data_bus[19]), .B1(n11649), 
        .B2(i_data_bus[915]), .ZN(n11412) );
  AOI22D1BWP30P140LVT U12001 ( .A1(n11651), .A2(i_data_bus[595]), .B1(n11657), 
        .B2(i_data_bus[627]), .ZN(n11411) );
  AOI22D1BWP30P140LVT U12002 ( .A1(n11671), .A2(i_data_bus[755]), .B1(n11685), 
        .B2(i_data_bus[371]), .ZN(n11410) );
  AOI22D1BWP30P140LVT U12003 ( .A1(n11684), .A2(i_data_bus[179]), .B1(n11675), 
        .B2(i_data_bus[211]), .ZN(n11409) );
  ND4D1BWP30P140LVT U12004 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(n11423) );
  AOI22D1BWP30P140LVT U12005 ( .A1(n11674), .A2(i_data_bus[403]), .B1(n11661), 
        .B2(i_data_bus[307]), .ZN(n11416) );
  AOI22D1BWP30P140LVT U12006 ( .A1(n11682), .A2(i_data_bus[147]), .B1(n11687), 
        .B2(i_data_bus[339]), .ZN(n11415) );
  AOI22D1BWP30P140LVT U12007 ( .A1(n11688), .A2(i_data_bus[243]), .B1(n11673), 
        .B2(i_data_bus[819]), .ZN(n11414) );
  AOI22D1BWP30P140LVT U12008 ( .A1(n11672), .A2(i_data_bus[659]), .B1(n11670), 
        .B2(i_data_bus[787]), .ZN(n11413) );
  ND4D1BWP30P140LVT U12009 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(n11422) );
  AOI22D1BWP30P140LVT U12010 ( .A1(n11676), .A2(i_data_bus[851]), .B1(n11681), 
        .B2(i_data_bus[883]), .ZN(n11420) );
  AOI22D1BWP30P140LVT U12011 ( .A1(n11664), .A2(i_data_bus[499]), .B1(n11683), 
        .B2(i_data_bus[691]), .ZN(n11419) );
  AOI22D1BWP30P140LVT U12012 ( .A1(n11662), .A2(i_data_bus[435]), .B1(n11669), 
        .B2(i_data_bus[723]), .ZN(n11418) );
  AOI22D1BWP30P140LVT U12013 ( .A1(n11686), .A2(i_data_bus[467]), .B1(n11663), 
        .B2(i_data_bus[275]), .ZN(n11417) );
  ND4D1BWP30P140LVT U12014 ( .A1(n11420), .A2(n11419), .A3(n11418), .A4(n11417), .ZN(n11421) );
  OR4D1BWP30P140LVT U12015 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .Z(o_data_bus[51]) );
  AOI22D1BWP30P140LVT U12016 ( .A1(n11658), .A2(i_data_bus[532]), .B1(n11651), 
        .B2(i_data_bus[596]), .ZN(n11428) );
  AOI22D1BWP30P140LVT U12017 ( .A1(n11648), .A2(i_data_bus[52]), .B1(n11647), 
        .B2(i_data_bus[980]), .ZN(n11427) );
  AOI22D1BWP30P140LVT U12018 ( .A1(n11646), .A2(i_data_bus[1012]), .B1(n11650), 
        .B2(i_data_bus[564]), .ZN(n11426) );
  AOI22D1BWP30P140LVT U12019 ( .A1(n11652), .A2(i_data_bus[20]), .B1(n11657), 
        .B2(i_data_bus[628]), .ZN(n11425) );
  ND4D1BWP30P140LVT U12020 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(n11444) );
  AOI22D1BWP30P140LVT U12021 ( .A1(n11659), .A2(i_data_bus[948]), .B1(n11645), 
        .B2(i_data_bus[84]), .ZN(n11432) );
  AOI22D1BWP30P140LVT U12022 ( .A1(n11660), .A2(i_data_bus[116]), .B1(n11649), 
        .B2(i_data_bus[916]), .ZN(n11431) );
  AOI22D1BWP30P140LVT U12023 ( .A1(n11669), .A2(i_data_bus[724]), .B1(n11675), 
        .B2(i_data_bus[212]), .ZN(n11430) );
  AOI22D1BWP30P140LVT U12024 ( .A1(n11688), .A2(i_data_bus[244]), .B1(n11687), 
        .B2(i_data_bus[340]), .ZN(n11429) );
  ND4D1BWP30P140LVT U12025 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(n11443) );
  AOI22D1BWP30P140LVT U12026 ( .A1(n11684), .A2(i_data_bus[180]), .B1(n11673), 
        .B2(i_data_bus[820]), .ZN(n11436) );
  AOI22D1BWP30P140LVT U12027 ( .A1(n11676), .A2(i_data_bus[852]), .B1(n11670), 
        .B2(i_data_bus[788]), .ZN(n11435) );
  AOI22D1BWP30P140LVT U12028 ( .A1(n11671), .A2(i_data_bus[756]), .B1(n11663), 
        .B2(i_data_bus[276]), .ZN(n11434) );
  AOI22D1BWP30P140LVT U12029 ( .A1(n11672), .A2(i_data_bus[660]), .B1(n11681), 
        .B2(i_data_bus[884]), .ZN(n11433) );
  ND4D1BWP30P140LVT U12030 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(n11442) );
  AOI22D1BWP30P140LVT U12031 ( .A1(n11674), .A2(i_data_bus[404]), .B1(n11662), 
        .B2(i_data_bus[436]), .ZN(n11440) );
  AOI22D1BWP30P140LVT U12032 ( .A1(n11686), .A2(i_data_bus[468]), .B1(n11683), 
        .B2(i_data_bus[692]), .ZN(n11439) );
  AOI22D1BWP30P140LVT U12033 ( .A1(n11682), .A2(i_data_bus[148]), .B1(n11661), 
        .B2(i_data_bus[308]), .ZN(n11438) );
  AOI22D1BWP30P140LVT U12034 ( .A1(n11664), .A2(i_data_bus[500]), .B1(n11685), 
        .B2(i_data_bus[372]), .ZN(n11437) );
  ND4D1BWP30P140LVT U12035 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(n11441) );
  OR4D1BWP30P140LVT U12036 ( .A1(n11444), .A2(n11443), .A3(n11442), .A4(n11441), .Z(o_data_bus[52]) );
  AOI22D1BWP30P140LVT U12037 ( .A1(n11648), .A2(i_data_bus[53]), .B1(n11659), 
        .B2(i_data_bus[949]), .ZN(n11448) );
  AOI22D1BWP30P140LVT U12038 ( .A1(n11660), .A2(i_data_bus[117]), .B1(n11657), 
        .B2(i_data_bus[629]), .ZN(n11447) );
  AOI22D1BWP30P140LVT U12039 ( .A1(n11647), .A2(i_data_bus[981]), .B1(n11649), 
        .B2(i_data_bus[917]), .ZN(n11446) );
  AOI22D1BWP30P140LVT U12040 ( .A1(n11652), .A2(i_data_bus[21]), .B1(n11651), 
        .B2(i_data_bus[597]), .ZN(n11445) );
  ND4D1BWP30P140LVT U12041 ( .A1(n11448), .A2(n11447), .A3(n11446), .A4(n11445), .ZN(n11464) );
  AOI22D1BWP30P140LVT U12042 ( .A1(n11650), .A2(i_data_bus[565]), .B1(n11658), 
        .B2(i_data_bus[533]), .ZN(n11452) );
  AOI22D1BWP30P140LVT U12043 ( .A1(n11646), .A2(i_data_bus[1013]), .B1(n11645), 
        .B2(i_data_bus[85]), .ZN(n11451) );
  AOI22D1BWP30P140LVT U12044 ( .A1(n11672), .A2(i_data_bus[661]), .B1(n11671), 
        .B2(i_data_bus[757]), .ZN(n11450) );
  AOI22D1BWP30P140LVT U12045 ( .A1(n11676), .A2(i_data_bus[853]), .B1(n11687), 
        .B2(i_data_bus[341]), .ZN(n11449) );
  ND4D1BWP30P140LVT U12046 ( .A1(n11452), .A2(n11451), .A3(n11450), .A4(n11449), .ZN(n11463) );
  AOI22D1BWP30P140LVT U12047 ( .A1(n11670), .A2(i_data_bus[789]), .B1(n11682), 
        .B2(i_data_bus[149]), .ZN(n11456) );
  AOI22D1BWP30P140LVT U12048 ( .A1(n11684), .A2(i_data_bus[181]), .B1(n11673), 
        .B2(i_data_bus[821]), .ZN(n11455) );
  AOI22D1BWP30P140LVT U12049 ( .A1(n11664), .A2(i_data_bus[501]), .B1(n11662), 
        .B2(i_data_bus[437]), .ZN(n11454) );
  AOI22D1BWP30P140LVT U12050 ( .A1(n11669), .A2(i_data_bus[725]), .B1(n11675), 
        .B2(i_data_bus[213]), .ZN(n11453) );
  ND4D1BWP30P140LVT U12051 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(n11462) );
  AOI22D1BWP30P140LVT U12052 ( .A1(n11683), .A2(i_data_bus[693]), .B1(n11661), 
        .B2(i_data_bus[309]), .ZN(n11460) );
  AOI22D1BWP30P140LVT U12053 ( .A1(n11686), .A2(i_data_bus[469]), .B1(n11688), 
        .B2(i_data_bus[245]), .ZN(n11459) );
  AOI22D1BWP30P140LVT U12054 ( .A1(n11674), .A2(i_data_bus[405]), .B1(n11663), 
        .B2(i_data_bus[277]), .ZN(n11458) );
  AOI22D1BWP30P140LVT U12055 ( .A1(n11685), .A2(i_data_bus[373]), .B1(n11681), 
        .B2(i_data_bus[885]), .ZN(n11457) );
  ND4D1BWP30P140LVT U12056 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(n11461) );
  OR4D1BWP30P140LVT U12057 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .Z(o_data_bus[53]) );
  AOI22D1BWP30P140LVT U12058 ( .A1(n11646), .A2(i_data_bus[1014]), .B1(n11648), 
        .B2(i_data_bus[54]), .ZN(n11468) );
  AOI22D1BWP30P140LVT U12059 ( .A1(n11650), .A2(i_data_bus[566]), .B1(n11658), 
        .B2(i_data_bus[534]), .ZN(n11467) );
  AOI22D1BWP30P140LVT U12060 ( .A1(n11660), .A2(i_data_bus[118]), .B1(n11651), 
        .B2(i_data_bus[598]), .ZN(n11466) );
  AOI22D1BWP30P140LVT U12061 ( .A1(n11659), .A2(i_data_bus[950]), .B1(n11649), 
        .B2(i_data_bus[918]), .ZN(n11465) );
  ND4D1BWP30P140LVT U12062 ( .A1(n11468), .A2(n11467), .A3(n11466), .A4(n11465), .ZN(n11484) );
  AOI22D1BWP30P140LVT U12063 ( .A1(n11652), .A2(i_data_bus[22]), .B1(n11645), 
        .B2(i_data_bus[86]), .ZN(n11472) );
  AOI22D1BWP30P140LVT U12064 ( .A1(n11647), .A2(i_data_bus[982]), .B1(n11657), 
        .B2(i_data_bus[630]), .ZN(n11471) );
  AOI22D1BWP30P140LVT U12065 ( .A1(n11683), .A2(i_data_bus[694]), .B1(n11673), 
        .B2(i_data_bus[822]), .ZN(n11470) );
  AOI22D1BWP30P140LVT U12066 ( .A1(n11662), .A2(i_data_bus[438]), .B1(n11671), 
        .B2(i_data_bus[758]), .ZN(n11469) );
  ND4D1BWP30P140LVT U12067 ( .A1(n11472), .A2(n11471), .A3(n11470), .A4(n11469), .ZN(n11483) );
  AOI22D1BWP30P140LVT U12068 ( .A1(n11670), .A2(i_data_bus[790]), .B1(n11688), 
        .B2(i_data_bus[246]), .ZN(n11476) );
  AOI22D1BWP30P140LVT U12069 ( .A1(n11674), .A2(i_data_bus[406]), .B1(n11685), 
        .B2(i_data_bus[374]), .ZN(n11475) );
  AOI22D1BWP30P140LVT U12070 ( .A1(n11664), .A2(i_data_bus[502]), .B1(n11684), 
        .B2(i_data_bus[182]), .ZN(n11474) );
  AOI22D1BWP30P140LVT U12071 ( .A1(n11682), .A2(i_data_bus[150]), .B1(n11669), 
        .B2(i_data_bus[726]), .ZN(n11473) );
  ND4D1BWP30P140LVT U12072 ( .A1(n11476), .A2(n11475), .A3(n11474), .A4(n11473), .ZN(n11482) );
  AOI22D1BWP30P140LVT U12073 ( .A1(n11681), .A2(i_data_bus[886]), .B1(n11661), 
        .B2(i_data_bus[310]), .ZN(n11480) );
  AOI22D1BWP30P140LVT U12074 ( .A1(n11686), .A2(i_data_bus[470]), .B1(n11687), 
        .B2(i_data_bus[342]), .ZN(n11479) );
  AOI22D1BWP30P140LVT U12075 ( .A1(n11676), .A2(i_data_bus[854]), .B1(n11663), 
        .B2(i_data_bus[278]), .ZN(n11478) );
  AOI22D1BWP30P140LVT U12076 ( .A1(n11672), .A2(i_data_bus[662]), .B1(n11675), 
        .B2(i_data_bus[214]), .ZN(n11477) );
  ND4D1BWP30P140LVT U12077 ( .A1(n11480), .A2(n11479), .A3(n11478), .A4(n11477), .ZN(n11481) );
  OR4D1BWP30P140LVT U12078 ( .A1(n11484), .A2(n11483), .A3(n11482), .A4(n11481), .Z(o_data_bus[54]) );
  AOI22D1BWP30P140LVT U12079 ( .A1(n11652), .A2(i_data_bus[23]), .B1(n11657), 
        .B2(i_data_bus[631]), .ZN(n11488) );
  AOI22D1BWP30P140LVT U12080 ( .A1(n11646), .A2(i_data_bus[1015]), .B1(n11648), 
        .B2(i_data_bus[55]), .ZN(n11487) );
  AOI22D1BWP30P140LVT U12081 ( .A1(n11651), .A2(i_data_bus[599]), .B1(n11645), 
        .B2(i_data_bus[87]), .ZN(n11486) );
  AOI22D1BWP30P140LVT U12082 ( .A1(n11660), .A2(i_data_bus[119]), .B1(n11659), 
        .B2(i_data_bus[951]), .ZN(n11485) );
  ND4D1BWP30P140LVT U12083 ( .A1(n11488), .A2(n11487), .A3(n11486), .A4(n11485), .ZN(n11504) );
  AOI22D1BWP30P140LVT U12084 ( .A1(n11658), .A2(i_data_bus[535]), .B1(n11647), 
        .B2(i_data_bus[983]), .ZN(n11492) );
  AOI22D1BWP30P140LVT U12085 ( .A1(n11650), .A2(i_data_bus[567]), .B1(n11649), 
        .B2(i_data_bus[919]), .ZN(n11491) );
  AOI22D1BWP30P140LVT U12086 ( .A1(n11683), .A2(i_data_bus[695]), .B1(n11688), 
        .B2(i_data_bus[247]), .ZN(n11490) );
  AOI22D1BWP30P140LVT U12087 ( .A1(n11686), .A2(i_data_bus[471]), .B1(n11681), 
        .B2(i_data_bus[887]), .ZN(n11489) );
  ND4D1BWP30P140LVT U12088 ( .A1(n11492), .A2(n11491), .A3(n11490), .A4(n11489), .ZN(n11503) );
  AOI22D1BWP30P140LVT U12089 ( .A1(n11684), .A2(i_data_bus[183]), .B1(n11661), 
        .B2(i_data_bus[311]), .ZN(n11496) );
  AOI22D1BWP30P140LVT U12090 ( .A1(n11671), .A2(i_data_bus[759]), .B1(n11663), 
        .B2(i_data_bus[279]), .ZN(n11495) );
  AOI22D1BWP30P140LVT U12091 ( .A1(n11664), .A2(i_data_bus[503]), .B1(n11675), 
        .B2(i_data_bus[215]), .ZN(n11494) );
  AOI22D1BWP30P140LVT U12092 ( .A1(n11662), .A2(i_data_bus[439]), .B1(n11669), 
        .B2(i_data_bus[727]), .ZN(n11493) );
  ND4D1BWP30P140LVT U12093 ( .A1(n11496), .A2(n11495), .A3(n11494), .A4(n11493), .ZN(n11502) );
  AOI22D1BWP30P140LVT U12094 ( .A1(n11674), .A2(i_data_bus[407]), .B1(n11682), 
        .B2(i_data_bus[151]), .ZN(n11500) );
  AOI22D1BWP30P140LVT U12095 ( .A1(n11672), .A2(i_data_bus[663]), .B1(n11673), 
        .B2(i_data_bus[823]), .ZN(n11499) );
  AOI22D1BWP30P140LVT U12096 ( .A1(n11670), .A2(i_data_bus[791]), .B1(n11685), 
        .B2(i_data_bus[375]), .ZN(n11498) );
  AOI22D1BWP30P140LVT U12097 ( .A1(n11676), .A2(i_data_bus[855]), .B1(n11687), 
        .B2(i_data_bus[343]), .ZN(n11497) );
  ND4D1BWP30P140LVT U12098 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(n11501) );
  OR4D1BWP30P140LVT U12099 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .Z(o_data_bus[55]) );
  AOI22D1BWP30P140LVT U12100 ( .A1(n11647), .A2(i_data_bus[984]), .B1(n11657), 
        .B2(i_data_bus[632]), .ZN(n11508) );
  AOI22D1BWP30P140LVT U12101 ( .A1(n11660), .A2(i_data_bus[120]), .B1(n11645), 
        .B2(i_data_bus[88]), .ZN(n11507) );
  AOI22D1BWP30P140LVT U12102 ( .A1(n11646), .A2(i_data_bus[1016]), .B1(n11651), 
        .B2(i_data_bus[600]), .ZN(n11506) );
  AOI22D1BWP30P140LVT U12103 ( .A1(n11658), .A2(i_data_bus[536]), .B1(n11652), 
        .B2(i_data_bus[24]), .ZN(n11505) );
  ND4D1BWP30P140LVT U12104 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(n11524) );
  AOI22D1BWP30P140LVT U12105 ( .A1(n11648), .A2(i_data_bus[56]), .B1(n11659), 
        .B2(i_data_bus[952]), .ZN(n11512) );
  AOI22D1BWP30P140LVT U12106 ( .A1(n11650), .A2(i_data_bus[568]), .B1(n11649), 
        .B2(i_data_bus[920]), .ZN(n11511) );
  AOI22D1BWP30P140LVT U12107 ( .A1(n11670), .A2(i_data_bus[792]), .B1(n11663), 
        .B2(i_data_bus[280]), .ZN(n11510) );
  AOI22D1BWP30P140LVT U12108 ( .A1(n11683), .A2(i_data_bus[696]), .B1(n11688), 
        .B2(i_data_bus[248]), .ZN(n11509) );
  ND4D1BWP30P140LVT U12109 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(n11523) );
  AOI22D1BWP30P140LVT U12110 ( .A1(n11674), .A2(i_data_bus[408]), .B1(n11687), 
        .B2(i_data_bus[344]), .ZN(n11516) );
  AOI22D1BWP30P140LVT U12111 ( .A1(n11662), .A2(i_data_bus[440]), .B1(n11676), 
        .B2(i_data_bus[856]), .ZN(n11515) );
  AOI22D1BWP30P140LVT U12112 ( .A1(n11672), .A2(i_data_bus[664]), .B1(n11673), 
        .B2(i_data_bus[824]), .ZN(n11514) );
  AOI22D1BWP30P140LVT U12113 ( .A1(n11685), .A2(i_data_bus[376]), .B1(n11669), 
        .B2(i_data_bus[728]), .ZN(n11513) );
  ND4D1BWP30P140LVT U12114 ( .A1(n11516), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(n11522) );
  AOI22D1BWP30P140LVT U12115 ( .A1(n11682), .A2(i_data_bus[152]), .B1(n11681), 
        .B2(i_data_bus[888]), .ZN(n11520) );
  AOI22D1BWP30P140LVT U12116 ( .A1(n11684), .A2(i_data_bus[184]), .B1(n11686), 
        .B2(i_data_bus[472]), .ZN(n11519) );
  AOI22D1BWP30P140LVT U12117 ( .A1(n11664), .A2(i_data_bus[504]), .B1(n11675), 
        .B2(i_data_bus[216]), .ZN(n11518) );
  AOI22D1BWP30P140LVT U12118 ( .A1(n11671), .A2(i_data_bus[760]), .B1(n11661), 
        .B2(i_data_bus[312]), .ZN(n11517) );
  ND4D1BWP30P140LVT U12119 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(n11521) );
  OR4D1BWP30P140LVT U12120 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .Z(o_data_bus[56]) );
  AOI22D1BWP30P140LVT U12121 ( .A1(n11646), .A2(i_data_bus[1017]), .B1(n11648), 
        .B2(i_data_bus[57]), .ZN(n11528) );
  AOI22D1BWP30P140LVT U12122 ( .A1(n11650), .A2(i_data_bus[569]), .B1(n11649), 
        .B2(i_data_bus[921]), .ZN(n11527) );
  AOI22D1BWP30P140LVT U12123 ( .A1(n11651), .A2(i_data_bus[601]), .B1(n11657), 
        .B2(i_data_bus[633]), .ZN(n11526) );
  AOI22D1BWP30P140LVT U12124 ( .A1(n11660), .A2(i_data_bus[121]), .B1(n11658), 
        .B2(i_data_bus[537]), .ZN(n11525) );
  ND4D1BWP30P140LVT U12125 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(n11544) );
  AOI22D1BWP30P140LVT U12126 ( .A1(n11652), .A2(i_data_bus[25]), .B1(n11647), 
        .B2(i_data_bus[985]), .ZN(n11532) );
  AOI22D1BWP30P140LVT U12127 ( .A1(n11659), .A2(i_data_bus[953]), .B1(n11645), 
        .B2(i_data_bus[89]), .ZN(n11531) );
  AOI22D1BWP30P140LVT U12128 ( .A1(n11669), .A2(i_data_bus[729]), .B1(n11673), 
        .B2(i_data_bus[825]), .ZN(n11530) );
  AOI22D1BWP30P140LVT U12129 ( .A1(n11672), .A2(i_data_bus[665]), .B1(n11683), 
        .B2(i_data_bus[697]), .ZN(n11529) );
  ND4D1BWP30P140LVT U12130 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(n11543) );
  AOI22D1BWP30P140LVT U12131 ( .A1(n11684), .A2(i_data_bus[185]), .B1(n11687), 
        .B2(i_data_bus[345]), .ZN(n11536) );
  AOI22D1BWP30P140LVT U12132 ( .A1(n11670), .A2(i_data_bus[793]), .B1(n11685), 
        .B2(i_data_bus[377]), .ZN(n11535) );
  AOI22D1BWP30P140LVT U12133 ( .A1(n11671), .A2(i_data_bus[761]), .B1(n11686), 
        .B2(i_data_bus[473]), .ZN(n11534) );
  AOI22D1BWP30P140LVT U12134 ( .A1(n11682), .A2(i_data_bus[153]), .B1(n11663), 
        .B2(i_data_bus[281]), .ZN(n11533) );
  ND4D1BWP30P140LVT U12135 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(n11542) );
  AOI22D1BWP30P140LVT U12136 ( .A1(n11674), .A2(i_data_bus[409]), .B1(n11675), 
        .B2(i_data_bus[217]), .ZN(n11540) );
  AOI22D1BWP30P140LVT U12137 ( .A1(n11681), .A2(i_data_bus[889]), .B1(n11661), 
        .B2(i_data_bus[313]), .ZN(n11539) );
  AOI22D1BWP30P140LVT U12138 ( .A1(n11664), .A2(i_data_bus[505]), .B1(n11676), 
        .B2(i_data_bus[857]), .ZN(n11538) );
  AOI22D1BWP30P140LVT U12139 ( .A1(n11662), .A2(i_data_bus[441]), .B1(n11688), 
        .B2(i_data_bus[249]), .ZN(n11537) );
  ND4D1BWP30P140LVT U12140 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(n11541) );
  OR4D1BWP30P140LVT U12141 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .Z(o_data_bus[57]) );
  AOI22D1BWP30P140LVT U12142 ( .A1(n11660), .A2(i_data_bus[122]), .B1(n11651), 
        .B2(i_data_bus[602]), .ZN(n11548) );
  AOI22D1BWP30P140LVT U12143 ( .A1(n11646), .A2(i_data_bus[1018]), .B1(n11645), 
        .B2(i_data_bus[90]), .ZN(n11547) );
  AOI22D1BWP30P140LVT U12144 ( .A1(n11659), .A2(i_data_bus[954]), .B1(n11647), 
        .B2(i_data_bus[986]), .ZN(n11546) );
  AOI22D1BWP30P140LVT U12145 ( .A1(n11658), .A2(i_data_bus[538]), .B1(n11649), 
        .B2(i_data_bus[922]), .ZN(n11545) );
  ND4D1BWP30P140LVT U12146 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(n11564) );
  AOI22D1BWP30P140LVT U12147 ( .A1(n11650), .A2(i_data_bus[570]), .B1(n11657), 
        .B2(i_data_bus[634]), .ZN(n11552) );
  AOI22D1BWP30P140LVT U12148 ( .A1(n11648), .A2(i_data_bus[58]), .B1(n11652), 
        .B2(i_data_bus[26]), .ZN(n11551) );
  AOI22D1BWP30P140LVT U12149 ( .A1(n11662), .A2(i_data_bus[442]), .B1(n11675), 
        .B2(i_data_bus[218]), .ZN(n11550) );
  AOI22D1BWP30P140LVT U12150 ( .A1(n11681), .A2(i_data_bus[890]), .B1(n11673), 
        .B2(i_data_bus[826]), .ZN(n11549) );
  ND4D1BWP30P140LVT U12151 ( .A1(n11552), .A2(n11551), .A3(n11550), .A4(n11549), .ZN(n11563) );
  AOI22D1BWP30P140LVT U12152 ( .A1(n11676), .A2(i_data_bus[858]), .B1(n11661), 
        .B2(i_data_bus[314]), .ZN(n11556) );
  AOI22D1BWP30P140LVT U12153 ( .A1(n11683), .A2(i_data_bus[698]), .B1(n11687), 
        .B2(i_data_bus[346]), .ZN(n11555) );
  AOI22D1BWP30P140LVT U12154 ( .A1(n11684), .A2(i_data_bus[186]), .B1(n11663), 
        .B2(i_data_bus[282]), .ZN(n11554) );
  AOI22D1BWP30P140LVT U12155 ( .A1(n11671), .A2(i_data_bus[762]), .B1(n11670), 
        .B2(i_data_bus[794]), .ZN(n11553) );
  ND4D1BWP30P140LVT U12156 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(n11562) );
  AOI22D1BWP30P140LVT U12157 ( .A1(n11664), .A2(i_data_bus[506]), .B1(n11688), 
        .B2(i_data_bus[250]), .ZN(n11560) );
  AOI22D1BWP30P140LVT U12158 ( .A1(n11674), .A2(i_data_bus[410]), .B1(n11672), 
        .B2(i_data_bus[666]), .ZN(n11559) );
  AOI22D1BWP30P140LVT U12159 ( .A1(n11682), .A2(i_data_bus[154]), .B1(n11669), 
        .B2(i_data_bus[730]), .ZN(n11558) );
  AOI22D1BWP30P140LVT U12160 ( .A1(n11686), .A2(i_data_bus[474]), .B1(n11685), 
        .B2(i_data_bus[378]), .ZN(n11557) );
  ND4D1BWP30P140LVT U12161 ( .A1(n11560), .A2(n11559), .A3(n11558), .A4(n11557), .ZN(n11561) );
  OR4D1BWP30P140LVT U12162 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .Z(o_data_bus[58]) );
  AOI22D1BWP30P140LVT U12163 ( .A1(n11660), .A2(i_data_bus[123]), .B1(n11647), 
        .B2(i_data_bus[987]), .ZN(n11568) );
  AOI22D1BWP30P140LVT U12164 ( .A1(n11646), .A2(i_data_bus[1019]), .B1(n11650), 
        .B2(i_data_bus[571]), .ZN(n11567) );
  AOI22D1BWP30P140LVT U12165 ( .A1(n11658), .A2(i_data_bus[539]), .B1(n11651), 
        .B2(i_data_bus[603]), .ZN(n11566) );
  AOI22D1BWP30P140LVT U12166 ( .A1(n11645), .A2(i_data_bus[91]), .B1(n11657), 
        .B2(i_data_bus[635]), .ZN(n11565) );
  ND4D1BWP30P140LVT U12167 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(n11584) );
  AOI22D1BWP30P140LVT U12168 ( .A1(n11652), .A2(i_data_bus[27]), .B1(n11649), 
        .B2(i_data_bus[923]), .ZN(n11572) );
  AOI22D1BWP30P140LVT U12169 ( .A1(n11648), .A2(i_data_bus[59]), .B1(n11659), 
        .B2(i_data_bus[955]), .ZN(n11571) );
  AOI22D1BWP30P140LVT U12170 ( .A1(n11674), .A2(i_data_bus[411]), .B1(n11664), 
        .B2(i_data_bus[507]), .ZN(n11570) );
  AOI22D1BWP30P140LVT U12171 ( .A1(n11669), .A2(i_data_bus[731]), .B1(n11673), 
        .B2(i_data_bus[827]), .ZN(n11569) );
  ND4D1BWP30P140LVT U12172 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(n11583) );
  AOI22D1BWP30P140LVT U12173 ( .A1(n11662), .A2(i_data_bus[443]), .B1(n11682), 
        .B2(i_data_bus[155]), .ZN(n11576) );
  AOI22D1BWP30P140LVT U12174 ( .A1(n11681), .A2(i_data_bus[891]), .B1(n11661), 
        .B2(i_data_bus[315]), .ZN(n11575) );
  AOI22D1BWP30P140LVT U12175 ( .A1(n11685), .A2(i_data_bus[379]), .B1(n11675), 
        .B2(i_data_bus[219]), .ZN(n11574) );
  AOI22D1BWP30P140LVT U12176 ( .A1(n11688), .A2(i_data_bus[251]), .B1(n11663), 
        .B2(i_data_bus[283]), .ZN(n11573) );
  ND4D1BWP30P140LVT U12177 ( .A1(n11576), .A2(n11575), .A3(n11574), .A4(n11573), .ZN(n11582) );
  AOI22D1BWP30P140LVT U12178 ( .A1(n11671), .A2(i_data_bus[763]), .B1(n11670), 
        .B2(i_data_bus[795]), .ZN(n11580) );
  AOI22D1BWP30P140LVT U12179 ( .A1(n11672), .A2(i_data_bus[667]), .B1(n11686), 
        .B2(i_data_bus[475]), .ZN(n11579) );
  AOI22D1BWP30P140LVT U12180 ( .A1(n11676), .A2(i_data_bus[859]), .B1(n11687), 
        .B2(i_data_bus[347]), .ZN(n11578) );
  AOI22D1BWP30P140LVT U12181 ( .A1(n11684), .A2(i_data_bus[187]), .B1(n11683), 
        .B2(i_data_bus[699]), .ZN(n11577) );
  ND4D1BWP30P140LVT U12182 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(n11581) );
  OR4D1BWP30P140LVT U12183 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .Z(o_data_bus[59]) );
  AOI22D1BWP30P140LVT U12184 ( .A1(n11658), .A2(i_data_bus[540]), .B1(n11647), 
        .B2(i_data_bus[988]), .ZN(n11588) );
  AOI22D1BWP30P140LVT U12185 ( .A1(n11659), .A2(i_data_bus[956]), .B1(n11649), 
        .B2(i_data_bus[924]), .ZN(n11587) );
  AOI22D1BWP30P140LVT U12186 ( .A1(n11651), .A2(i_data_bus[604]), .B1(n11657), 
        .B2(i_data_bus[636]), .ZN(n11586) );
  AOI22D1BWP30P140LVT U12187 ( .A1(n11660), .A2(i_data_bus[124]), .B1(n11645), 
        .B2(i_data_bus[92]), .ZN(n11585) );
  ND4D1BWP30P140LVT U12188 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(n11604) );
  AOI22D1BWP30P140LVT U12189 ( .A1(n11650), .A2(i_data_bus[572]), .B1(n11652), 
        .B2(i_data_bus[28]), .ZN(n11592) );
  AOI22D1BWP30P140LVT U12190 ( .A1(n11646), .A2(i_data_bus[1020]), .B1(n11648), 
        .B2(i_data_bus[60]), .ZN(n11591) );
  AOI22D1BWP30P140LVT U12191 ( .A1(n11685), .A2(i_data_bus[380]), .B1(n11687), 
        .B2(i_data_bus[348]), .ZN(n11590) );
  AOI22D1BWP30P140LVT U12192 ( .A1(n11662), .A2(i_data_bus[444]), .B1(n11670), 
        .B2(i_data_bus[796]), .ZN(n11589) );
  ND4D1BWP30P140LVT U12193 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(n11603) );
  AOI22D1BWP30P140LVT U12194 ( .A1(n11669), .A2(i_data_bus[732]), .B1(n11688), 
        .B2(i_data_bus[252]), .ZN(n11596) );
  AOI22D1BWP30P140LVT U12195 ( .A1(n11664), .A2(i_data_bus[508]), .B1(n11681), 
        .B2(i_data_bus[892]), .ZN(n11595) );
  AOI22D1BWP30P140LVT U12196 ( .A1(n11682), .A2(i_data_bus[156]), .B1(n11673), 
        .B2(i_data_bus[828]), .ZN(n11594) );
  AOI22D1BWP30P140LVT U12197 ( .A1(n11674), .A2(i_data_bus[412]), .B1(n11675), 
        .B2(i_data_bus[220]), .ZN(n11593) );
  ND4D1BWP30P140LVT U12198 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(n11602) );
  AOI22D1BWP30P140LVT U12199 ( .A1(n11672), .A2(i_data_bus[668]), .B1(n11671), 
        .B2(i_data_bus[764]), .ZN(n11600) );
  AOI22D1BWP30P140LVT U12200 ( .A1(n11676), .A2(i_data_bus[860]), .B1(n11684), 
        .B2(i_data_bus[188]), .ZN(n11599) );
  AOI22D1BWP30P140LVT U12201 ( .A1(n11686), .A2(i_data_bus[476]), .B1(n11683), 
        .B2(i_data_bus[700]), .ZN(n11598) );
  AOI22D1BWP30P140LVT U12202 ( .A1(n11661), .A2(i_data_bus[316]), .B1(n11663), 
        .B2(i_data_bus[284]), .ZN(n11597) );
  ND4D1BWP30P140LVT U12203 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(n11601) );
  OR4D1BWP30P140LVT U12204 ( .A1(n11604), .A2(n11603), .A3(n11602), .A4(n11601), .Z(o_data_bus[60]) );
  AOI22D1BWP30P140LVT U12205 ( .A1(n11659), .A2(i_data_bus[957]), .B1(n11649), 
        .B2(i_data_bus[925]), .ZN(n11608) );
  AOI22D1BWP30P140LVT U12206 ( .A1(n11650), .A2(i_data_bus[573]), .B1(n11652), 
        .B2(i_data_bus[29]), .ZN(n11607) );
  AOI22D1BWP30P140LVT U12207 ( .A1(n11647), .A2(i_data_bus[989]), .B1(n11657), 
        .B2(i_data_bus[637]), .ZN(n11606) );
  AOI22D1BWP30P140LVT U12208 ( .A1(n11646), .A2(i_data_bus[1021]), .B1(n11660), 
        .B2(i_data_bus[125]), .ZN(n11605) );
  ND4D1BWP30P140LVT U12209 ( .A1(n11608), .A2(n11607), .A3(n11606), .A4(n11605), .ZN(n11624) );
  AOI22D1BWP30P140LVT U12210 ( .A1(n11658), .A2(i_data_bus[541]), .B1(n11651), 
        .B2(i_data_bus[605]), .ZN(n11612) );
  AOI22D1BWP30P140LVT U12211 ( .A1(n11648), .A2(i_data_bus[61]), .B1(n11645), 
        .B2(i_data_bus[93]), .ZN(n11611) );
  AOI22D1BWP30P140LVT U12212 ( .A1(n11682), .A2(i_data_bus[157]), .B1(n11683), 
        .B2(i_data_bus[701]), .ZN(n11610) );
  AOI22D1BWP30P140LVT U12213 ( .A1(n11662), .A2(i_data_bus[445]), .B1(n11672), 
        .B2(i_data_bus[669]), .ZN(n11609) );
  ND4D1BWP30P140LVT U12214 ( .A1(n11612), .A2(n11611), .A3(n11610), .A4(n11609), .ZN(n11623) );
  AOI22D1BWP30P140LVT U12215 ( .A1(n11671), .A2(i_data_bus[765]), .B1(n11661), 
        .B2(i_data_bus[317]), .ZN(n11616) );
  AOI22D1BWP30P140LVT U12216 ( .A1(n11664), .A2(i_data_bus[509]), .B1(n11684), 
        .B2(i_data_bus[189]), .ZN(n11615) );
  AOI22D1BWP30P140LVT U12217 ( .A1(n11670), .A2(i_data_bus[797]), .B1(n11687), 
        .B2(i_data_bus[349]), .ZN(n11614) );
  AOI22D1BWP30P140LVT U12218 ( .A1(n11686), .A2(i_data_bus[477]), .B1(n11669), 
        .B2(i_data_bus[733]), .ZN(n11613) );
  ND4D1BWP30P140LVT U12219 ( .A1(n11616), .A2(n11615), .A3(n11614), .A4(n11613), .ZN(n11622) );
  AOI22D1BWP30P140LVT U12220 ( .A1(n11674), .A2(i_data_bus[413]), .B1(n11685), 
        .B2(i_data_bus[381]), .ZN(n11620) );
  AOI22D1BWP30P140LVT U12221 ( .A1(n11688), .A2(i_data_bus[253]), .B1(n11663), 
        .B2(i_data_bus[285]), .ZN(n11619) );
  AOI22D1BWP30P140LVT U12222 ( .A1(n11676), .A2(i_data_bus[861]), .B1(n11673), 
        .B2(i_data_bus[829]), .ZN(n11618) );
  AOI22D1BWP30P140LVT U12223 ( .A1(n11675), .A2(i_data_bus[221]), .B1(n11681), 
        .B2(i_data_bus[893]), .ZN(n11617) );
  ND4D1BWP30P140LVT U12224 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(n11621) );
  OR4D1BWP30P140LVT U12225 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .Z(o_data_bus[61]) );
  AOI22D1BWP30P140LVT U12226 ( .A1(n11648), .A2(i_data_bus[62]), .B1(n11649), 
        .B2(i_data_bus[926]), .ZN(n11628) );
  AOI22D1BWP30P140LVT U12227 ( .A1(n11658), .A2(i_data_bus[542]), .B1(n11659), 
        .B2(i_data_bus[958]), .ZN(n11627) );
  AOI22D1BWP30P140LVT U12228 ( .A1(n11650), .A2(i_data_bus[574]), .B1(n11660), 
        .B2(i_data_bus[126]), .ZN(n11626) );
  AOI22D1BWP30P140LVT U12229 ( .A1(n11646), .A2(i_data_bus[1022]), .B1(n11647), 
        .B2(i_data_bus[990]), .ZN(n11625) );
  ND4D1BWP30P140LVT U12230 ( .A1(n11628), .A2(n11627), .A3(n11626), .A4(n11625), .ZN(n11644) );
  AOI22D1BWP30P140LVT U12231 ( .A1(n11652), .A2(i_data_bus[30]), .B1(n11645), 
        .B2(i_data_bus[94]), .ZN(n11632) );
  AOI22D1BWP30P140LVT U12232 ( .A1(n11651), .A2(i_data_bus[606]), .B1(n11657), 
        .B2(i_data_bus[638]), .ZN(n11631) );
  AOI22D1BWP30P140LVT U12233 ( .A1(n11672), .A2(i_data_bus[670]), .B1(n11675), 
        .B2(i_data_bus[222]), .ZN(n11630) );
  AOI22D1BWP30P140LVT U12234 ( .A1(n11662), .A2(i_data_bus[446]), .B1(n11687), 
        .B2(i_data_bus[350]), .ZN(n11629) );
  ND4D1BWP30P140LVT U12235 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(n11643) );
  AOI22D1BWP30P140LVT U12236 ( .A1(n11676), .A2(i_data_bus[862]), .B1(n11661), 
        .B2(i_data_bus[318]), .ZN(n11636) );
  AOI22D1BWP30P140LVT U12237 ( .A1(n11670), .A2(i_data_bus[798]), .B1(n11663), 
        .B2(i_data_bus[286]), .ZN(n11635) );
  AOI22D1BWP30P140LVT U12238 ( .A1(n11671), .A2(i_data_bus[766]), .B1(n11684), 
        .B2(i_data_bus[190]), .ZN(n11634) );
  AOI22D1BWP30P140LVT U12239 ( .A1(n11688), .A2(i_data_bus[254]), .B1(n11673), 
        .B2(i_data_bus[830]), .ZN(n11633) );
  ND4D1BWP30P140LVT U12240 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(n11642) );
  AOI22D1BWP30P140LVT U12241 ( .A1(n11674), .A2(i_data_bus[414]), .B1(n11686), 
        .B2(i_data_bus[478]), .ZN(n11640) );
  AOI22D1BWP30P140LVT U12242 ( .A1(n11664), .A2(i_data_bus[510]), .B1(n11683), 
        .B2(i_data_bus[702]), .ZN(n11639) );
  AOI22D1BWP30P140LVT U12243 ( .A1(n11685), .A2(i_data_bus[382]), .B1(n11669), 
        .B2(i_data_bus[734]), .ZN(n11638) );
  AOI22D1BWP30P140LVT U12244 ( .A1(n11682), .A2(i_data_bus[158]), .B1(n11681), 
        .B2(i_data_bus[894]), .ZN(n11637) );
  ND4D1BWP30P140LVT U12245 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(n11641) );
  OR4D1BWP30P140LVT U12246 ( .A1(n11644), .A2(n11643), .A3(n11642), .A4(n11641), .Z(o_data_bus[62]) );
  AOI22D1BWP30P140LVT U12247 ( .A1(n11646), .A2(i_data_bus[1023]), .B1(n11645), 
        .B2(i_data_bus[95]), .ZN(n11656) );
  AOI22D1BWP30P140LVT U12248 ( .A1(n11648), .A2(i_data_bus[63]), .B1(n11647), 
        .B2(i_data_bus[991]), .ZN(n11655) );
  AOI22D1BWP30P140LVT U12249 ( .A1(n11650), .A2(i_data_bus[575]), .B1(n11649), 
        .B2(i_data_bus[927]), .ZN(n11654) );
  AOI22D1BWP30P140LVT U12250 ( .A1(n11652), .A2(i_data_bus[31]), .B1(n11651), 
        .B2(i_data_bus[607]), .ZN(n11653) );
  ND4D1BWP30P140LVT U12251 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(n11696) );
  AOI22D1BWP30P140LVT U12252 ( .A1(n11658), .A2(i_data_bus[543]), .B1(n11657), 
        .B2(i_data_bus[639]), .ZN(n11668) );
  AOI22D1BWP30P140LVT U12253 ( .A1(n11660), .A2(i_data_bus[127]), .B1(n11659), 
        .B2(i_data_bus[959]), .ZN(n11667) );
  AOI22D1BWP30P140LVT U12254 ( .A1(n11662), .A2(i_data_bus[447]), .B1(n11661), 
        .B2(i_data_bus[319]), .ZN(n11666) );
  AOI22D1BWP30P140LVT U12255 ( .A1(n11664), .A2(i_data_bus[511]), .B1(n11663), 
        .B2(i_data_bus[287]), .ZN(n11665) );
  ND4D1BWP30P140LVT U12256 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(n11695) );
  AOI22D1BWP30P140LVT U12257 ( .A1(n11670), .A2(i_data_bus[799]), .B1(n11669), 
        .B2(i_data_bus[735]), .ZN(n11680) );
  AOI22D1BWP30P140LVT U12258 ( .A1(n11672), .A2(i_data_bus[671]), .B1(n11671), 
        .B2(i_data_bus[767]), .ZN(n11679) );
  AOI22D1BWP30P140LVT U12259 ( .A1(n11674), .A2(i_data_bus[415]), .B1(n11673), 
        .B2(i_data_bus[831]), .ZN(n11678) );
  AOI22D1BWP30P140LVT U12260 ( .A1(n11676), .A2(i_data_bus[863]), .B1(n11675), 
        .B2(i_data_bus[223]), .ZN(n11677) );
  ND4D1BWP30P140LVT U12261 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(n11694) );
  AOI22D1BWP30P140LVT U12262 ( .A1(n11682), .A2(i_data_bus[159]), .B1(n11681), 
        .B2(i_data_bus[895]), .ZN(n11692) );
  AOI22D1BWP30P140LVT U12263 ( .A1(n11684), .A2(i_data_bus[191]), .B1(n11683), 
        .B2(i_data_bus[703]), .ZN(n11691) );
  AOI22D1BWP30P140LVT U12264 ( .A1(n11686), .A2(i_data_bus[479]), .B1(n11685), 
        .B2(i_data_bus[383]), .ZN(n11690) );
  AOI22D1BWP30P140LVT U12265 ( .A1(n11688), .A2(i_data_bus[255]), .B1(n11687), 
        .B2(i_data_bus[351]), .ZN(n11689) );
  ND4D1BWP30P140LVT U12266 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(n11693) );
  OR4D1BWP30P140LVT U12267 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .Z(o_data_bus[63]) );
  INR3D0BWP30P140LVT U12268 ( .A1(i_cmd[155]), .B1(n11697), .B2(n11732), .ZN(
        n12366) );
  INR3D0BWP30P140LVT U12269 ( .A1(i_cmd[107]), .B1(n11698), .B2(n11718), .ZN(
        n12377) );
  AOI22D1BWP30P140LVT U12270 ( .A1(i_data_bus[608]), .A2(n12366), .B1(
        i_data_bus[416]), .B2(n12377), .ZN(n11710) );
  INR3D0BWP30P140LVT U12271 ( .A1(i_cmd[19]), .B1(n11699), .B2(n11736), .ZN(
        n12382) );
  INR3D0BWP30P140LVT U12272 ( .A1(i_cmd[83]), .B1(n11700), .B2(n11730), .ZN(
        n12369) );
  AOI22D1BWP30P140LVT U12273 ( .A1(i_data_bus[64]), .A2(n12382), .B1(
        i_data_bus[320]), .B2(n12369), .ZN(n11709) );
  INR3D0BWP30P140LVT U12274 ( .A1(i_cmd[139]), .B1(n11701), .B2(n11732), .ZN(
        n12381) );
  NR3D0P7BWP30P140LVT U12275 ( .A1(n11703), .A2(n11702), .A3(n11736), .ZN(
        n12393) );
  AOI22D1BWP30P140LVT U12276 ( .A1(i_data_bus[544]), .A2(n12381), .B1(
        i_data_bus[0]), .B2(n12393), .ZN(n11708) );
  INVD1BWP30P140LVT U12277 ( .I(i_cmd[99]), .ZN(n11704) );
  NR3D0P7BWP30P140LVT U12278 ( .A1(n11705), .A2(n11704), .A3(n11718), .ZN(
        n12365) );
  INR3D0BWP30P140LVT U12279 ( .A1(i_cmd[115]), .B1(n11706), .B2(n11718), .ZN(
        n12391) );
  AOI22D1BWP30P140LVT U12280 ( .A1(i_data_bus[384]), .A2(n12365), .B1(
        i_data_bus[448]), .B2(n12391), .ZN(n11707) );
  ND4D1BWP30P140LVT U12281 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(n11764) );
  AN3D1BWP30P140LVT U12282 ( .A1(i_valid[7]), .A2(i_cmd[59]), .A3(n11729), .Z(
        n12367) );
  INR3D0BWP30P140LVT U12283 ( .A1(i_cmd[75]), .B1(n11711), .B2(n11730), .ZN(
        n12378) );
  AOI22D1BWP30P140LVT U12284 ( .A1(i_data_bus[224]), .A2(n12367), .B1(
        i_data_bus[288]), .B2(n12378), .ZN(n11725) );
  NR3D0P7BWP30P140LVT U12285 ( .A1(n11713), .A2(n11712), .A3(n11732), .ZN(
        n12384) );
  NR3D0P7BWP30P140LVT U12286 ( .A1(n11715), .A2(n11714), .A3(n11738), .ZN(
        n12380) );
  AOI22D1BWP30P140LVT U12287 ( .A1(i_data_bus[512]), .A2(n12384), .B1(
        i_data_bus[960]), .B2(n12380), .ZN(n11724) );
  NR3D0P7BWP30P140LVT U12288 ( .A1(n11717), .A2(n11716), .A3(n11738), .ZN(
        n12394) );
  INR3D0BWP30P140LVT U12289 ( .A1(i_cmd[123]), .B1(n11719), .B2(n11718), .ZN(
        n12390) );
  AOI22D1BWP30P140LVT U12290 ( .A1(i_data_bus[992]), .A2(n12394), .B1(
        i_data_bus[480]), .B2(n12390), .ZN(n11723) );
  INR3D0BWP30P140LVT U12291 ( .A1(n11729), .B1(n11721), .B2(n11720), .ZN(
        n12395) );
  AN3D1BWP30P140LVT U12292 ( .A1(i_valid[6]), .A2(i_cmd[51]), .A3(n11729), .Z(
        n12372) );
  AOI22D1BWP30P140LVT U12293 ( .A1(i_data_bus[128]), .A2(n12395), .B1(
        i_data_bus[192]), .B2(n12372), .ZN(n11722) );
  ND4D1BWP30P140LVT U12294 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(n11763) );
  INR3D0BWP30P140LVT U12295 ( .A1(i_cmd[27]), .B1(n11726), .B2(n11736), .ZN(
        n12396) );
  INVD1BWP30P140LVT U12296 ( .I(i_cmd[67]), .ZN(n11727) );
  NR3D0P7BWP30P140LVT U12297 ( .A1(n11728), .A2(n11727), .A3(n11730), .ZN(
        n12389) );
  AOI22D1BWP30P140LVT U12298 ( .A1(i_data_bus[96]), .A2(n12396), .B1(
        i_data_bus[256]), .B2(n12389), .ZN(n11744) );
  AN3D1BWP30P140LVT U12299 ( .A1(i_valid[5]), .A2(i_cmd[43]), .A3(n11729), .Z(
        n12371) );
  INR3D0BWP30P140LVT U12300 ( .A1(i_cmd[91]), .B1(n11731), .B2(n11730), .ZN(
        n12383) );
  AOI22D1BWP30P140LVT U12301 ( .A1(i_data_bus[160]), .A2(n12371), .B1(
        i_data_bus[352]), .B2(n12383), .ZN(n11743) );
  INR3D0BWP30P140LVT U12302 ( .A1(i_cmd[147]), .B1(n11733), .B2(n11732), .ZN(
        n12368) );
  NR3D0P7BWP30P140LVT U12303 ( .A1(n11735), .A2(n11734), .A3(n11738), .ZN(
        n12392) );
  AOI22D1BWP30P140LVT U12304 ( .A1(i_data_bus[576]), .A2(n12368), .B1(
        i_data_bus[896]), .B2(n12392), .ZN(n11742) );
  INR3D0BWP30P140LVT U12305 ( .A1(i_cmd[11]), .B1(n11737), .B2(n11736), .ZN(
        n12370) );
  NR3D0P7BWP30P140LVT U12306 ( .A1(n11740), .A2(n11739), .A3(n11738), .ZN(
        n12379) );
  AOI22D1BWP30P140LVT U12307 ( .A1(i_data_bus[32]), .A2(n12370), .B1(
        i_data_bus[928]), .B2(n12379), .ZN(n11741) );
  ND4D1BWP30P140LVT U12308 ( .A1(n11744), .A2(n11743), .A3(n11742), .A4(n11741), .ZN(n11762) );
  INR3D0BWP30P140LVT U12309 ( .A1(i_cmd[211]), .B1(n11745), .B2(n11752), .ZN(
        n12408) );
  NR3D0P7BWP30P140LVT U12310 ( .A1(n11747), .A2(n11746), .A3(n11755), .ZN(
        n12404) );
  AOI22D1BWP30P140LVT U12311 ( .A1(i_data_bus[832]), .A2(n12408), .B1(
        i_data_bus[640]), .B2(n12404), .ZN(n11760) );
  INR3D0BWP30P140LVT U12312 ( .A1(i_cmd[179]), .B1(n11748), .B2(n11755), .ZN(
        n12402) );
  INR3D0BWP30P140LVT U12313 ( .A1(i_cmd[219]), .B1(n11749), .B2(n11752), .ZN(
        n12401) );
  AOI22D1BWP30P140LVT U12314 ( .A1(i_data_bus[704]), .A2(n12402), .B1(
        i_data_bus[864]), .B2(n12401), .ZN(n11759) );
  INR3D0BWP30P140LVT U12315 ( .A1(i_cmd[187]), .B1(n11750), .B2(n11755), .ZN(
        n12405) );
  INR3D0BWP30P140LVT U12316 ( .A1(i_cmd[203]), .B1(n11751), .B2(n11752), .ZN(
        n12403) );
  AOI22D1BWP30P140LVT U12317 ( .A1(i_data_bus[736]), .A2(n12405), .B1(
        i_data_bus[800]), .B2(n12403), .ZN(n11758) );
  INVD1BWP30P140LVT U12318 ( .I(i_cmd[195]), .ZN(n11753) );
  NR3D0P7BWP30P140LVT U12319 ( .A1(n11754), .A2(n11753), .A3(n11752), .ZN(
        n12406) );
  INR3D0BWP30P140LVT U12320 ( .A1(i_cmd[171]), .B1(n11756), .B2(n11755), .ZN(
        n12407) );
  AOI22D1BWP30P140LVT U12321 ( .A1(i_data_bus[768]), .A2(n12406), .B1(
        i_data_bus[672]), .B2(n12407), .ZN(n11757) );
  ND4D1BWP30P140LVT U12322 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(n11761) );
  OR4D1BWP30P140LVT U12323 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .Z(o_data_bus[96]) );
  AOI22D1BWP30P140LVT U12324 ( .A1(i_data_bus[385]), .A2(n12365), .B1(
        i_data_bus[225]), .B2(n12367), .ZN(n11768) );
  AOI22D1BWP30P140LVT U12325 ( .A1(i_data_bus[65]), .A2(n12382), .B1(
        i_data_bus[513]), .B2(n12384), .ZN(n11767) );
  AOI22D1BWP30P140LVT U12326 ( .A1(i_data_bus[929]), .A2(n12379), .B1(
        i_data_bus[129]), .B2(n12395), .ZN(n11766) );
  AOI22D1BWP30P140LVT U12327 ( .A1(i_data_bus[33]), .A2(n12370), .B1(
        i_data_bus[161]), .B2(n12371), .ZN(n11765) );
  ND4D1BWP30P140LVT U12328 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(n11784) );
  AOI22D1BWP30P140LVT U12329 ( .A1(i_data_bus[97]), .A2(n12396), .B1(
        i_data_bus[1]), .B2(n12393), .ZN(n11772) );
  AOI22D1BWP30P140LVT U12330 ( .A1(i_data_bus[257]), .A2(n12389), .B1(
        i_data_bus[449]), .B2(n12391), .ZN(n11771) );
  AOI22D1BWP30P140LVT U12331 ( .A1(i_data_bus[897]), .A2(n12392), .B1(
        i_data_bus[481]), .B2(n12390), .ZN(n11770) );
  AOI22D1BWP30P140LVT U12332 ( .A1(i_data_bus[289]), .A2(n12378), .B1(
        i_data_bus[321]), .B2(n12369), .ZN(n11769) );
  ND4D1BWP30P140LVT U12333 ( .A1(n11772), .A2(n11771), .A3(n11770), .A4(n11769), .ZN(n11783) );
  AOI22D1BWP30P140LVT U12334 ( .A1(i_data_bus[993]), .A2(n12394), .B1(
        i_data_bus[609]), .B2(n12366), .ZN(n11776) );
  AOI22D1BWP30P140LVT U12335 ( .A1(i_data_bus[961]), .A2(n12380), .B1(
        i_data_bus[193]), .B2(n12372), .ZN(n11775) );
  AOI22D1BWP30P140LVT U12336 ( .A1(i_data_bus[577]), .A2(n12368), .B1(
        i_data_bus[417]), .B2(n12377), .ZN(n11774) );
  AOI22D1BWP30P140LVT U12337 ( .A1(i_data_bus[545]), .A2(n12381), .B1(
        i_data_bus[353]), .B2(n12383), .ZN(n11773) );
  ND4D1BWP30P140LVT U12338 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(n11782) );
  AOI22D1BWP30P140LVT U12339 ( .A1(i_data_bus[769]), .A2(n12406), .B1(
        i_data_bus[737]), .B2(n12405), .ZN(n11780) );
  AOI22D1BWP30P140LVT U12340 ( .A1(i_data_bus[705]), .A2(n12402), .B1(
        i_data_bus[641]), .B2(n12404), .ZN(n11779) );
  AOI22D1BWP30P140LVT U12341 ( .A1(i_data_bus[673]), .A2(n12407), .B1(
        i_data_bus[865]), .B2(n12401), .ZN(n11778) );
  AOI22D1BWP30P140LVT U12342 ( .A1(i_data_bus[801]), .A2(n12403), .B1(
        i_data_bus[833]), .B2(n12408), .ZN(n11777) );
  ND4D1BWP30P140LVT U12343 ( .A1(n11780), .A2(n11779), .A3(n11778), .A4(n11777), .ZN(n11781) );
  OR4D1BWP30P140LVT U12344 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .Z(o_data_bus[97]) );
  AOI22D1BWP30P140LVT U12345 ( .A1(i_data_bus[546]), .A2(n12381), .B1(
        i_data_bus[226]), .B2(n12367), .ZN(n11788) );
  AOI22D1BWP30P140LVT U12346 ( .A1(i_data_bus[578]), .A2(n12368), .B1(
        i_data_bus[130]), .B2(n12395), .ZN(n11787) );
  AOI22D1BWP30P140LVT U12347 ( .A1(i_data_bus[2]), .A2(n12393), .B1(
        i_data_bus[194]), .B2(n12372), .ZN(n11786) );
  AOI22D1BWP30P140LVT U12348 ( .A1(i_data_bus[162]), .A2(n12371), .B1(
        i_data_bus[450]), .B2(n12391), .ZN(n11785) );
  ND4D1BWP30P140LVT U12349 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(n11804) );
  AOI22D1BWP30P140LVT U12350 ( .A1(i_data_bus[482]), .A2(n12390), .B1(
        i_data_bus[258]), .B2(n12389), .ZN(n11792) );
  AOI22D1BWP30P140LVT U12351 ( .A1(i_data_bus[994]), .A2(n12394), .B1(
        i_data_bus[354]), .B2(n12383), .ZN(n11791) );
  AOI22D1BWP30P140LVT U12352 ( .A1(i_data_bus[98]), .A2(n12396), .B1(
        i_data_bus[418]), .B2(n12377), .ZN(n11790) );
  AOI22D1BWP30P140LVT U12353 ( .A1(i_data_bus[930]), .A2(n12379), .B1(
        i_data_bus[290]), .B2(n12378), .ZN(n11789) );
  ND4D1BWP30P140LVT U12354 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(n11803) );
  AOI22D1BWP30P140LVT U12355 ( .A1(i_data_bus[898]), .A2(n12392), .B1(
        i_data_bus[514]), .B2(n12384), .ZN(n11796) );
  AOI22D1BWP30P140LVT U12356 ( .A1(i_data_bus[386]), .A2(n12365), .B1(
        i_data_bus[322]), .B2(n12369), .ZN(n11795) );
  AOI22D1BWP30P140LVT U12357 ( .A1(i_data_bus[66]), .A2(n12382), .B1(
        i_data_bus[610]), .B2(n12366), .ZN(n11794) );
  AOI22D1BWP30P140LVT U12358 ( .A1(i_data_bus[962]), .A2(n12380), .B1(
        i_data_bus[34]), .B2(n12370), .ZN(n11793) );
  ND4D1BWP30P140LVT U12359 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(n11802) );
  AOI22D1BWP30P140LVT U12360 ( .A1(i_data_bus[834]), .A2(n12408), .B1(
        i_data_bus[642]), .B2(n12404), .ZN(n11800) );
  AOI22D1BWP30P140LVT U12361 ( .A1(i_data_bus[866]), .A2(n12401), .B1(
        i_data_bus[738]), .B2(n12405), .ZN(n11799) );
  AOI22D1BWP30P140LVT U12362 ( .A1(i_data_bus[674]), .A2(n12407), .B1(
        i_data_bus[706]), .B2(n12402), .ZN(n11798) );
  AOI22D1BWP30P140LVT U12363 ( .A1(i_data_bus[802]), .A2(n12403), .B1(
        i_data_bus[770]), .B2(n12406), .ZN(n11797) );
  ND4D1BWP30P140LVT U12364 ( .A1(n11800), .A2(n11799), .A3(n11798), .A4(n11797), .ZN(n11801) );
  OR4D1BWP30P140LVT U12365 ( .A1(n11804), .A2(n11803), .A3(n11802), .A4(n11801), .Z(o_data_bus[98]) );
  AOI22D1BWP30P140LVT U12366 ( .A1(i_data_bus[67]), .A2(n12382), .B1(
        i_data_bus[899]), .B2(n12392), .ZN(n11808) );
  AOI22D1BWP30P140LVT U12367 ( .A1(i_data_bus[35]), .A2(n12370), .B1(
        i_data_bus[451]), .B2(n12391), .ZN(n11807) );
  AOI22D1BWP30P140LVT U12368 ( .A1(i_data_bus[963]), .A2(n12380), .B1(
        i_data_bus[163]), .B2(n12371), .ZN(n11806) );
  AOI22D1BWP30P140LVT U12369 ( .A1(i_data_bus[259]), .A2(n12389), .B1(
        i_data_bus[227]), .B2(n12367), .ZN(n11805) );
  ND4D1BWP30P140LVT U12370 ( .A1(n11808), .A2(n11807), .A3(n11806), .A4(n11805), .ZN(n11824) );
  AOI22D1BWP30P140LVT U12371 ( .A1(i_data_bus[579]), .A2(n12368), .B1(
        i_data_bus[3]), .B2(n12393), .ZN(n11812) );
  AOI22D1BWP30P140LVT U12372 ( .A1(i_data_bus[515]), .A2(n12384), .B1(
        i_data_bus[547]), .B2(n12381), .ZN(n11811) );
  AOI22D1BWP30P140LVT U12373 ( .A1(i_data_bus[995]), .A2(n12394), .B1(
        i_data_bus[483]), .B2(n12390), .ZN(n11810) );
  AOI22D1BWP30P140LVT U12374 ( .A1(i_data_bus[419]), .A2(n12377), .B1(
        i_data_bus[323]), .B2(n12369), .ZN(n11809) );
  ND4D1BWP30P140LVT U12375 ( .A1(n11812), .A2(n11811), .A3(n11810), .A4(n11809), .ZN(n11823) );
  AOI22D1BWP30P140LVT U12376 ( .A1(i_data_bus[931]), .A2(n12379), .B1(
        i_data_bus[355]), .B2(n12383), .ZN(n11816) );
  AOI22D1BWP30P140LVT U12377 ( .A1(i_data_bus[611]), .A2(n12366), .B1(
        i_data_bus[291]), .B2(n12378), .ZN(n11815) );
  AOI22D1BWP30P140LVT U12378 ( .A1(i_data_bus[387]), .A2(n12365), .B1(
        i_data_bus[195]), .B2(n12372), .ZN(n11814) );
  AOI22D1BWP30P140LVT U12379 ( .A1(i_data_bus[99]), .A2(n12396), .B1(
        i_data_bus[131]), .B2(n12395), .ZN(n11813) );
  ND4D1BWP30P140LVT U12380 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(n11822) );
  AOI22D1BWP30P140LVT U12381 ( .A1(i_data_bus[835]), .A2(n12408), .B1(
        i_data_bus[739]), .B2(n12405), .ZN(n11820) );
  AOI22D1BWP30P140LVT U12382 ( .A1(i_data_bus[771]), .A2(n12406), .B1(
        i_data_bus[803]), .B2(n12403), .ZN(n11819) );
  AOI22D1BWP30P140LVT U12383 ( .A1(i_data_bus[643]), .A2(n12404), .B1(
        i_data_bus[707]), .B2(n12402), .ZN(n11818) );
  AOI22D1BWP30P140LVT U12384 ( .A1(i_data_bus[675]), .A2(n12407), .B1(
        i_data_bus[867]), .B2(n12401), .ZN(n11817) );
  ND4D1BWP30P140LVT U12385 ( .A1(n11820), .A2(n11819), .A3(n11818), .A4(n11817), .ZN(n11821) );
  OR4D1BWP30P140LVT U12386 ( .A1(n11824), .A2(n11823), .A3(n11822), .A4(n11821), .Z(o_data_bus[99]) );
  AOI22D1BWP30P140LVT U12387 ( .A1(i_data_bus[548]), .A2(n12381), .B1(
        i_data_bus[36]), .B2(n12370), .ZN(n11828) );
  AOI22D1BWP30P140LVT U12388 ( .A1(i_data_bus[900]), .A2(n12392), .B1(
        i_data_bus[356]), .B2(n12383), .ZN(n11827) );
  AOI22D1BWP30P140LVT U12389 ( .A1(i_data_bus[964]), .A2(n12380), .B1(
        i_data_bus[68]), .B2(n12382), .ZN(n11826) );
  AOI22D1BWP30P140LVT U12390 ( .A1(i_data_bus[996]), .A2(n12394), .B1(
        i_data_bus[484]), .B2(n12390), .ZN(n11825) );
  ND4D1BWP30P140LVT U12391 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(n11844) );
  AOI22D1BWP30P140LVT U12392 ( .A1(i_data_bus[516]), .A2(n12384), .B1(
        i_data_bus[420]), .B2(n12377), .ZN(n11832) );
  AOI22D1BWP30P140LVT U12393 ( .A1(i_data_bus[324]), .A2(n12369), .B1(
        i_data_bus[260]), .B2(n12389), .ZN(n11831) );
  AOI22D1BWP30P140LVT U12394 ( .A1(i_data_bus[932]), .A2(n12379), .B1(
        i_data_bus[164]), .B2(n12371), .ZN(n11830) );
  AOI22D1BWP30P140LVT U12395 ( .A1(i_data_bus[100]), .A2(n12396), .B1(
        i_data_bus[196]), .B2(n12372), .ZN(n11829) );
  ND4D1BWP30P140LVT U12396 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(n11843) );
  AOI22D1BWP30P140LVT U12397 ( .A1(i_data_bus[228]), .A2(n12367), .B1(
        i_data_bus[452]), .B2(n12391), .ZN(n11836) );
  AOI22D1BWP30P140LVT U12398 ( .A1(i_data_bus[612]), .A2(n12366), .B1(
        i_data_bus[292]), .B2(n12378), .ZN(n11835) );
  AOI22D1BWP30P140LVT U12399 ( .A1(i_data_bus[4]), .A2(n12393), .B1(
        i_data_bus[580]), .B2(n12368), .ZN(n11834) );
  AOI22D1BWP30P140LVT U12400 ( .A1(i_data_bus[132]), .A2(n12395), .B1(
        i_data_bus[388]), .B2(n12365), .ZN(n11833) );
  ND4D1BWP30P140LVT U12401 ( .A1(n11836), .A2(n11835), .A3(n11834), .A4(n11833), .ZN(n11842) );
  AOI22D1BWP30P140LVT U12402 ( .A1(i_data_bus[740]), .A2(n12405), .B1(
        i_data_bus[772]), .B2(n12406), .ZN(n11840) );
  AOI22D1BWP30P140LVT U12403 ( .A1(i_data_bus[836]), .A2(n12408), .B1(
        i_data_bus[804]), .B2(n12403), .ZN(n11839) );
  AOI22D1BWP30P140LVT U12404 ( .A1(i_data_bus[708]), .A2(n12402), .B1(
        i_data_bus[644]), .B2(n12404), .ZN(n11838) );
  AOI22D1BWP30P140LVT U12405 ( .A1(i_data_bus[868]), .A2(n12401), .B1(
        i_data_bus[676]), .B2(n12407), .ZN(n11837) );
  ND4D1BWP30P140LVT U12406 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(n11841) );
  OR4D1BWP30P140LVT U12407 ( .A1(n11844), .A2(n11843), .A3(n11842), .A4(n11841), .Z(o_data_bus[100]) );
  AOI22D1BWP30P140LVT U12408 ( .A1(i_data_bus[133]), .A2(n12395), .B1(
        i_data_bus[229]), .B2(n12367), .ZN(n11848) );
  AOI22D1BWP30P140LVT U12409 ( .A1(i_data_bus[933]), .A2(n12379), .B1(
        i_data_bus[613]), .B2(n12366), .ZN(n11847) );
  AOI22D1BWP30P140LVT U12410 ( .A1(i_data_bus[997]), .A2(n12394), .B1(
        i_data_bus[261]), .B2(n12389), .ZN(n11846) );
  AOI22D1BWP30P140LVT U12411 ( .A1(i_data_bus[101]), .A2(n12396), .B1(
        i_data_bus[965]), .B2(n12380), .ZN(n11845) );
  ND4D1BWP30P140LVT U12412 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(n11864) );
  AOI22D1BWP30P140LVT U12413 ( .A1(i_data_bus[581]), .A2(n12368), .B1(
        i_data_bus[421]), .B2(n12377), .ZN(n11852) );
  AOI22D1BWP30P140LVT U12414 ( .A1(i_data_bus[197]), .A2(n12372), .B1(
        i_data_bus[453]), .B2(n12391), .ZN(n11851) );
  AOI22D1BWP30P140LVT U12415 ( .A1(i_data_bus[517]), .A2(n12384), .B1(
        i_data_bus[549]), .B2(n12381), .ZN(n11850) );
  AOI22D1BWP30P140LVT U12416 ( .A1(i_data_bus[485]), .A2(n12390), .B1(
        i_data_bus[293]), .B2(n12378), .ZN(n11849) );
  ND4D1BWP30P140LVT U12417 ( .A1(n11852), .A2(n11851), .A3(n11850), .A4(n11849), .ZN(n11863) );
  AOI22D1BWP30P140LVT U12418 ( .A1(i_data_bus[69]), .A2(n12382), .B1(
        i_data_bus[357]), .B2(n12383), .ZN(n11856) );
  AOI22D1BWP30P140LVT U12419 ( .A1(i_data_bus[5]), .A2(n12393), .B1(
        i_data_bus[325]), .B2(n12369), .ZN(n11855) );
  AOI22D1BWP30P140LVT U12420 ( .A1(i_data_bus[37]), .A2(n12370), .B1(
        i_data_bus[389]), .B2(n12365), .ZN(n11854) );
  AOI22D1BWP30P140LVT U12421 ( .A1(i_data_bus[901]), .A2(n12392), .B1(
        i_data_bus[165]), .B2(n12371), .ZN(n11853) );
  ND4D1BWP30P140LVT U12422 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(n11862) );
  AOI22D1BWP30P140LVT U12423 ( .A1(i_data_bus[773]), .A2(n12406), .B1(
        i_data_bus[837]), .B2(n12408), .ZN(n11860) );
  AOI22D1BWP30P140LVT U12424 ( .A1(i_data_bus[869]), .A2(n12401), .B1(
        i_data_bus[741]), .B2(n12405), .ZN(n11859) );
  AOI22D1BWP30P140LVT U12425 ( .A1(i_data_bus[677]), .A2(n12407), .B1(
        i_data_bus[805]), .B2(n12403), .ZN(n11858) );
  AOI22D1BWP30P140LVT U12426 ( .A1(i_data_bus[645]), .A2(n12404), .B1(
        i_data_bus[709]), .B2(n12402), .ZN(n11857) );
  ND4D1BWP30P140LVT U12427 ( .A1(n11860), .A2(n11859), .A3(n11858), .A4(n11857), .ZN(n11861) );
  OR4D1BWP30P140LVT U12428 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11861), .Z(o_data_bus[101]) );
  AOI22D1BWP30P140LVT U12429 ( .A1(i_data_bus[966]), .A2(n12380), .B1(
        i_data_bus[518]), .B2(n12384), .ZN(n11868) );
  AOI22D1BWP30P140LVT U12430 ( .A1(i_data_bus[6]), .A2(n12393), .B1(
        i_data_bus[102]), .B2(n12396), .ZN(n11867) );
  AOI22D1BWP30P140LVT U12431 ( .A1(i_data_bus[902]), .A2(n12392), .B1(
        i_data_bus[326]), .B2(n12369), .ZN(n11866) );
  AOI22D1BWP30P140LVT U12432 ( .A1(i_data_bus[582]), .A2(n12368), .B1(
        i_data_bus[38]), .B2(n12370), .ZN(n11865) );
  ND4D1BWP30P140LVT U12433 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(n11884) );
  AOI22D1BWP30P140LVT U12434 ( .A1(i_data_bus[358]), .A2(n12383), .B1(
        i_data_bus[294]), .B2(n12378), .ZN(n11872) );
  AOI22D1BWP30P140LVT U12435 ( .A1(i_data_bus[166]), .A2(n12371), .B1(
        i_data_bus[422]), .B2(n12377), .ZN(n11871) );
  AOI22D1BWP30P140LVT U12436 ( .A1(i_data_bus[486]), .A2(n12390), .B1(
        i_data_bus[390]), .B2(n12365), .ZN(n11870) );
  AOI22D1BWP30P140LVT U12437 ( .A1(i_data_bus[550]), .A2(n12381), .B1(
        i_data_bus[230]), .B2(n12367), .ZN(n11869) );
  ND4D1BWP30P140LVT U12438 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(n11883) );
  AOI22D1BWP30P140LVT U12439 ( .A1(i_data_bus[998]), .A2(n12394), .B1(
        i_data_bus[262]), .B2(n12389), .ZN(n11876) );
  AOI22D1BWP30P140LVT U12440 ( .A1(i_data_bus[614]), .A2(n12366), .B1(
        i_data_bus[934]), .B2(n12379), .ZN(n11875) );
  AOI22D1BWP30P140LVT U12441 ( .A1(i_data_bus[198]), .A2(n12372), .B1(
        i_data_bus[134]), .B2(n12395), .ZN(n11874) );
  AOI22D1BWP30P140LVT U12442 ( .A1(i_data_bus[70]), .A2(n12382), .B1(
        i_data_bus[454]), .B2(n12391), .ZN(n11873) );
  ND4D1BWP30P140LVT U12443 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(n11882) );
  AOI22D1BWP30P140LVT U12444 ( .A1(i_data_bus[838]), .A2(n12408), .B1(
        i_data_bus[646]), .B2(n12404), .ZN(n11880) );
  AOI22D1BWP30P140LVT U12445 ( .A1(i_data_bus[870]), .A2(n12401), .B1(
        i_data_bus[678]), .B2(n12407), .ZN(n11879) );
  AOI22D1BWP30P140LVT U12446 ( .A1(i_data_bus[742]), .A2(n12405), .B1(
        i_data_bus[774]), .B2(n12406), .ZN(n11878) );
  AOI22D1BWP30P140LVT U12447 ( .A1(i_data_bus[806]), .A2(n12403), .B1(
        i_data_bus[710]), .B2(n12402), .ZN(n11877) );
  ND4D1BWP30P140LVT U12448 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(n11881) );
  OR4D1BWP30P140LVT U12449 ( .A1(n11884), .A2(n11883), .A3(n11882), .A4(n11881), .Z(o_data_bus[102]) );
  AOI22D1BWP30P140LVT U12450 ( .A1(i_data_bus[551]), .A2(n12381), .B1(
        i_data_bus[135]), .B2(n12395), .ZN(n11888) );
  AOI22D1BWP30P140LVT U12451 ( .A1(i_data_bus[39]), .A2(n12370), .B1(
        i_data_bus[999]), .B2(n12394), .ZN(n11887) );
  AOI22D1BWP30P140LVT U12452 ( .A1(i_data_bus[295]), .A2(n12378), .B1(
        i_data_bus[199]), .B2(n12372), .ZN(n11886) );
  AOI22D1BWP30P140LVT U12453 ( .A1(i_data_bus[903]), .A2(n12392), .B1(
        i_data_bus[167]), .B2(n12371), .ZN(n11885) );
  ND4D1BWP30P140LVT U12454 ( .A1(n11888), .A2(n11887), .A3(n11886), .A4(n11885), .ZN(n11904) );
  AOI22D1BWP30P140LVT U12455 ( .A1(i_data_bus[519]), .A2(n12384), .B1(
        i_data_bus[487]), .B2(n12390), .ZN(n11892) );
  AOI22D1BWP30P140LVT U12456 ( .A1(i_data_bus[103]), .A2(n12396), .B1(
        i_data_bus[935]), .B2(n12379), .ZN(n11891) );
  AOI22D1BWP30P140LVT U12457 ( .A1(i_data_bus[583]), .A2(n12368), .B1(
        i_data_bus[263]), .B2(n12389), .ZN(n11890) );
  AOI22D1BWP30P140LVT U12458 ( .A1(i_data_bus[455]), .A2(n12391), .B1(
        i_data_bus[231]), .B2(n12367), .ZN(n11889) );
  ND4D1BWP30P140LVT U12459 ( .A1(n11892), .A2(n11891), .A3(n11890), .A4(n11889), .ZN(n11903) );
  AOI22D1BWP30P140LVT U12460 ( .A1(i_data_bus[391]), .A2(n12365), .B1(
        i_data_bus[423]), .B2(n12377), .ZN(n11896) );
  AOI22D1BWP30P140LVT U12461 ( .A1(i_data_bus[615]), .A2(n12366), .B1(
        i_data_bus[7]), .B2(n12393), .ZN(n11895) );
  AOI22D1BWP30P140LVT U12462 ( .A1(i_data_bus[967]), .A2(n12380), .B1(
        i_data_bus[71]), .B2(n12382), .ZN(n11894) );
  AOI22D1BWP30P140LVT U12463 ( .A1(i_data_bus[359]), .A2(n12383), .B1(
        i_data_bus[327]), .B2(n12369), .ZN(n11893) );
  ND4D1BWP30P140LVT U12464 ( .A1(n11896), .A2(n11895), .A3(n11894), .A4(n11893), .ZN(n11902) );
  AOI22D1BWP30P140LVT U12465 ( .A1(i_data_bus[743]), .A2(n12405), .B1(
        i_data_bus[775]), .B2(n12406), .ZN(n11900) );
  AOI22D1BWP30P140LVT U12466 ( .A1(i_data_bus[807]), .A2(n12403), .B1(
        i_data_bus[647]), .B2(n12404), .ZN(n11899) );
  AOI22D1BWP30P140LVT U12467 ( .A1(i_data_bus[679]), .A2(n12407), .B1(
        i_data_bus[711]), .B2(n12402), .ZN(n11898) );
  AOI22D1BWP30P140LVT U12468 ( .A1(i_data_bus[871]), .A2(n12401), .B1(
        i_data_bus[839]), .B2(n12408), .ZN(n11897) );
  ND4D1BWP30P140LVT U12469 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(n11901) );
  OR4D1BWP30P140LVT U12470 ( .A1(n11904), .A2(n11903), .A3(n11902), .A4(n11901), .Z(o_data_bus[103]) );
  AOI22D1BWP30P140LVT U12471 ( .A1(i_data_bus[584]), .A2(n12368), .B1(
        i_data_bus[200]), .B2(n12372), .ZN(n11908) );
  AOI22D1BWP30P140LVT U12472 ( .A1(i_data_bus[104]), .A2(n12396), .B1(
        i_data_bus[168]), .B2(n12371), .ZN(n11907) );
  AOI22D1BWP30P140LVT U12473 ( .A1(i_data_bus[520]), .A2(n12384), .B1(
        i_data_bus[456]), .B2(n12391), .ZN(n11906) );
  AOI22D1BWP30P140LVT U12474 ( .A1(i_data_bus[968]), .A2(n12380), .B1(
        i_data_bus[424]), .B2(n12377), .ZN(n11905) );
  ND4D1BWP30P140LVT U12475 ( .A1(n11908), .A2(n11907), .A3(n11906), .A4(n11905), .ZN(n11924) );
  AOI22D1BWP30P140LVT U12476 ( .A1(i_data_bus[360]), .A2(n12383), .B1(
        i_data_bus[232]), .B2(n12367), .ZN(n11912) );
  AOI22D1BWP30P140LVT U12477 ( .A1(i_data_bus[1000]), .A2(n12394), .B1(
        i_data_bus[136]), .B2(n12395), .ZN(n11911) );
  AOI22D1BWP30P140LVT U12478 ( .A1(i_data_bus[8]), .A2(n12393), .B1(
        i_data_bus[488]), .B2(n12390), .ZN(n11910) );
  AOI22D1BWP30P140LVT U12479 ( .A1(i_data_bus[936]), .A2(n12379), .B1(
        i_data_bus[392]), .B2(n12365), .ZN(n11909) );
  ND4D1BWP30P140LVT U12480 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(n11923) );
  AOI22D1BWP30P140LVT U12481 ( .A1(i_data_bus[616]), .A2(n12366), .B1(
        i_data_bus[328]), .B2(n12369), .ZN(n11916) );
  AOI22D1BWP30P140LVT U12482 ( .A1(i_data_bus[264]), .A2(n12389), .B1(
        i_data_bus[296]), .B2(n12378), .ZN(n11915) );
  AOI22D1BWP30P140LVT U12483 ( .A1(i_data_bus[904]), .A2(n12392), .B1(
        i_data_bus[72]), .B2(n12382), .ZN(n11914) );
  AOI22D1BWP30P140LVT U12484 ( .A1(i_data_bus[552]), .A2(n12381), .B1(
        i_data_bus[40]), .B2(n12370), .ZN(n11913) );
  ND4D1BWP30P140LVT U12485 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(n11922) );
  AOI22D1BWP30P140LVT U12486 ( .A1(i_data_bus[680]), .A2(n12407), .B1(
        i_data_bus[808]), .B2(n12403), .ZN(n11920) );
  AOI22D1BWP30P140LVT U12487 ( .A1(i_data_bus[712]), .A2(n12402), .B1(
        i_data_bus[776]), .B2(n12406), .ZN(n11919) );
  AOI22D1BWP30P140LVT U12488 ( .A1(i_data_bus[744]), .A2(n12405), .B1(
        i_data_bus[648]), .B2(n12404), .ZN(n11918) );
  AOI22D1BWP30P140LVT U12489 ( .A1(i_data_bus[840]), .A2(n12408), .B1(
        i_data_bus[872]), .B2(n12401), .ZN(n11917) );
  ND4D1BWP30P140LVT U12490 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(n11921) );
  OR4D1BWP30P140LVT U12491 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .Z(o_data_bus[104]) );
  AOI22D1BWP30P140LVT U12492 ( .A1(i_data_bus[521]), .A2(n12384), .B1(
        i_data_bus[73]), .B2(n12382), .ZN(n11928) );
  AOI22D1BWP30P140LVT U12493 ( .A1(i_data_bus[1001]), .A2(n12394), .B1(
        i_data_bus[169]), .B2(n12371), .ZN(n11927) );
  AOI22D1BWP30P140LVT U12494 ( .A1(i_data_bus[905]), .A2(n12392), .B1(
        i_data_bus[41]), .B2(n12370), .ZN(n11926) );
  AOI22D1BWP30P140LVT U12495 ( .A1(i_data_bus[489]), .A2(n12390), .B1(
        i_data_bus[137]), .B2(n12395), .ZN(n11925) );
  ND4D1BWP30P140LVT U12496 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(n11944) );
  AOI22D1BWP30P140LVT U12497 ( .A1(i_data_bus[617]), .A2(n12366), .B1(
        i_data_bus[297]), .B2(n12378), .ZN(n11932) );
  AOI22D1BWP30P140LVT U12498 ( .A1(i_data_bus[105]), .A2(n12396), .B1(
        i_data_bus[457]), .B2(n12391), .ZN(n11931) );
  AOI22D1BWP30P140LVT U12499 ( .A1(i_data_bus[969]), .A2(n12380), .B1(
        i_data_bus[329]), .B2(n12369), .ZN(n11930) );
  AOI22D1BWP30P140LVT U12500 ( .A1(i_data_bus[585]), .A2(n12368), .B1(
        i_data_bus[361]), .B2(n12383), .ZN(n11929) );
  ND4D1BWP30P140LVT U12501 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(n11943) );
  AOI22D1BWP30P140LVT U12502 ( .A1(i_data_bus[937]), .A2(n12379), .B1(
        i_data_bus[425]), .B2(n12377), .ZN(n11936) );
  AOI22D1BWP30P140LVT U12503 ( .A1(i_data_bus[201]), .A2(n12372), .B1(
        i_data_bus[265]), .B2(n12389), .ZN(n11935) );
  AOI22D1BWP30P140LVT U12504 ( .A1(i_data_bus[9]), .A2(n12393), .B1(
        i_data_bus[553]), .B2(n12381), .ZN(n11934) );
  AOI22D1BWP30P140LVT U12505 ( .A1(i_data_bus[233]), .A2(n12367), .B1(
        i_data_bus[393]), .B2(n12365), .ZN(n11933) );
  ND4D1BWP30P140LVT U12506 ( .A1(n11936), .A2(n11935), .A3(n11934), .A4(n11933), .ZN(n11942) );
  AOI22D1BWP30P140LVT U12507 ( .A1(i_data_bus[873]), .A2(n12401), .B1(
        i_data_bus[841]), .B2(n12408), .ZN(n11940) );
  AOI22D1BWP30P140LVT U12508 ( .A1(i_data_bus[809]), .A2(n12403), .B1(
        i_data_bus[777]), .B2(n12406), .ZN(n11939) );
  AOI22D1BWP30P140LVT U12509 ( .A1(i_data_bus[681]), .A2(n12407), .B1(
        i_data_bus[713]), .B2(n12402), .ZN(n11938) );
  AOI22D1BWP30P140LVT U12510 ( .A1(i_data_bus[745]), .A2(n12405), .B1(
        i_data_bus[649]), .B2(n12404), .ZN(n11937) );
  ND4D1BWP30P140LVT U12511 ( .A1(n11940), .A2(n11939), .A3(n11938), .A4(n11937), .ZN(n11941) );
  OR4D1BWP30P140LVT U12512 ( .A1(n11944), .A2(n11943), .A3(n11942), .A4(n11941), .Z(o_data_bus[105]) );
  AOI22D1BWP30P140LVT U12513 ( .A1(i_data_bus[906]), .A2(n12392), .B1(
        i_data_bus[394]), .B2(n12365), .ZN(n11948) );
  AOI22D1BWP30P140LVT U12514 ( .A1(i_data_bus[106]), .A2(n12396), .B1(
        i_data_bus[938]), .B2(n12379), .ZN(n11947) );
  AOI22D1BWP30P140LVT U12515 ( .A1(i_data_bus[202]), .A2(n12372), .B1(
        i_data_bus[298]), .B2(n12378), .ZN(n11946) );
  AOI22D1BWP30P140LVT U12516 ( .A1(i_data_bus[490]), .A2(n12390), .B1(
        i_data_bus[266]), .B2(n12389), .ZN(n11945) );
  ND4D1BWP30P140LVT U12517 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(n11964) );
  AOI22D1BWP30P140LVT U12518 ( .A1(i_data_bus[554]), .A2(n12381), .B1(
        i_data_bus[458]), .B2(n12391), .ZN(n11952) );
  AOI22D1BWP30P140LVT U12519 ( .A1(i_data_bus[234]), .A2(n12367), .B1(
        i_data_bus[426]), .B2(n12377), .ZN(n11951) );
  AOI22D1BWP30P140LVT U12520 ( .A1(i_data_bus[1002]), .A2(n12394), .B1(
        i_data_bus[138]), .B2(n12395), .ZN(n11950) );
  AOI22D1BWP30P140LVT U12521 ( .A1(i_data_bus[970]), .A2(n12380), .B1(
        i_data_bus[362]), .B2(n12383), .ZN(n11949) );
  ND4D1BWP30P140LVT U12522 ( .A1(n11952), .A2(n11951), .A3(n11950), .A4(n11949), .ZN(n11963) );
  AOI22D1BWP30P140LVT U12523 ( .A1(i_data_bus[74]), .A2(n12382), .B1(
        i_data_bus[522]), .B2(n12384), .ZN(n11956) );
  AOI22D1BWP30P140LVT U12524 ( .A1(i_data_bus[586]), .A2(n12368), .B1(
        i_data_bus[330]), .B2(n12369), .ZN(n11955) );
  AOI22D1BWP30P140LVT U12525 ( .A1(i_data_bus[10]), .A2(n12393), .B1(
        i_data_bus[618]), .B2(n12366), .ZN(n11954) );
  AOI22D1BWP30P140LVT U12526 ( .A1(i_data_bus[42]), .A2(n12370), .B1(
        i_data_bus[170]), .B2(n12371), .ZN(n11953) );
  ND4D1BWP30P140LVT U12527 ( .A1(n11956), .A2(n11955), .A3(n11954), .A4(n11953), .ZN(n11962) );
  AOI22D1BWP30P140LVT U12528 ( .A1(i_data_bus[874]), .A2(n12401), .B1(
        i_data_bus[714]), .B2(n12402), .ZN(n11960) );
  AOI22D1BWP30P140LVT U12529 ( .A1(i_data_bus[842]), .A2(n12408), .B1(
        i_data_bus[682]), .B2(n12407), .ZN(n11959) );
  AOI22D1BWP30P140LVT U12530 ( .A1(i_data_bus[778]), .A2(n12406), .B1(
        i_data_bus[810]), .B2(n12403), .ZN(n11958) );
  AOI22D1BWP30P140LVT U12531 ( .A1(i_data_bus[650]), .A2(n12404), .B1(
        i_data_bus[746]), .B2(n12405), .ZN(n11957) );
  ND4D1BWP30P140LVT U12532 ( .A1(n11960), .A2(n11959), .A3(n11958), .A4(n11957), .ZN(n11961) );
  OR4D1BWP30P140LVT U12533 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .Z(o_data_bus[106]) );
  AOI22D1BWP30P140LVT U12534 ( .A1(i_data_bus[523]), .A2(n12384), .B1(
        i_data_bus[203]), .B2(n12372), .ZN(n11968) );
  AOI22D1BWP30P140LVT U12535 ( .A1(i_data_bus[555]), .A2(n12381), .B1(
        i_data_bus[139]), .B2(n12395), .ZN(n11967) );
  AOI22D1BWP30P140LVT U12536 ( .A1(i_data_bus[43]), .A2(n12370), .B1(
        i_data_bus[171]), .B2(n12371), .ZN(n11966) );
  AOI22D1BWP30P140LVT U12537 ( .A1(i_data_bus[427]), .A2(n12377), .B1(
        i_data_bus[299]), .B2(n12378), .ZN(n11965) );
  ND4D1BWP30P140LVT U12538 ( .A1(n11968), .A2(n11967), .A3(n11966), .A4(n11965), .ZN(n11984) );
  AOI22D1BWP30P140LVT U12539 ( .A1(i_data_bus[235]), .A2(n12367), .B1(
        i_data_bus[267]), .B2(n12389), .ZN(n11972) );
  AOI22D1BWP30P140LVT U12540 ( .A1(i_data_bus[907]), .A2(n12392), .B1(
        i_data_bus[363]), .B2(n12383), .ZN(n11971) );
  AOI22D1BWP30P140LVT U12541 ( .A1(i_data_bus[1003]), .A2(n12394), .B1(
        i_data_bus[491]), .B2(n12390), .ZN(n11970) );
  AOI22D1BWP30P140LVT U12542 ( .A1(i_data_bus[587]), .A2(n12368), .B1(
        i_data_bus[395]), .B2(n12365), .ZN(n11969) );
  ND4D1BWP30P140LVT U12543 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(n11983) );
  AOI22D1BWP30P140LVT U12544 ( .A1(i_data_bus[11]), .A2(n12393), .B1(
        i_data_bus[459]), .B2(n12391), .ZN(n11976) );
  AOI22D1BWP30P140LVT U12545 ( .A1(i_data_bus[619]), .A2(n12366), .B1(
        i_data_bus[331]), .B2(n12369), .ZN(n11975) );
  AOI22D1BWP30P140LVT U12546 ( .A1(i_data_bus[939]), .A2(n12379), .B1(
        i_data_bus[107]), .B2(n12396), .ZN(n11974) );
  AOI22D1BWP30P140LVT U12547 ( .A1(i_data_bus[971]), .A2(n12380), .B1(
        i_data_bus[75]), .B2(n12382), .ZN(n11973) );
  ND4D1BWP30P140LVT U12548 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(n11982) );
  AOI22D1BWP30P140LVT U12549 ( .A1(i_data_bus[843]), .A2(n12408), .B1(
        i_data_bus[779]), .B2(n12406), .ZN(n11980) );
  AOI22D1BWP30P140LVT U12550 ( .A1(i_data_bus[875]), .A2(n12401), .B1(
        i_data_bus[715]), .B2(n12402), .ZN(n11979) );
  AOI22D1BWP30P140LVT U12551 ( .A1(i_data_bus[811]), .A2(n12403), .B1(
        i_data_bus[683]), .B2(n12407), .ZN(n11978) );
  AOI22D1BWP30P140LVT U12552 ( .A1(i_data_bus[747]), .A2(n12405), .B1(
        i_data_bus[651]), .B2(n12404), .ZN(n11977) );
  ND4D1BWP30P140LVT U12553 ( .A1(n11980), .A2(n11979), .A3(n11978), .A4(n11977), .ZN(n11981) );
  OR4D1BWP30P140LVT U12554 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .Z(o_data_bus[107]) );
  AOI22D1BWP30P140LVT U12555 ( .A1(i_data_bus[556]), .A2(n12381), .B1(
        i_data_bus[588]), .B2(n12368), .ZN(n11988) );
  AOI22D1BWP30P140LVT U12556 ( .A1(i_data_bus[1004]), .A2(n12394), .B1(
        i_data_bus[364]), .B2(n12383), .ZN(n11987) );
  AOI22D1BWP30P140LVT U12557 ( .A1(i_data_bus[428]), .A2(n12377), .B1(
        i_data_bus[204]), .B2(n12372), .ZN(n11986) );
  AOI22D1BWP30P140LVT U12558 ( .A1(i_data_bus[12]), .A2(n12393), .B1(
        i_data_bus[908]), .B2(n12392), .ZN(n11985) );
  ND4D1BWP30P140LVT U12559 ( .A1(n11988), .A2(n11987), .A3(n11986), .A4(n11985), .ZN(n12004) );
  AOI22D1BWP30P140LVT U12560 ( .A1(i_data_bus[972]), .A2(n12380), .B1(
        i_data_bus[108]), .B2(n12396), .ZN(n11992) );
  AOI22D1BWP30P140LVT U12561 ( .A1(i_data_bus[140]), .A2(n12395), .B1(
        i_data_bus[396]), .B2(n12365), .ZN(n11991) );
  AOI22D1BWP30P140LVT U12562 ( .A1(i_data_bus[236]), .A2(n12367), .B1(
        i_data_bus[172]), .B2(n12371), .ZN(n11990) );
  AOI22D1BWP30P140LVT U12563 ( .A1(i_data_bus[460]), .A2(n12391), .B1(
        i_data_bus[268]), .B2(n12389), .ZN(n11989) );
  ND4D1BWP30P140LVT U12564 ( .A1(n11992), .A2(n11991), .A3(n11990), .A4(n11989), .ZN(n12003) );
  AOI22D1BWP30P140LVT U12565 ( .A1(i_data_bus[300]), .A2(n12378), .B1(
        i_data_bus[332]), .B2(n12369), .ZN(n11996) );
  AOI22D1BWP30P140LVT U12566 ( .A1(i_data_bus[76]), .A2(n12382), .B1(
        i_data_bus[492]), .B2(n12390), .ZN(n11995) );
  AOI22D1BWP30P140LVT U12567 ( .A1(i_data_bus[620]), .A2(n12366), .B1(
        i_data_bus[44]), .B2(n12370), .ZN(n11994) );
  AOI22D1BWP30P140LVT U12568 ( .A1(i_data_bus[940]), .A2(n12379), .B1(
        i_data_bus[524]), .B2(n12384), .ZN(n11993) );
  ND4D1BWP30P140LVT U12569 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(n12002) );
  AOI22D1BWP30P140LVT U12570 ( .A1(i_data_bus[780]), .A2(n12406), .B1(
        i_data_bus[652]), .B2(n12404), .ZN(n12000) );
  AOI22D1BWP30P140LVT U12571 ( .A1(i_data_bus[812]), .A2(n12403), .B1(
        i_data_bus[876]), .B2(n12401), .ZN(n11999) );
  AOI22D1BWP30P140LVT U12572 ( .A1(i_data_bus[684]), .A2(n12407), .B1(
        i_data_bus[844]), .B2(n12408), .ZN(n11998) );
  AOI22D1BWP30P140LVT U12573 ( .A1(i_data_bus[716]), .A2(n12402), .B1(
        i_data_bus[748]), .B2(n12405), .ZN(n11997) );
  ND4D1BWP30P140LVT U12574 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(n12001) );
  OR4D1BWP30P140LVT U12575 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .Z(o_data_bus[108]) );
  AOI22D1BWP30P140LVT U12576 ( .A1(i_data_bus[973]), .A2(n12380), .B1(
        i_data_bus[493]), .B2(n12390), .ZN(n12008) );
  AOI22D1BWP30P140LVT U12577 ( .A1(i_data_bus[397]), .A2(n12365), .B1(
        i_data_bus[365]), .B2(n12383), .ZN(n12007) );
  AOI22D1BWP30P140LVT U12578 ( .A1(i_data_bus[621]), .A2(n12366), .B1(
        i_data_bus[141]), .B2(n12395), .ZN(n12006) );
  AOI22D1BWP30P140LVT U12579 ( .A1(i_data_bus[589]), .A2(n12368), .B1(
        i_data_bus[13]), .B2(n12393), .ZN(n12005) );
  ND4D1BWP30P140LVT U12580 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(n12024) );
  AOI22D1BWP30P140LVT U12581 ( .A1(i_data_bus[45]), .A2(n12370), .B1(
        i_data_bus[525]), .B2(n12384), .ZN(n12012) );
  AOI22D1BWP30P140LVT U12582 ( .A1(i_data_bus[941]), .A2(n12379), .B1(
        i_data_bus[461]), .B2(n12391), .ZN(n12011) );
  AOI22D1BWP30P140LVT U12583 ( .A1(i_data_bus[909]), .A2(n12392), .B1(
        i_data_bus[109]), .B2(n12396), .ZN(n12010) );
  AOI22D1BWP30P140LVT U12584 ( .A1(i_data_bus[77]), .A2(n12382), .B1(
        i_data_bus[205]), .B2(n12372), .ZN(n12009) );
  ND4D1BWP30P140LVT U12585 ( .A1(n12012), .A2(n12011), .A3(n12010), .A4(n12009), .ZN(n12023) );
  AOI22D1BWP30P140LVT U12586 ( .A1(i_data_bus[429]), .A2(n12377), .B1(
        i_data_bus[301]), .B2(n12378), .ZN(n12016) );
  AOI22D1BWP30P140LVT U12587 ( .A1(i_data_bus[237]), .A2(n12367), .B1(
        i_data_bus[269]), .B2(n12389), .ZN(n12015) );
  AOI22D1BWP30P140LVT U12588 ( .A1(i_data_bus[1005]), .A2(n12394), .B1(
        i_data_bus[173]), .B2(n12371), .ZN(n12014) );
  AOI22D1BWP30P140LVT U12589 ( .A1(i_data_bus[557]), .A2(n12381), .B1(
        i_data_bus[333]), .B2(n12369), .ZN(n12013) );
  ND4D1BWP30P140LVT U12590 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(n12022) );
  AOI22D1BWP30P140LVT U12591 ( .A1(i_data_bus[877]), .A2(n12401), .B1(
        i_data_bus[717]), .B2(n12402), .ZN(n12020) );
  AOI22D1BWP30P140LVT U12592 ( .A1(i_data_bus[781]), .A2(n12406), .B1(
        i_data_bus[813]), .B2(n12403), .ZN(n12019) );
  AOI22D1BWP30P140LVT U12593 ( .A1(i_data_bus[749]), .A2(n12405), .B1(
        i_data_bus[685]), .B2(n12407), .ZN(n12018) );
  AOI22D1BWP30P140LVT U12594 ( .A1(i_data_bus[845]), .A2(n12408), .B1(
        i_data_bus[653]), .B2(n12404), .ZN(n12017) );
  ND4D1BWP30P140LVT U12595 ( .A1(n12020), .A2(n12019), .A3(n12018), .A4(n12017), .ZN(n12021) );
  OR4D1BWP30P140LVT U12596 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .Z(o_data_bus[109]) );
  AOI22D1BWP30P140LVT U12597 ( .A1(i_data_bus[14]), .A2(n12393), .B1(
        i_data_bus[398]), .B2(n12365), .ZN(n12028) );
  AOI22D1BWP30P140LVT U12598 ( .A1(i_data_bus[910]), .A2(n12392), .B1(
        i_data_bus[974]), .B2(n12380), .ZN(n12027) );
  AOI22D1BWP30P140LVT U12599 ( .A1(i_data_bus[558]), .A2(n12381), .B1(
        i_data_bus[302]), .B2(n12378), .ZN(n12026) );
  AOI22D1BWP30P140LVT U12600 ( .A1(i_data_bus[174]), .A2(n12371), .B1(
        i_data_bus[334]), .B2(n12369), .ZN(n12025) );
  ND4D1BWP30P140LVT U12601 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(n12044) );
  AOI22D1BWP30P140LVT U12602 ( .A1(i_data_bus[622]), .A2(n12366), .B1(
        i_data_bus[270]), .B2(n12389), .ZN(n12032) );
  AOI22D1BWP30P140LVT U12603 ( .A1(i_data_bus[78]), .A2(n12382), .B1(
        i_data_bus[46]), .B2(n12370), .ZN(n12031) );
  AOI22D1BWP30P140LVT U12604 ( .A1(i_data_bus[590]), .A2(n12368), .B1(
        i_data_bus[238]), .B2(n12367), .ZN(n12030) );
  AOI22D1BWP30P140LVT U12605 ( .A1(i_data_bus[110]), .A2(n12396), .B1(
        i_data_bus[142]), .B2(n12395), .ZN(n12029) );
  ND4D1BWP30P140LVT U12606 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(n12043) );
  AOI22D1BWP30P140LVT U12607 ( .A1(i_data_bus[942]), .A2(n12379), .B1(
        i_data_bus[462]), .B2(n12391), .ZN(n12036) );
  AOI22D1BWP30P140LVT U12608 ( .A1(i_data_bus[1006]), .A2(n12394), .B1(
        i_data_bus[430]), .B2(n12377), .ZN(n12035) );
  AOI22D1BWP30P140LVT U12609 ( .A1(i_data_bus[206]), .A2(n12372), .B1(
        i_data_bus[494]), .B2(n12390), .ZN(n12034) );
  AOI22D1BWP30P140LVT U12610 ( .A1(i_data_bus[526]), .A2(n12384), .B1(
        i_data_bus[366]), .B2(n12383), .ZN(n12033) );
  ND4D1BWP30P140LVT U12611 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(n12042) );
  AOI22D1BWP30P140LVT U12612 ( .A1(i_data_bus[846]), .A2(n12408), .B1(
        i_data_bus[750]), .B2(n12405), .ZN(n12040) );
  AOI22D1BWP30P140LVT U12613 ( .A1(i_data_bus[782]), .A2(n12406), .B1(
        i_data_bus[878]), .B2(n12401), .ZN(n12039) );
  AOI22D1BWP30P140LVT U12614 ( .A1(i_data_bus[686]), .A2(n12407), .B1(
        i_data_bus[654]), .B2(n12404), .ZN(n12038) );
  AOI22D1BWP30P140LVT U12615 ( .A1(i_data_bus[814]), .A2(n12403), .B1(
        i_data_bus[718]), .B2(n12402), .ZN(n12037) );
  ND4D1BWP30P140LVT U12616 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(n12041) );
  OR4D1BWP30P140LVT U12617 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .Z(o_data_bus[110]) );
  AOI22D1BWP30P140LVT U12618 ( .A1(i_data_bus[911]), .A2(n12392), .B1(
        i_data_bus[1007]), .B2(n12394), .ZN(n12048) );
  AOI22D1BWP30P140LVT U12619 ( .A1(i_data_bus[111]), .A2(n12396), .B1(
        i_data_bus[175]), .B2(n12371), .ZN(n12047) );
  AOI22D1BWP30P140LVT U12620 ( .A1(i_data_bus[591]), .A2(n12368), .B1(
        i_data_bus[239]), .B2(n12367), .ZN(n12046) );
  AOI22D1BWP30P140LVT U12621 ( .A1(i_data_bus[975]), .A2(n12380), .B1(
        i_data_bus[79]), .B2(n12382), .ZN(n12045) );
  ND4D1BWP30P140LVT U12622 ( .A1(n12048), .A2(n12047), .A3(n12046), .A4(n12045), .ZN(n12064) );
  AOI22D1BWP30P140LVT U12623 ( .A1(i_data_bus[47]), .A2(n12370), .B1(
        i_data_bus[303]), .B2(n12378), .ZN(n12052) );
  AOI22D1BWP30P140LVT U12624 ( .A1(i_data_bus[527]), .A2(n12384), .B1(
        i_data_bus[335]), .B2(n12369), .ZN(n12051) );
  AOI22D1BWP30P140LVT U12625 ( .A1(i_data_bus[207]), .A2(n12372), .B1(
        i_data_bus[367]), .B2(n12383), .ZN(n12050) );
  AOI22D1BWP30P140LVT U12626 ( .A1(i_data_bus[271]), .A2(n12389), .B1(
        i_data_bus[143]), .B2(n12395), .ZN(n12049) );
  ND4D1BWP30P140LVT U12627 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(n12063) );
  AOI22D1BWP30P140LVT U12628 ( .A1(i_data_bus[559]), .A2(n12381), .B1(
        i_data_bus[15]), .B2(n12393), .ZN(n12056) );
  AOI22D1BWP30P140LVT U12629 ( .A1(i_data_bus[431]), .A2(n12377), .B1(
        i_data_bus[463]), .B2(n12391), .ZN(n12055) );
  AOI22D1BWP30P140LVT U12630 ( .A1(i_data_bus[943]), .A2(n12379), .B1(
        i_data_bus[399]), .B2(n12365), .ZN(n12054) );
  AOI22D1BWP30P140LVT U12631 ( .A1(i_data_bus[623]), .A2(n12366), .B1(
        i_data_bus[495]), .B2(n12390), .ZN(n12053) );
  ND4D1BWP30P140LVT U12632 ( .A1(n12056), .A2(n12055), .A3(n12054), .A4(n12053), .ZN(n12062) );
  AOI22D1BWP30P140LVT U12633 ( .A1(i_data_bus[655]), .A2(n12404), .B1(
        i_data_bus[879]), .B2(n12401), .ZN(n12060) );
  AOI22D1BWP30P140LVT U12634 ( .A1(i_data_bus[719]), .A2(n12402), .B1(
        i_data_bus[687]), .B2(n12407), .ZN(n12059) );
  AOI22D1BWP30P140LVT U12635 ( .A1(i_data_bus[847]), .A2(n12408), .B1(
        i_data_bus[783]), .B2(n12406), .ZN(n12058) );
  AOI22D1BWP30P140LVT U12636 ( .A1(i_data_bus[751]), .A2(n12405), .B1(
        i_data_bus[815]), .B2(n12403), .ZN(n12057) );
  ND4D1BWP30P140LVT U12637 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(n12061) );
  OR4D1BWP30P140LVT U12638 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .Z(o_data_bus[111]) );
  AOI22D1BWP30P140LVT U12639 ( .A1(i_data_bus[80]), .A2(n12382), .B1(
        i_data_bus[368]), .B2(n12383), .ZN(n12068) );
  AOI22D1BWP30P140LVT U12640 ( .A1(i_data_bus[1008]), .A2(n12394), .B1(
        i_data_bus[240]), .B2(n12367), .ZN(n12067) );
  AOI22D1BWP30P140LVT U12641 ( .A1(i_data_bus[912]), .A2(n12392), .B1(
        i_data_bus[112]), .B2(n12396), .ZN(n12066) );
  AOI22D1BWP30P140LVT U12642 ( .A1(i_data_bus[560]), .A2(n12381), .B1(
        i_data_bus[528]), .B2(n12384), .ZN(n12065) );
  ND4D1BWP30P140LVT U12643 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(n12084) );
  AOI22D1BWP30P140LVT U12644 ( .A1(i_data_bus[48]), .A2(n12370), .B1(
        i_data_bus[208]), .B2(n12372), .ZN(n12072) );
  AOI22D1BWP30P140LVT U12645 ( .A1(i_data_bus[336]), .A2(n12369), .B1(
        i_data_bus[144]), .B2(n12395), .ZN(n12071) );
  AOI22D1BWP30P140LVT U12646 ( .A1(i_data_bus[592]), .A2(n12368), .B1(
        i_data_bus[304]), .B2(n12378), .ZN(n12070) );
  AOI22D1BWP30P140LVT U12647 ( .A1(i_data_bus[496]), .A2(n12390), .B1(
        i_data_bus[272]), .B2(n12389), .ZN(n12069) );
  ND4D1BWP30P140LVT U12648 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(n12083) );
  AOI22D1BWP30P140LVT U12649 ( .A1(i_data_bus[16]), .A2(n12393), .B1(
        i_data_bus[464]), .B2(n12391), .ZN(n12076) );
  AOI22D1BWP30P140LVT U12650 ( .A1(i_data_bus[624]), .A2(n12366), .B1(
        i_data_bus[400]), .B2(n12365), .ZN(n12075) );
  AOI22D1BWP30P140LVT U12651 ( .A1(i_data_bus[944]), .A2(n12379), .B1(
        i_data_bus[432]), .B2(n12377), .ZN(n12074) );
  AOI22D1BWP30P140LVT U12652 ( .A1(i_data_bus[976]), .A2(n12380), .B1(
        i_data_bus[176]), .B2(n12371), .ZN(n12073) );
  ND4D1BWP30P140LVT U12653 ( .A1(n12076), .A2(n12075), .A3(n12074), .A4(n12073), .ZN(n12082) );
  AOI22D1BWP30P140LVT U12654 ( .A1(i_data_bus[656]), .A2(n12404), .B1(
        i_data_bus[848]), .B2(n12408), .ZN(n12080) );
  AOI22D1BWP30P140LVT U12655 ( .A1(i_data_bus[880]), .A2(n12401), .B1(
        i_data_bus[688]), .B2(n12407), .ZN(n12079) );
  AOI22D1BWP30P140LVT U12656 ( .A1(i_data_bus[752]), .A2(n12405), .B1(
        i_data_bus[720]), .B2(n12402), .ZN(n12078) );
  AOI22D1BWP30P140LVT U12657 ( .A1(i_data_bus[784]), .A2(n12406), .B1(
        i_data_bus[816]), .B2(n12403), .ZN(n12077) );
  ND4D1BWP30P140LVT U12658 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(n12081) );
  OR4D1BWP30P140LVT U12659 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .Z(o_data_bus[112]) );
  AOI22D1BWP30P140LVT U12660 ( .A1(i_data_bus[1009]), .A2(n12394), .B1(
        i_data_bus[593]), .B2(n12368), .ZN(n12088) );
  AOI22D1BWP30P140LVT U12661 ( .A1(i_data_bus[305]), .A2(n12378), .B1(
        i_data_bus[497]), .B2(n12390), .ZN(n12087) );
  AOI22D1BWP30P140LVT U12662 ( .A1(i_data_bus[113]), .A2(n12396), .B1(
        i_data_bus[273]), .B2(n12389), .ZN(n12086) );
  AOI22D1BWP30P140LVT U12663 ( .A1(i_data_bus[561]), .A2(n12381), .B1(
        i_data_bus[241]), .B2(n12367), .ZN(n12085) );
  ND4D1BWP30P140LVT U12664 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(n12104) );
  AOI22D1BWP30P140LVT U12665 ( .A1(i_data_bus[81]), .A2(n12382), .B1(
        i_data_bus[945]), .B2(n12379), .ZN(n12092) );
  AOI22D1BWP30P140LVT U12666 ( .A1(i_data_bus[401]), .A2(n12365), .B1(
        i_data_bus[209]), .B2(n12372), .ZN(n12091) );
  AOI22D1BWP30P140LVT U12667 ( .A1(i_data_bus[977]), .A2(n12380), .B1(
        i_data_bus[433]), .B2(n12377), .ZN(n12090) );
  AOI22D1BWP30P140LVT U12668 ( .A1(i_data_bus[49]), .A2(n12370), .B1(
        i_data_bus[913]), .B2(n12392), .ZN(n12089) );
  ND4D1BWP30P140LVT U12669 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(n12103) );
  AOI22D1BWP30P140LVT U12670 ( .A1(i_data_bus[145]), .A2(n12395), .B1(
        i_data_bus[177]), .B2(n12371), .ZN(n12096) );
  AOI22D1BWP30P140LVT U12671 ( .A1(i_data_bus[17]), .A2(n12393), .B1(
        i_data_bus[465]), .B2(n12391), .ZN(n12095) );
  AOI22D1BWP30P140LVT U12672 ( .A1(i_data_bus[625]), .A2(n12366), .B1(
        i_data_bus[529]), .B2(n12384), .ZN(n12094) );
  AOI22D1BWP30P140LVT U12673 ( .A1(i_data_bus[337]), .A2(n12369), .B1(
        i_data_bus[369]), .B2(n12383), .ZN(n12093) );
  ND4D1BWP30P140LVT U12674 ( .A1(n12096), .A2(n12095), .A3(n12094), .A4(n12093), .ZN(n12102) );
  AOI22D1BWP30P140LVT U12675 ( .A1(i_data_bus[881]), .A2(n12401), .B1(
        i_data_bus[817]), .B2(n12403), .ZN(n12100) );
  AOI22D1BWP30P140LVT U12676 ( .A1(i_data_bus[785]), .A2(n12406), .B1(
        i_data_bus[657]), .B2(n12404), .ZN(n12099) );
  AOI22D1BWP30P140LVT U12677 ( .A1(i_data_bus[689]), .A2(n12407), .B1(
        i_data_bus[753]), .B2(n12405), .ZN(n12098) );
  AOI22D1BWP30P140LVT U12678 ( .A1(i_data_bus[849]), .A2(n12408), .B1(
        i_data_bus[721]), .B2(n12402), .ZN(n12097) );
  ND4D1BWP30P140LVT U12679 ( .A1(n12100), .A2(n12099), .A3(n12098), .A4(n12097), .ZN(n12101) );
  OR4D1BWP30P140LVT U12680 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .Z(o_data_bus[113]) );
  AOI22D1BWP30P140LVT U12681 ( .A1(i_data_bus[402]), .A2(n12365), .B1(
        i_data_bus[146]), .B2(n12395), .ZN(n12108) );
  AOI22D1BWP30P140LVT U12682 ( .A1(i_data_bus[242]), .A2(n12367), .B1(
        i_data_bus[210]), .B2(n12372), .ZN(n12107) );
  AOI22D1BWP30P140LVT U12683 ( .A1(i_data_bus[530]), .A2(n12384), .B1(
        i_data_bus[82]), .B2(n12382), .ZN(n12106) );
  AOI22D1BWP30P140LVT U12684 ( .A1(i_data_bus[594]), .A2(n12368), .B1(
        i_data_bus[466]), .B2(n12391), .ZN(n12105) );
  ND4D1BWP30P140LVT U12685 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(n12124) );
  AOI22D1BWP30P140LVT U12686 ( .A1(i_data_bus[626]), .A2(n12366), .B1(
        i_data_bus[178]), .B2(n12371), .ZN(n12112) );
  AOI22D1BWP30P140LVT U12687 ( .A1(i_data_bus[914]), .A2(n12392), .B1(
        i_data_bus[370]), .B2(n12383), .ZN(n12111) );
  AOI22D1BWP30P140LVT U12688 ( .A1(i_data_bus[562]), .A2(n12381), .B1(
        i_data_bus[338]), .B2(n12369), .ZN(n12110) );
  AOI22D1BWP30P140LVT U12689 ( .A1(i_data_bus[50]), .A2(n12370), .B1(
        i_data_bus[498]), .B2(n12390), .ZN(n12109) );
  ND4D1BWP30P140LVT U12690 ( .A1(n12112), .A2(n12111), .A3(n12110), .A4(n12109), .ZN(n12123) );
  AOI22D1BWP30P140LVT U12691 ( .A1(i_data_bus[978]), .A2(n12380), .B1(
        i_data_bus[1010]), .B2(n12394), .ZN(n12116) );
  AOI22D1BWP30P140LVT U12692 ( .A1(i_data_bus[274]), .A2(n12389), .B1(
        i_data_bus[434]), .B2(n12377), .ZN(n12115) );
  AOI22D1BWP30P140LVT U12693 ( .A1(i_data_bus[18]), .A2(n12393), .B1(
        i_data_bus[306]), .B2(n12378), .ZN(n12114) );
  AOI22D1BWP30P140LVT U12694 ( .A1(i_data_bus[114]), .A2(n12396), .B1(
        i_data_bus[946]), .B2(n12379), .ZN(n12113) );
  ND4D1BWP30P140LVT U12695 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(n12122) );
  AOI22D1BWP30P140LVT U12696 ( .A1(i_data_bus[882]), .A2(n12401), .B1(
        i_data_bus[850]), .B2(n12408), .ZN(n12120) );
  AOI22D1BWP30P140LVT U12697 ( .A1(i_data_bus[722]), .A2(n12402), .B1(
        i_data_bus[818]), .B2(n12403), .ZN(n12119) );
  AOI22D1BWP30P140LVT U12698 ( .A1(i_data_bus[690]), .A2(n12407), .B1(
        i_data_bus[754]), .B2(n12405), .ZN(n12118) );
  AOI22D1BWP30P140LVT U12699 ( .A1(i_data_bus[658]), .A2(n12404), .B1(
        i_data_bus[786]), .B2(n12406), .ZN(n12117) );
  ND4D1BWP30P140LVT U12700 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(n12121) );
  OR4D1BWP30P140LVT U12701 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .Z(o_data_bus[114]) );
  AOI22D1BWP30P140LVT U12702 ( .A1(i_data_bus[147]), .A2(n12395), .B1(
        i_data_bus[275]), .B2(n12389), .ZN(n12128) );
  AOI22D1BWP30P140LVT U12703 ( .A1(i_data_bus[595]), .A2(n12368), .B1(
        i_data_bus[179]), .B2(n12371), .ZN(n12127) );
  AOI22D1BWP30P140LVT U12704 ( .A1(i_data_bus[339]), .A2(n12369), .B1(
        i_data_bus[435]), .B2(n12377), .ZN(n12126) );
  AOI22D1BWP30P140LVT U12705 ( .A1(i_data_bus[1011]), .A2(n12394), .B1(
        i_data_bus[947]), .B2(n12379), .ZN(n12125) );
  ND4D1BWP30P140LVT U12706 ( .A1(n12128), .A2(n12127), .A3(n12126), .A4(n12125), .ZN(n12144) );
  AOI22D1BWP30P140LVT U12707 ( .A1(i_data_bus[979]), .A2(n12380), .B1(
        i_data_bus[211]), .B2(n12372), .ZN(n12132) );
  AOI22D1BWP30P140LVT U12708 ( .A1(i_data_bus[83]), .A2(n12382), .B1(
        i_data_bus[915]), .B2(n12392), .ZN(n12131) );
  AOI22D1BWP30P140LVT U12709 ( .A1(i_data_bus[627]), .A2(n12366), .B1(
        i_data_bus[371]), .B2(n12383), .ZN(n12130) );
  AOI22D1BWP30P140LVT U12710 ( .A1(i_data_bus[307]), .A2(n12378), .B1(
        i_data_bus[403]), .B2(n12365), .ZN(n12129) );
  ND4D1BWP30P140LVT U12711 ( .A1(n12132), .A2(n12131), .A3(n12130), .A4(n12129), .ZN(n12143) );
  AOI22D1BWP30P140LVT U12712 ( .A1(i_data_bus[563]), .A2(n12381), .B1(
        i_data_bus[531]), .B2(n12384), .ZN(n12136) );
  AOI22D1BWP30P140LVT U12713 ( .A1(i_data_bus[243]), .A2(n12367), .B1(
        i_data_bus[467]), .B2(n12391), .ZN(n12135) );
  AOI22D1BWP30P140LVT U12714 ( .A1(i_data_bus[51]), .A2(n12370), .B1(
        i_data_bus[115]), .B2(n12396), .ZN(n12134) );
  AOI22D1BWP30P140LVT U12715 ( .A1(i_data_bus[19]), .A2(n12393), .B1(
        i_data_bus[499]), .B2(n12390), .ZN(n12133) );
  ND4D1BWP30P140LVT U12716 ( .A1(n12136), .A2(n12135), .A3(n12134), .A4(n12133), .ZN(n12142) );
  AOI22D1BWP30P140LVT U12717 ( .A1(i_data_bus[883]), .A2(n12401), .B1(
        i_data_bus[851]), .B2(n12408), .ZN(n12140) );
  AOI22D1BWP30P140LVT U12718 ( .A1(i_data_bus[819]), .A2(n12403), .B1(
        i_data_bus[787]), .B2(n12406), .ZN(n12139) );
  AOI22D1BWP30P140LVT U12719 ( .A1(i_data_bus[755]), .A2(n12405), .B1(
        i_data_bus[659]), .B2(n12404), .ZN(n12138) );
  AOI22D1BWP30P140LVT U12720 ( .A1(i_data_bus[691]), .A2(n12407), .B1(
        i_data_bus[723]), .B2(n12402), .ZN(n12137) );
  ND4D1BWP30P140LVT U12721 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(n12141) );
  OR4D1BWP30P140LVT U12722 ( .A1(n12144), .A2(n12143), .A3(n12142), .A4(n12141), .Z(o_data_bus[115]) );
  AOI22D1BWP30P140LVT U12723 ( .A1(i_data_bus[916]), .A2(n12392), .B1(
        i_data_bus[276]), .B2(n12389), .ZN(n12148) );
  AOI22D1BWP30P140LVT U12724 ( .A1(i_data_bus[980]), .A2(n12380), .B1(
        i_data_bus[436]), .B2(n12377), .ZN(n12147) );
  AOI22D1BWP30P140LVT U12725 ( .A1(i_data_bus[340]), .A2(n12369), .B1(
        i_data_bus[468]), .B2(n12391), .ZN(n12146) );
  AOI22D1BWP30P140LVT U12726 ( .A1(i_data_bus[116]), .A2(n12396), .B1(
        i_data_bus[404]), .B2(n12365), .ZN(n12145) );
  ND4D1BWP30P140LVT U12727 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(n12164) );
  AOI22D1BWP30P140LVT U12728 ( .A1(i_data_bus[20]), .A2(n12393), .B1(
        i_data_bus[180]), .B2(n12371), .ZN(n12152) );
  AOI22D1BWP30P140LVT U12729 ( .A1(i_data_bus[564]), .A2(n12381), .B1(
        i_data_bus[212]), .B2(n12372), .ZN(n12151) );
  AOI22D1BWP30P140LVT U12730 ( .A1(i_data_bus[628]), .A2(n12366), .B1(
        i_data_bus[948]), .B2(n12379), .ZN(n12150) );
  AOI22D1BWP30P140LVT U12731 ( .A1(i_data_bus[84]), .A2(n12382), .B1(
        i_data_bus[372]), .B2(n12383), .ZN(n12149) );
  ND4D1BWP30P140LVT U12732 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(n12163) );
  AOI22D1BWP30P140LVT U12733 ( .A1(i_data_bus[244]), .A2(n12367), .B1(
        i_data_bus[148]), .B2(n12395), .ZN(n12156) );
  AOI22D1BWP30P140LVT U12734 ( .A1(i_data_bus[532]), .A2(n12384), .B1(
        i_data_bus[308]), .B2(n12378), .ZN(n12155) );
  AOI22D1BWP30P140LVT U12735 ( .A1(i_data_bus[52]), .A2(n12370), .B1(
        i_data_bus[1012]), .B2(n12394), .ZN(n12154) );
  AOI22D1BWP30P140LVT U12736 ( .A1(i_data_bus[596]), .A2(n12368), .B1(
        i_data_bus[500]), .B2(n12390), .ZN(n12153) );
  ND4D1BWP30P140LVT U12737 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(n12162) );
  AOI22D1BWP30P140LVT U12738 ( .A1(i_data_bus[756]), .A2(n12405), .B1(
        i_data_bus[884]), .B2(n12401), .ZN(n12160) );
  AOI22D1BWP30P140LVT U12739 ( .A1(i_data_bus[660]), .A2(n12404), .B1(
        i_data_bus[692]), .B2(n12407), .ZN(n12159) );
  AOI22D1BWP30P140LVT U12740 ( .A1(i_data_bus[724]), .A2(n12402), .B1(
        i_data_bus[820]), .B2(n12403), .ZN(n12158) );
  AOI22D1BWP30P140LVT U12741 ( .A1(i_data_bus[788]), .A2(n12406), .B1(
        i_data_bus[852]), .B2(n12408), .ZN(n12157) );
  ND4D1BWP30P140LVT U12742 ( .A1(n12160), .A2(n12159), .A3(n12158), .A4(n12157), .ZN(n12161) );
  OR4D1BWP30P140LVT U12743 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .Z(o_data_bus[116]) );
  AOI22D1BWP30P140LVT U12744 ( .A1(i_data_bus[533]), .A2(n12384), .B1(
        i_data_bus[373]), .B2(n12383), .ZN(n12168) );
  AOI22D1BWP30P140LVT U12745 ( .A1(i_data_bus[1013]), .A2(n12394), .B1(
        i_data_bus[469]), .B2(n12391), .ZN(n12167) );
  AOI22D1BWP30P140LVT U12746 ( .A1(i_data_bus[181]), .A2(n12371), .B1(
        i_data_bus[501]), .B2(n12390), .ZN(n12166) );
  AOI22D1BWP30P140LVT U12747 ( .A1(i_data_bus[277]), .A2(n12389), .B1(
        i_data_bus[405]), .B2(n12365), .ZN(n12165) );
  ND4D1BWP30P140LVT U12748 ( .A1(n12168), .A2(n12167), .A3(n12166), .A4(n12165), .ZN(n12184) );
  AOI22D1BWP30P140LVT U12749 ( .A1(i_data_bus[213]), .A2(n12372), .B1(
        i_data_bus[245]), .B2(n12367), .ZN(n12172) );
  AOI22D1BWP30P140LVT U12750 ( .A1(i_data_bus[917]), .A2(n12392), .B1(
        i_data_bus[21]), .B2(n12393), .ZN(n12171) );
  AOI22D1BWP30P140LVT U12751 ( .A1(i_data_bus[629]), .A2(n12366), .B1(
        i_data_bus[85]), .B2(n12382), .ZN(n12170) );
  AOI22D1BWP30P140LVT U12752 ( .A1(i_data_bus[117]), .A2(n12396), .B1(
        i_data_bus[149]), .B2(n12395), .ZN(n12169) );
  ND4D1BWP30P140LVT U12753 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(n12183) );
  AOI22D1BWP30P140LVT U12754 ( .A1(i_data_bus[53]), .A2(n12370), .B1(
        i_data_bus[341]), .B2(n12369), .ZN(n12176) );
  AOI22D1BWP30P140LVT U12755 ( .A1(i_data_bus[949]), .A2(n12379), .B1(
        i_data_bus[981]), .B2(n12380), .ZN(n12175) );
  AOI22D1BWP30P140LVT U12756 ( .A1(i_data_bus[597]), .A2(n12368), .B1(
        i_data_bus[309]), .B2(n12378), .ZN(n12174) );
  AOI22D1BWP30P140LVT U12757 ( .A1(i_data_bus[565]), .A2(n12381), .B1(
        i_data_bus[437]), .B2(n12377), .ZN(n12173) );
  ND4D1BWP30P140LVT U12758 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(n12182) );
  AOI22D1BWP30P140LVT U12759 ( .A1(i_data_bus[789]), .A2(n12406), .B1(
        i_data_bus[725]), .B2(n12402), .ZN(n12180) );
  AOI22D1BWP30P140LVT U12760 ( .A1(i_data_bus[821]), .A2(n12403), .B1(
        i_data_bus[693]), .B2(n12407), .ZN(n12179) );
  AOI22D1BWP30P140LVT U12761 ( .A1(i_data_bus[757]), .A2(n12405), .B1(
        i_data_bus[853]), .B2(n12408), .ZN(n12178) );
  AOI22D1BWP30P140LVT U12762 ( .A1(i_data_bus[661]), .A2(n12404), .B1(
        i_data_bus[885]), .B2(n12401), .ZN(n12177) );
  ND4D1BWP30P140LVT U12763 ( .A1(n12180), .A2(n12179), .A3(n12178), .A4(n12177), .ZN(n12181) );
  OR4D1BWP30P140LVT U12764 ( .A1(n12184), .A2(n12183), .A3(n12182), .A4(n12181), .Z(o_data_bus[117]) );
  AOI22D1BWP30P140LVT U12765 ( .A1(i_data_bus[502]), .A2(n12390), .B1(
        i_data_bus[214]), .B2(n12372), .ZN(n12188) );
  AOI22D1BWP30P140LVT U12766 ( .A1(i_data_bus[406]), .A2(n12365), .B1(
        i_data_bus[342]), .B2(n12369), .ZN(n12187) );
  AOI22D1BWP30P140LVT U12767 ( .A1(i_data_bus[150]), .A2(n12395), .B1(
        i_data_bus[278]), .B2(n12389), .ZN(n12186) );
  AOI22D1BWP30P140LVT U12768 ( .A1(i_data_bus[630]), .A2(n12366), .B1(
        i_data_bus[982]), .B2(n12380), .ZN(n12185) );
  ND4D1BWP30P140LVT U12769 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(n12204) );
  AOI22D1BWP30P140LVT U12770 ( .A1(i_data_bus[118]), .A2(n12396), .B1(
        i_data_bus[950]), .B2(n12379), .ZN(n12192) );
  AOI22D1BWP30P140LVT U12771 ( .A1(i_data_bus[598]), .A2(n12368), .B1(
        i_data_bus[86]), .B2(n12382), .ZN(n12191) );
  AOI22D1BWP30P140LVT U12772 ( .A1(i_data_bus[1014]), .A2(n12394), .B1(
        i_data_bus[534]), .B2(n12384), .ZN(n12190) );
  AOI22D1BWP30P140LVT U12773 ( .A1(i_data_bus[566]), .A2(n12381), .B1(
        i_data_bus[374]), .B2(n12383), .ZN(n12189) );
  ND4D1BWP30P140LVT U12774 ( .A1(n12192), .A2(n12191), .A3(n12190), .A4(n12189), .ZN(n12203) );
  AOI22D1BWP30P140LVT U12775 ( .A1(i_data_bus[54]), .A2(n12370), .B1(
        i_data_bus[438]), .B2(n12377), .ZN(n12196) );
  AOI22D1BWP30P140LVT U12776 ( .A1(i_data_bus[22]), .A2(n12393), .B1(
        i_data_bus[470]), .B2(n12391), .ZN(n12195) );
  AOI22D1BWP30P140LVT U12777 ( .A1(i_data_bus[246]), .A2(n12367), .B1(
        i_data_bus[182]), .B2(n12371), .ZN(n12194) );
  AOI22D1BWP30P140LVT U12778 ( .A1(i_data_bus[918]), .A2(n12392), .B1(
        i_data_bus[310]), .B2(n12378), .ZN(n12193) );
  ND4D1BWP30P140LVT U12779 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(n12202) );
  AOI22D1BWP30P140LVT U12780 ( .A1(i_data_bus[694]), .A2(n12407), .B1(
        i_data_bus[758]), .B2(n12405), .ZN(n12200) );
  AOI22D1BWP30P140LVT U12781 ( .A1(i_data_bus[726]), .A2(n12402), .B1(
        i_data_bus[854]), .B2(n12408), .ZN(n12199) );
  AOI22D1BWP30P140LVT U12782 ( .A1(i_data_bus[886]), .A2(n12401), .B1(
        i_data_bus[662]), .B2(n12404), .ZN(n12198) );
  AOI22D1BWP30P140LVT U12783 ( .A1(i_data_bus[822]), .A2(n12403), .B1(
        i_data_bus[790]), .B2(n12406), .ZN(n12197) );
  ND4D1BWP30P140LVT U12784 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(n12201) );
  OR4D1BWP30P140LVT U12785 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .Z(o_data_bus[118]) );
  AOI22D1BWP30P140LVT U12786 ( .A1(i_data_bus[471]), .A2(n12391), .B1(
        i_data_bus[439]), .B2(n12377), .ZN(n12208) );
  AOI22D1BWP30P140LVT U12787 ( .A1(i_data_bus[311]), .A2(n12378), .B1(
        i_data_bus[279]), .B2(n12389), .ZN(n12207) );
  AOI22D1BWP30P140LVT U12788 ( .A1(i_data_bus[1015]), .A2(n12394), .B1(
        i_data_bus[87]), .B2(n12382), .ZN(n12206) );
  AOI22D1BWP30P140LVT U12789 ( .A1(i_data_bus[599]), .A2(n12368), .B1(
        i_data_bus[343]), .B2(n12369), .ZN(n12205) );
  ND4D1BWP30P140LVT U12790 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(n12224) );
  AOI22D1BWP30P140LVT U12791 ( .A1(i_data_bus[247]), .A2(n12367), .B1(
        i_data_bus[375]), .B2(n12383), .ZN(n12212) );
  AOI22D1BWP30P140LVT U12792 ( .A1(i_data_bus[119]), .A2(n12396), .B1(
        i_data_bus[567]), .B2(n12381), .ZN(n12211) );
  AOI22D1BWP30P140LVT U12793 ( .A1(i_data_bus[151]), .A2(n12395), .B1(
        i_data_bus[407]), .B2(n12365), .ZN(n12210) );
  AOI22D1BWP30P140LVT U12794 ( .A1(i_data_bus[951]), .A2(n12379), .B1(
        i_data_bus[919]), .B2(n12392), .ZN(n12209) );
  ND4D1BWP30P140LVT U12795 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(n12223) );
  AOI22D1BWP30P140LVT U12796 ( .A1(i_data_bus[23]), .A2(n12393), .B1(
        i_data_bus[535]), .B2(n12384), .ZN(n12216) );
  AOI22D1BWP30P140LVT U12797 ( .A1(i_data_bus[983]), .A2(n12380), .B1(
        i_data_bus[215]), .B2(n12372), .ZN(n12215) );
  AOI22D1BWP30P140LVT U12798 ( .A1(i_data_bus[631]), .A2(n12366), .B1(
        i_data_bus[183]), .B2(n12371), .ZN(n12214) );
  AOI22D1BWP30P140LVT U12799 ( .A1(i_data_bus[55]), .A2(n12370), .B1(
        i_data_bus[503]), .B2(n12390), .ZN(n12213) );
  ND4D1BWP30P140LVT U12800 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(n12222) );
  AOI22D1BWP30P140LVT U12801 ( .A1(i_data_bus[887]), .A2(n12401), .B1(
        i_data_bus[663]), .B2(n12404), .ZN(n12220) );
  AOI22D1BWP30P140LVT U12802 ( .A1(i_data_bus[759]), .A2(n12405), .B1(
        i_data_bus[855]), .B2(n12408), .ZN(n12219) );
  AOI22D1BWP30P140LVT U12803 ( .A1(i_data_bus[727]), .A2(n12402), .B1(
        i_data_bus[823]), .B2(n12403), .ZN(n12218) );
  AOI22D1BWP30P140LVT U12804 ( .A1(i_data_bus[695]), .A2(n12407), .B1(
        i_data_bus[791]), .B2(n12406), .ZN(n12217) );
  ND4D1BWP30P140LVT U12805 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(n12221) );
  OR4D1BWP30P140LVT U12806 ( .A1(n12224), .A2(n12223), .A3(n12222), .A4(n12221), .Z(o_data_bus[119]) );
  AOI22D1BWP30P140LVT U12807 ( .A1(i_data_bus[600]), .A2(n12368), .B1(
        i_data_bus[952]), .B2(n12379), .ZN(n12228) );
  AOI22D1BWP30P140LVT U12808 ( .A1(i_data_bus[536]), .A2(n12384), .B1(
        i_data_bus[248]), .B2(n12367), .ZN(n12227) );
  AOI22D1BWP30P140LVT U12809 ( .A1(i_data_bus[920]), .A2(n12392), .B1(
        i_data_bus[376]), .B2(n12383), .ZN(n12226) );
  AOI22D1BWP30P140LVT U12810 ( .A1(i_data_bus[88]), .A2(n12382), .B1(
        i_data_bus[344]), .B2(n12369), .ZN(n12225) );
  ND4D1BWP30P140LVT U12811 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(n12244) );
  AOI22D1BWP30P140LVT U12812 ( .A1(i_data_bus[56]), .A2(n12370), .B1(
        i_data_bus[216]), .B2(n12372), .ZN(n12232) );
  AOI22D1BWP30P140LVT U12813 ( .A1(i_data_bus[440]), .A2(n12377), .B1(
        i_data_bus[152]), .B2(n12395), .ZN(n12231) );
  AOI22D1BWP30P140LVT U12814 ( .A1(i_data_bus[280]), .A2(n12389), .B1(
        i_data_bus[504]), .B2(n12390), .ZN(n12230) );
  AOI22D1BWP30P140LVT U12815 ( .A1(i_data_bus[1016]), .A2(n12394), .B1(
        i_data_bus[184]), .B2(n12371), .ZN(n12229) );
  ND4D1BWP30P140LVT U12816 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(n12243) );
  AOI22D1BWP30P140LVT U12817 ( .A1(i_data_bus[24]), .A2(n12393), .B1(
        i_data_bus[568]), .B2(n12381), .ZN(n12236) );
  AOI22D1BWP30P140LVT U12818 ( .A1(i_data_bus[984]), .A2(n12380), .B1(
        i_data_bus[472]), .B2(n12391), .ZN(n12235) );
  AOI22D1BWP30P140LVT U12819 ( .A1(i_data_bus[632]), .A2(n12366), .B1(
        i_data_bus[408]), .B2(n12365), .ZN(n12234) );
  AOI22D1BWP30P140LVT U12820 ( .A1(i_data_bus[120]), .A2(n12396), .B1(
        i_data_bus[312]), .B2(n12378), .ZN(n12233) );
  ND4D1BWP30P140LVT U12821 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(n12242) );
  AOI22D1BWP30P140LVT U12822 ( .A1(i_data_bus[824]), .A2(n12403), .B1(
        i_data_bus[760]), .B2(n12405), .ZN(n12240) );
  AOI22D1BWP30P140LVT U12823 ( .A1(i_data_bus[856]), .A2(n12408), .B1(
        i_data_bus[664]), .B2(n12404), .ZN(n12239) );
  AOI22D1BWP30P140LVT U12824 ( .A1(i_data_bus[728]), .A2(n12402), .B1(
        i_data_bus[888]), .B2(n12401), .ZN(n12238) );
  AOI22D1BWP30P140LVT U12825 ( .A1(i_data_bus[792]), .A2(n12406), .B1(
        i_data_bus[696]), .B2(n12407), .ZN(n12237) );
  ND4D1BWP30P140LVT U12826 ( .A1(n12240), .A2(n12239), .A3(n12238), .A4(n12237), .ZN(n12241) );
  OR4D1BWP30P140LVT U12827 ( .A1(n12244), .A2(n12243), .A3(n12242), .A4(n12241), .Z(o_data_bus[120]) );
  AOI22D1BWP30P140LVT U12828 ( .A1(i_data_bus[281]), .A2(n12389), .B1(
        i_data_bus[249]), .B2(n12367), .ZN(n12248) );
  AOI22D1BWP30P140LVT U12829 ( .A1(i_data_bus[345]), .A2(n12369), .B1(
        i_data_bus[441]), .B2(n12377), .ZN(n12247) );
  AOI22D1BWP30P140LVT U12830 ( .A1(i_data_bus[1017]), .A2(n12394), .B1(
        i_data_bus[313]), .B2(n12378), .ZN(n12246) );
  AOI22D1BWP30P140LVT U12831 ( .A1(i_data_bus[921]), .A2(n12392), .B1(
        i_data_bus[121]), .B2(n12396), .ZN(n12245) );
  ND4D1BWP30P140LVT U12832 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(n12264) );
  AOI22D1BWP30P140LVT U12833 ( .A1(i_data_bus[89]), .A2(n12382), .B1(
        i_data_bus[217]), .B2(n12372), .ZN(n12252) );
  AOI22D1BWP30P140LVT U12834 ( .A1(i_data_bus[953]), .A2(n12379), .B1(
        i_data_bus[185]), .B2(n12371), .ZN(n12251) );
  AOI22D1BWP30P140LVT U12835 ( .A1(i_data_bus[57]), .A2(n12370), .B1(
        i_data_bus[601]), .B2(n12368), .ZN(n12250) );
  AOI22D1BWP30P140LVT U12836 ( .A1(i_data_bus[537]), .A2(n12384), .B1(
        i_data_bus[153]), .B2(n12395), .ZN(n12249) );
  ND4D1BWP30P140LVT U12837 ( .A1(n12252), .A2(n12251), .A3(n12250), .A4(n12249), .ZN(n12263) );
  AOI22D1BWP30P140LVT U12838 ( .A1(i_data_bus[377]), .A2(n12383), .B1(
        i_data_bus[505]), .B2(n12390), .ZN(n12256) );
  AOI22D1BWP30P140LVT U12839 ( .A1(i_data_bus[633]), .A2(n12366), .B1(
        i_data_bus[473]), .B2(n12391), .ZN(n12255) );
  AOI22D1BWP30P140LVT U12840 ( .A1(i_data_bus[985]), .A2(n12380), .B1(
        i_data_bus[25]), .B2(n12393), .ZN(n12254) );
  AOI22D1BWP30P140LVT U12841 ( .A1(i_data_bus[569]), .A2(n12381), .B1(
        i_data_bus[409]), .B2(n12365), .ZN(n12253) );
  ND4D1BWP30P140LVT U12842 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12253), .ZN(n12262) );
  AOI22D1BWP30P140LVT U12843 ( .A1(i_data_bus[825]), .A2(n12403), .B1(
        i_data_bus[793]), .B2(n12406), .ZN(n12260) );
  AOI22D1BWP30P140LVT U12844 ( .A1(i_data_bus[761]), .A2(n12405), .B1(
        i_data_bus[857]), .B2(n12408), .ZN(n12259) );
  AOI22D1BWP30P140LVT U12845 ( .A1(i_data_bus[729]), .A2(n12402), .B1(
        i_data_bus[665]), .B2(n12404), .ZN(n12258) );
  AOI22D1BWP30P140LVT U12846 ( .A1(i_data_bus[697]), .A2(n12407), .B1(
        i_data_bus[889]), .B2(n12401), .ZN(n12257) );
  ND4D1BWP30P140LVT U12847 ( .A1(n12260), .A2(n12259), .A3(n12258), .A4(n12257), .ZN(n12261) );
  OR4D1BWP30P140LVT U12848 ( .A1(n12264), .A2(n12263), .A3(n12262), .A4(n12261), .Z(o_data_bus[121]) );
  AOI22D1BWP30P140LVT U12849 ( .A1(i_data_bus[634]), .A2(n12366), .B1(
        i_data_bus[314]), .B2(n12378), .ZN(n12268) );
  AOI22D1BWP30P140LVT U12850 ( .A1(i_data_bus[954]), .A2(n12379), .B1(
        i_data_bus[506]), .B2(n12390), .ZN(n12267) );
  AOI22D1BWP30P140LVT U12851 ( .A1(i_data_bus[442]), .A2(n12377), .B1(
        i_data_bus[378]), .B2(n12383), .ZN(n12266) );
  AOI22D1BWP30P140LVT U12852 ( .A1(i_data_bus[570]), .A2(n12381), .B1(
        i_data_bus[218]), .B2(n12372), .ZN(n12265) );
  ND4D1BWP30P140LVT U12853 ( .A1(n12268), .A2(n12267), .A3(n12266), .A4(n12265), .ZN(n12284) );
  AOI22D1BWP30P140LVT U12854 ( .A1(i_data_bus[90]), .A2(n12382), .B1(
        i_data_bus[474]), .B2(n12391), .ZN(n12272) );
  AOI22D1BWP30P140LVT U12855 ( .A1(i_data_bus[122]), .A2(n12396), .B1(
        i_data_bus[538]), .B2(n12384), .ZN(n12271) );
  AOI22D1BWP30P140LVT U12856 ( .A1(i_data_bus[602]), .A2(n12368), .B1(
        i_data_bus[986]), .B2(n12380), .ZN(n12270) );
  AOI22D1BWP30P140LVT U12857 ( .A1(i_data_bus[58]), .A2(n12370), .B1(
        i_data_bus[186]), .B2(n12371), .ZN(n12269) );
  ND4D1BWP30P140LVT U12858 ( .A1(n12272), .A2(n12271), .A3(n12270), .A4(n12269), .ZN(n12283) );
  AOI22D1BWP30P140LVT U12859 ( .A1(i_data_bus[26]), .A2(n12393), .B1(
        i_data_bus[346]), .B2(n12369), .ZN(n12276) );
  AOI22D1BWP30P140LVT U12860 ( .A1(i_data_bus[922]), .A2(n12392), .B1(
        i_data_bus[282]), .B2(n12389), .ZN(n12275) );
  AOI22D1BWP30P140LVT U12861 ( .A1(i_data_bus[1018]), .A2(n12394), .B1(
        i_data_bus[154]), .B2(n12395), .ZN(n12274) );
  AOI22D1BWP30P140LVT U12862 ( .A1(i_data_bus[250]), .A2(n12367), .B1(
        i_data_bus[410]), .B2(n12365), .ZN(n12273) );
  ND4D1BWP30P140LVT U12863 ( .A1(n12276), .A2(n12275), .A3(n12274), .A4(n12273), .ZN(n12282) );
  AOI22D1BWP30P140LVT U12864 ( .A1(i_data_bus[858]), .A2(n12408), .B1(
        i_data_bus[762]), .B2(n12405), .ZN(n12280) );
  AOI22D1BWP30P140LVT U12865 ( .A1(i_data_bus[826]), .A2(n12403), .B1(
        i_data_bus[730]), .B2(n12402), .ZN(n12279) );
  AOI22D1BWP30P140LVT U12866 ( .A1(i_data_bus[890]), .A2(n12401), .B1(
        i_data_bus[698]), .B2(n12407), .ZN(n12278) );
  AOI22D1BWP30P140LVT U12867 ( .A1(i_data_bus[794]), .A2(n12406), .B1(
        i_data_bus[666]), .B2(n12404), .ZN(n12277) );
  ND4D1BWP30P140LVT U12868 ( .A1(n12280), .A2(n12279), .A3(n12278), .A4(n12277), .ZN(n12281) );
  OR4D1BWP30P140LVT U12869 ( .A1(n12284), .A2(n12283), .A3(n12282), .A4(n12281), .Z(o_data_bus[122]) );
  AOI22D1BWP30P140LVT U12870 ( .A1(i_data_bus[603]), .A2(n12368), .B1(
        i_data_bus[923]), .B2(n12392), .ZN(n12288) );
  AOI22D1BWP30P140LVT U12871 ( .A1(i_data_bus[411]), .A2(n12365), .B1(
        i_data_bus[283]), .B2(n12389), .ZN(n12287) );
  AOI22D1BWP30P140LVT U12872 ( .A1(i_data_bus[123]), .A2(n12396), .B1(
        i_data_bus[475]), .B2(n12391), .ZN(n12286) );
  AOI22D1BWP30P140LVT U12873 ( .A1(i_data_bus[987]), .A2(n12380), .B1(
        i_data_bus[347]), .B2(n12369), .ZN(n12285) );
  ND4D1BWP30P140LVT U12874 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(n12304) );
  AOI22D1BWP30P140LVT U12875 ( .A1(i_data_bus[635]), .A2(n12366), .B1(
        i_data_bus[219]), .B2(n12372), .ZN(n12292) );
  AOI22D1BWP30P140LVT U12876 ( .A1(i_data_bus[1019]), .A2(n12394), .B1(
        i_data_bus[155]), .B2(n12395), .ZN(n12291) );
  AOI22D1BWP30P140LVT U12877 ( .A1(i_data_bus[91]), .A2(n12382), .B1(
        i_data_bus[379]), .B2(n12383), .ZN(n12290) );
  AOI22D1BWP30P140LVT U12878 ( .A1(i_data_bus[571]), .A2(n12381), .B1(
        i_data_bus[443]), .B2(n12377), .ZN(n12289) );
  ND4D1BWP30P140LVT U12879 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(n12303) );
  AOI22D1BWP30P140LVT U12880 ( .A1(i_data_bus[27]), .A2(n12393), .B1(
        i_data_bus[59]), .B2(n12370), .ZN(n12296) );
  AOI22D1BWP30P140LVT U12881 ( .A1(i_data_bus[539]), .A2(n12384), .B1(
        i_data_bus[955]), .B2(n12379), .ZN(n12295) );
  AOI22D1BWP30P140LVT U12882 ( .A1(i_data_bus[507]), .A2(n12390), .B1(
        i_data_bus[187]), .B2(n12371), .ZN(n12294) );
  AOI22D1BWP30P140LVT U12883 ( .A1(i_data_bus[315]), .A2(n12378), .B1(
        i_data_bus[251]), .B2(n12367), .ZN(n12293) );
  ND4D1BWP30P140LVT U12884 ( .A1(n12296), .A2(n12295), .A3(n12294), .A4(n12293), .ZN(n12302) );
  AOI22D1BWP30P140LVT U12885 ( .A1(i_data_bus[827]), .A2(n12403), .B1(
        i_data_bus[763]), .B2(n12405), .ZN(n12300) );
  AOI22D1BWP30P140LVT U12886 ( .A1(i_data_bus[731]), .A2(n12402), .B1(
        i_data_bus[699]), .B2(n12407), .ZN(n12299) );
  AOI22D1BWP30P140LVT U12887 ( .A1(i_data_bus[891]), .A2(n12401), .B1(
        i_data_bus[667]), .B2(n12404), .ZN(n12298) );
  AOI22D1BWP30P140LVT U12888 ( .A1(i_data_bus[795]), .A2(n12406), .B1(
        i_data_bus[859]), .B2(n12408), .ZN(n12297) );
  ND4D1BWP30P140LVT U12889 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(n12301) );
  OR4D1BWP30P140LVT U12890 ( .A1(n12304), .A2(n12303), .A3(n12302), .A4(n12301), .Z(o_data_bus[123]) );
  AOI22D1BWP30P140LVT U12891 ( .A1(i_data_bus[124]), .A2(n12396), .B1(
        i_data_bus[1020]), .B2(n12394), .ZN(n12308) );
  AOI22D1BWP30P140LVT U12892 ( .A1(i_data_bus[636]), .A2(n12366), .B1(
        i_data_bus[444]), .B2(n12377), .ZN(n12307) );
  AOI22D1BWP30P140LVT U12893 ( .A1(i_data_bus[92]), .A2(n12382), .B1(
        i_data_bus[28]), .B2(n12393), .ZN(n12306) );
  AOI22D1BWP30P140LVT U12894 ( .A1(i_data_bus[988]), .A2(n12380), .B1(
        i_data_bus[316]), .B2(n12378), .ZN(n12305) );
  ND4D1BWP30P140LVT U12895 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(n12324) );
  AOI22D1BWP30P140LVT U12896 ( .A1(i_data_bus[572]), .A2(n12381), .B1(
        i_data_bus[380]), .B2(n12383), .ZN(n12312) );
  AOI22D1BWP30P140LVT U12897 ( .A1(i_data_bus[956]), .A2(n12379), .B1(
        i_data_bus[412]), .B2(n12365), .ZN(n12311) );
  AOI22D1BWP30P140LVT U12898 ( .A1(i_data_bus[60]), .A2(n12370), .B1(
        i_data_bus[188]), .B2(n12371), .ZN(n12310) );
  AOI22D1BWP30P140LVT U12899 ( .A1(i_data_bus[252]), .A2(n12367), .B1(
        i_data_bus[284]), .B2(n12389), .ZN(n12309) );
  ND4D1BWP30P140LVT U12900 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(n12323) );
  AOI22D1BWP30P140LVT U12901 ( .A1(i_data_bus[156]), .A2(n12395), .B1(
        i_data_bus[220]), .B2(n12372), .ZN(n12316) );
  AOI22D1BWP30P140LVT U12902 ( .A1(i_data_bus[540]), .A2(n12384), .B1(
        i_data_bus[348]), .B2(n12369), .ZN(n12315) );
  AOI22D1BWP30P140LVT U12903 ( .A1(i_data_bus[924]), .A2(n12392), .B1(
        i_data_bus[476]), .B2(n12391), .ZN(n12314) );
  AOI22D1BWP30P140LVT U12904 ( .A1(i_data_bus[604]), .A2(n12368), .B1(
        i_data_bus[508]), .B2(n12390), .ZN(n12313) );
  ND4D1BWP30P140LVT U12905 ( .A1(n12316), .A2(n12315), .A3(n12314), .A4(n12313), .ZN(n12322) );
  AOI22D1BWP30P140LVT U12906 ( .A1(i_data_bus[764]), .A2(n12405), .B1(
        i_data_bus[860]), .B2(n12408), .ZN(n12320) );
  AOI22D1BWP30P140LVT U12907 ( .A1(i_data_bus[796]), .A2(n12406), .B1(
        i_data_bus[828]), .B2(n12403), .ZN(n12319) );
  AOI22D1BWP30P140LVT U12908 ( .A1(i_data_bus[892]), .A2(n12401), .B1(
        i_data_bus[700]), .B2(n12407), .ZN(n12318) );
  AOI22D1BWP30P140LVT U12909 ( .A1(i_data_bus[732]), .A2(n12402), .B1(
        i_data_bus[668]), .B2(n12404), .ZN(n12317) );
  ND4D1BWP30P140LVT U12910 ( .A1(n12320), .A2(n12319), .A3(n12318), .A4(n12317), .ZN(n12321) );
  OR4D1BWP30P140LVT U12911 ( .A1(n12324), .A2(n12323), .A3(n12322), .A4(n12321), .Z(o_data_bus[124]) );
  AOI22D1BWP30P140LVT U12912 ( .A1(i_data_bus[93]), .A2(n12382), .B1(
        i_data_bus[189]), .B2(n12371), .ZN(n12328) );
  AOI22D1BWP30P140LVT U12913 ( .A1(i_data_bus[29]), .A2(n12393), .B1(
        i_data_bus[477]), .B2(n12391), .ZN(n12327) );
  AOI22D1BWP30P140LVT U12914 ( .A1(i_data_bus[125]), .A2(n12396), .B1(
        i_data_bus[157]), .B2(n12395), .ZN(n12326) );
  AOI22D1BWP30P140LVT U12915 ( .A1(i_data_bus[637]), .A2(n12366), .B1(
        i_data_bus[221]), .B2(n12372), .ZN(n12325) );
  ND4D1BWP30P140LVT U12916 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(n12344) );
  AOI22D1BWP30P140LVT U12917 ( .A1(i_data_bus[573]), .A2(n12381), .B1(
        i_data_bus[1021]), .B2(n12394), .ZN(n12332) );
  AOI22D1BWP30P140LVT U12918 ( .A1(i_data_bus[989]), .A2(n12380), .B1(
        i_data_bus[285]), .B2(n12389), .ZN(n12331) );
  AOI22D1BWP30P140LVT U12919 ( .A1(i_data_bus[349]), .A2(n12369), .B1(
        i_data_bus[253]), .B2(n12367), .ZN(n12330) );
  AOI22D1BWP30P140LVT U12920 ( .A1(i_data_bus[605]), .A2(n12368), .B1(
        i_data_bus[317]), .B2(n12378), .ZN(n12329) );
  ND4D1BWP30P140LVT U12921 ( .A1(n12332), .A2(n12331), .A3(n12330), .A4(n12329), .ZN(n12343) );
  AOI22D1BWP30P140LVT U12922 ( .A1(i_data_bus[61]), .A2(n12370), .B1(
        i_data_bus[413]), .B2(n12365), .ZN(n12336) );
  AOI22D1BWP30P140LVT U12923 ( .A1(i_data_bus[445]), .A2(n12377), .B1(
        i_data_bus[509]), .B2(n12390), .ZN(n12335) );
  AOI22D1BWP30P140LVT U12924 ( .A1(i_data_bus[957]), .A2(n12379), .B1(
        i_data_bus[541]), .B2(n12384), .ZN(n12334) );
  AOI22D1BWP30P140LVT U12925 ( .A1(i_data_bus[925]), .A2(n12392), .B1(
        i_data_bus[381]), .B2(n12383), .ZN(n12333) );
  ND4D1BWP30P140LVT U12926 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(n12342) );
  AOI22D1BWP30P140LVT U12927 ( .A1(i_data_bus[669]), .A2(n12404), .B1(
        i_data_bus[797]), .B2(n12406), .ZN(n12340) );
  AOI22D1BWP30P140LVT U12928 ( .A1(i_data_bus[829]), .A2(n12403), .B1(
        i_data_bus[861]), .B2(n12408), .ZN(n12339) );
  AOI22D1BWP30P140LVT U12929 ( .A1(i_data_bus[765]), .A2(n12405), .B1(
        i_data_bus[733]), .B2(n12402), .ZN(n12338) );
  AOI22D1BWP30P140LVT U12930 ( .A1(i_data_bus[701]), .A2(n12407), .B1(
        i_data_bus[893]), .B2(n12401), .ZN(n12337) );
  ND4D1BWP30P140LVT U12931 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(n12341) );
  OR4D1BWP30P140LVT U12932 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12341), .Z(o_data_bus[125]) );
  AOI22D1BWP30P140LVT U12933 ( .A1(i_data_bus[958]), .A2(n12379), .B1(
        i_data_bus[606]), .B2(n12368), .ZN(n12348) );
  AOI22D1BWP30P140LVT U12934 ( .A1(i_data_bus[62]), .A2(n12370), .B1(
        i_data_bus[574]), .B2(n12381), .ZN(n12347) );
  AOI22D1BWP30P140LVT U12935 ( .A1(i_data_bus[126]), .A2(n12396), .B1(
        i_data_bus[478]), .B2(n12391), .ZN(n12346) );
  AOI22D1BWP30P140LVT U12936 ( .A1(i_data_bus[638]), .A2(n12366), .B1(
        i_data_bus[446]), .B2(n12377), .ZN(n12345) );
  ND4D1BWP30P140LVT U12937 ( .A1(n12348), .A2(n12347), .A3(n12346), .A4(n12345), .ZN(n12364) );
  AOI22D1BWP30P140LVT U12938 ( .A1(i_data_bus[542]), .A2(n12384), .B1(
        i_data_bus[382]), .B2(n12383), .ZN(n12352) );
  AOI22D1BWP30P140LVT U12939 ( .A1(i_data_bus[222]), .A2(n12372), .B1(
        i_data_bus[510]), .B2(n12390), .ZN(n12351) );
  AOI22D1BWP30P140LVT U12940 ( .A1(i_data_bus[30]), .A2(n12393), .B1(
        i_data_bus[158]), .B2(n12395), .ZN(n12350) );
  AOI22D1BWP30P140LVT U12941 ( .A1(i_data_bus[990]), .A2(n12380), .B1(
        i_data_bus[350]), .B2(n12369), .ZN(n12349) );
  ND4D1BWP30P140LVT U12942 ( .A1(n12352), .A2(n12351), .A3(n12350), .A4(n12349), .ZN(n12363) );
  AOI22D1BWP30P140LVT U12943 ( .A1(i_data_bus[318]), .A2(n12378), .B1(
        i_data_bus[190]), .B2(n12371), .ZN(n12356) );
  AOI22D1BWP30P140LVT U12944 ( .A1(i_data_bus[1022]), .A2(n12394), .B1(
        i_data_bus[254]), .B2(n12367), .ZN(n12355) );
  AOI22D1BWP30P140LVT U12945 ( .A1(i_data_bus[94]), .A2(n12382), .B1(
        i_data_bus[286]), .B2(n12389), .ZN(n12354) );
  AOI22D1BWP30P140LVT U12946 ( .A1(i_data_bus[926]), .A2(n12392), .B1(
        i_data_bus[414]), .B2(n12365), .ZN(n12353) );
  ND4D1BWP30P140LVT U12947 ( .A1(n12356), .A2(n12355), .A3(n12354), .A4(n12353), .ZN(n12362) );
  AOI22D1BWP30P140LVT U12948 ( .A1(i_data_bus[670]), .A2(n12404), .B1(
        i_data_bus[894]), .B2(n12401), .ZN(n12360) );
  AOI22D1BWP30P140LVT U12949 ( .A1(i_data_bus[798]), .A2(n12406), .B1(
        i_data_bus[830]), .B2(n12403), .ZN(n12359) );
  AOI22D1BWP30P140LVT U12950 ( .A1(i_data_bus[766]), .A2(n12405), .B1(
        i_data_bus[702]), .B2(n12407), .ZN(n12358) );
  AOI22D1BWP30P140LVT U12951 ( .A1(i_data_bus[862]), .A2(n12408), .B1(
        i_data_bus[734]), .B2(n12402), .ZN(n12357) );
  ND4D1BWP30P140LVT U12952 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12357), .ZN(n12361) );
  OR4D1BWP30P140LVT U12953 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .Z(o_data_bus[126]) );
  AOI22D1BWP30P140LVT U12954 ( .A1(i_data_bus[639]), .A2(n12366), .B1(
        i_data_bus[415]), .B2(n12365), .ZN(n12376) );
  AOI22D1BWP30P140LVT U12955 ( .A1(i_data_bus[607]), .A2(n12368), .B1(
        i_data_bus[255]), .B2(n12367), .ZN(n12375) );
  AOI22D1BWP30P140LVT U12956 ( .A1(i_data_bus[63]), .A2(n12370), .B1(
        i_data_bus[351]), .B2(n12369), .ZN(n12374) );
  AOI22D1BWP30P140LVT U12957 ( .A1(i_data_bus[223]), .A2(n12372), .B1(
        i_data_bus[191]), .B2(n12371), .ZN(n12373) );
  ND4D1BWP30P140LVT U12958 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(n12416) );
  AOI22D1BWP30P140LVT U12959 ( .A1(i_data_bus[319]), .A2(n12378), .B1(
        i_data_bus[447]), .B2(n12377), .ZN(n12388) );
  AOI22D1BWP30P140LVT U12960 ( .A1(i_data_bus[991]), .A2(n12380), .B1(
        i_data_bus[959]), .B2(n12379), .ZN(n12387) );
  AOI22D1BWP30P140LVT U12961 ( .A1(i_data_bus[95]), .A2(n12382), .B1(
        i_data_bus[575]), .B2(n12381), .ZN(n12386) );
  AOI22D1BWP30P140LVT U12962 ( .A1(i_data_bus[543]), .A2(n12384), .B1(
        i_data_bus[383]), .B2(n12383), .ZN(n12385) );
  ND4D1BWP30P140LVT U12963 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n12385), .ZN(n12415) );
  AOI22D1BWP30P140LVT U12964 ( .A1(i_data_bus[511]), .A2(n12390), .B1(
        i_data_bus[287]), .B2(n12389), .ZN(n12400) );
  AOI22D1BWP30P140LVT U12965 ( .A1(i_data_bus[927]), .A2(n12392), .B1(
        i_data_bus[479]), .B2(n12391), .ZN(n12399) );
  AOI22D1BWP30P140LVT U12966 ( .A1(i_data_bus[1023]), .A2(n12394), .B1(
        i_data_bus[31]), .B2(n12393), .ZN(n12398) );
  AOI22D1BWP30P140LVT U12967 ( .A1(i_data_bus[127]), .A2(n12396), .B1(
        i_data_bus[159]), .B2(n12395), .ZN(n12397) );
  ND4D1BWP30P140LVT U12968 ( .A1(n12400), .A2(n12399), .A3(n12398), .A4(n12397), .ZN(n12414) );
  AOI22D1BWP30P140LVT U12969 ( .A1(i_data_bus[735]), .A2(n12402), .B1(
        i_data_bus[895]), .B2(n12401), .ZN(n12412) );
  AOI22D1BWP30P140LVT U12970 ( .A1(i_data_bus[671]), .A2(n12404), .B1(
        i_data_bus[831]), .B2(n12403), .ZN(n12411) );
  AOI22D1BWP30P140LVT U12971 ( .A1(i_data_bus[799]), .A2(n12406), .B1(
        i_data_bus[767]), .B2(n12405), .ZN(n12410) );
  AOI22D1BWP30P140LVT U12972 ( .A1(i_data_bus[863]), .A2(n12408), .B1(
        i_data_bus[703]), .B2(n12407), .ZN(n12409) );
  ND4D1BWP30P140LVT U12973 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12409), .ZN(n12413) );
  OR4D1BWP30P140LVT U12974 ( .A1(n12416), .A2(n12415), .A3(n12414), .A4(n12413), .Z(o_data_bus[127]) );
  AOI22D1BWP30P140LVT U12975 ( .A1(i_data_bus[960]), .A2(n12482), .B1(
        i_data_bus[128]), .B2(n12502), .ZN(n12420) );
  AOI22D1BWP30P140LVT U12976 ( .A1(i_data_bus[544]), .A2(n12479), .B1(
        i_data_bus[608]), .B2(n12504), .ZN(n12419) );
  AOI22D1BWP30P140LVT U12977 ( .A1(i_data_bus[224]), .A2(n12493), .B1(
        i_data_bus[288]), .B2(n12505), .ZN(n12418) );
  AOI22D1BWP30P140LVT U12978 ( .A1(i_data_bus[480]), .A2(n12494), .B1(
        i_data_bus[416]), .B2(n12481), .ZN(n12417) );
  ND4D1BWP30P140LVT U12979 ( .A1(n12420), .A2(n12419), .A3(n12418), .A4(n12417), .ZN(n12436) );
  AOI22D1BWP30P140LVT U12980 ( .A1(i_data_bus[320]), .A2(n12508), .B1(
        i_data_bus[256]), .B2(n12503), .ZN(n12424) );
  AOI22D1BWP30P140LVT U12981 ( .A1(i_data_bus[384]), .A2(n12506), .B1(
        i_data_bus[448]), .B2(n12507), .ZN(n12423) );
  AOI22D1BWP30P140LVT U12982 ( .A1(i_data_bus[992]), .A2(n12496), .B1(
        i_data_bus[928]), .B2(n12492), .ZN(n12422) );
  AOI22D1BWP30P140LVT U12983 ( .A1(i_data_bus[0]), .A2(n12490), .B1(
        i_data_bus[64]), .B2(n12478), .ZN(n12421) );
  ND4D1BWP30P140LVT U12984 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(n12435) );
  AOI22D1BWP30P140LVT U12985 ( .A1(i_data_bus[512]), .A2(n12477), .B1(
        i_data_bus[192]), .B2(n12495), .ZN(n12428) );
  AOI22D1BWP30P140LVT U12986 ( .A1(i_data_bus[96]), .A2(n12489), .B1(
        i_data_bus[576]), .B2(n12480), .ZN(n12427) );
  AOI22D1BWP30P140LVT U12987 ( .A1(i_data_bus[32]), .A2(n12483), .B1(
        i_data_bus[352]), .B2(n12491), .ZN(n12426) );
  AOI22D1BWP30P140LVT U12988 ( .A1(i_data_bus[896]), .A2(n12484), .B1(
        i_data_bus[160]), .B2(n12501), .ZN(n12425) );
  ND4D1BWP30P140LVT U12989 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(n12434) );
  AOI22D1BWP30P140LVT U12990 ( .A1(i_data_bus[672]), .A2(n12515), .B1(
        i_data_bus[800]), .B2(n12517), .ZN(n12432) );
  AOI22D1BWP30P140LVT U12991 ( .A1(i_data_bus[768]), .A2(n12516), .B1(
        i_data_bus[864]), .B2(n12513), .ZN(n12431) );
  AOI22D1BWP30P140LVT U12992 ( .A1(i_data_bus[832]), .A2(n12514), .B1(
        i_data_bus[704]), .B2(n12519), .ZN(n12430) );
  AOI22D1BWP30P140LVT U12993 ( .A1(i_data_bus[640]), .A2(n12520), .B1(
        i_data_bus[736]), .B2(n12518), .ZN(n12429) );
  ND4D1BWP30P140LVT U12994 ( .A1(n12432), .A2(n12431), .A3(n12430), .A4(n12429), .ZN(n12433) );
  OR4D1BWP30P140LVT U12995 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n12433), .Z(o_data_bus[128]) );
  AOI22D1BWP30P140LVT U12996 ( .A1(i_data_bus[65]), .A2(n12478), .B1(
        i_data_bus[449]), .B2(n12507), .ZN(n12440) );
  AOI22D1BWP30P140LVT U12997 ( .A1(i_data_bus[33]), .A2(n12483), .B1(
        i_data_bus[161]), .B2(n12501), .ZN(n12439) );
  AOI22D1BWP30P140LVT U12998 ( .A1(i_data_bus[257]), .A2(n12503), .B1(
        i_data_bus[289]), .B2(n12505), .ZN(n12438) );
  AOI22D1BWP30P140LVT U12999 ( .A1(i_data_bus[609]), .A2(n12504), .B1(
        i_data_bus[1]), .B2(n12490), .ZN(n12437) );
  ND4D1BWP30P140LVT U13000 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(n12456) );
  AOI22D1BWP30P140LVT U13001 ( .A1(i_data_bus[225]), .A2(n12493), .B1(
        i_data_bus[129]), .B2(n12502), .ZN(n12444) );
  AOI22D1BWP30P140LVT U13002 ( .A1(i_data_bus[545]), .A2(n12479), .B1(
        i_data_bus[193]), .B2(n12495), .ZN(n12443) );
  AOI22D1BWP30P140LVT U13003 ( .A1(i_data_bus[577]), .A2(n12480), .B1(
        i_data_bus[321]), .B2(n12508), .ZN(n12442) );
  AOI22D1BWP30P140LVT U13004 ( .A1(i_data_bus[385]), .A2(n12506), .B1(
        i_data_bus[481]), .B2(n12494), .ZN(n12441) );
  ND4D1BWP30P140LVT U13005 ( .A1(n12444), .A2(n12443), .A3(n12442), .A4(n12441), .ZN(n12455) );
  AOI22D1BWP30P140LVT U13006 ( .A1(i_data_bus[97]), .A2(n12489), .B1(
        i_data_bus[993]), .B2(n12496), .ZN(n12448) );
  AOI22D1BWP30P140LVT U13007 ( .A1(i_data_bus[353]), .A2(n12491), .B1(
        i_data_bus[417]), .B2(n12481), .ZN(n12447) );
  AOI22D1BWP30P140LVT U13008 ( .A1(i_data_bus[961]), .A2(n12482), .B1(
        i_data_bus[513]), .B2(n12477), .ZN(n12446) );
  AOI22D1BWP30P140LVT U13009 ( .A1(i_data_bus[897]), .A2(n12484), .B1(
        i_data_bus[929]), .B2(n12492), .ZN(n12445) );
  ND4D1BWP30P140LVT U13010 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(n12454) );
  AOI22D1BWP30P140LVT U13011 ( .A1(i_data_bus[865]), .A2(n12513), .B1(
        i_data_bus[737]), .B2(n12518), .ZN(n12452) );
  AOI22D1BWP30P140LVT U13012 ( .A1(i_data_bus[641]), .A2(n12520), .B1(
        i_data_bus[801]), .B2(n12517), .ZN(n12451) );
  AOI22D1BWP30P140LVT U13013 ( .A1(i_data_bus[705]), .A2(n12519), .B1(
        i_data_bus[769]), .B2(n12516), .ZN(n12450) );
  AOI22D1BWP30P140LVT U13014 ( .A1(i_data_bus[673]), .A2(n12515), .B1(
        i_data_bus[833]), .B2(n12514), .ZN(n12449) );
  ND4D1BWP30P140LVT U13015 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(n12453) );
  OR4D1BWP30P140LVT U13016 ( .A1(n12456), .A2(n12455), .A3(n12454), .A4(n12453), .Z(o_data_bus[129]) );
  AOI22D1BWP30P140LVT U13017 ( .A1(i_data_bus[578]), .A2(n12480), .B1(
        i_data_bus[962]), .B2(n12482), .ZN(n12460) );
  AOI22D1BWP30P140LVT U13018 ( .A1(i_data_bus[418]), .A2(n12481), .B1(
        i_data_bus[450]), .B2(n12507), .ZN(n12459) );
  AOI22D1BWP30P140LVT U13019 ( .A1(i_data_bus[66]), .A2(n12478), .B1(
        i_data_bus[930]), .B2(n12492), .ZN(n12458) );
  AOI22D1BWP30P140LVT U13020 ( .A1(i_data_bus[994]), .A2(n12496), .B1(
        i_data_bus[258]), .B2(n12503), .ZN(n12457) );
  ND4D1BWP30P140LVT U13021 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(n12476) );
  AOI22D1BWP30P140LVT U13022 ( .A1(i_data_bus[290]), .A2(n12505), .B1(
        i_data_bus[354]), .B2(n12491), .ZN(n12464) );
  AOI22D1BWP30P140LVT U13023 ( .A1(i_data_bus[162]), .A2(n12501), .B1(
        i_data_bus[130]), .B2(n12502), .ZN(n12463) );
  AOI22D1BWP30P140LVT U13024 ( .A1(i_data_bus[194]), .A2(n12495), .B1(
        i_data_bus[482]), .B2(n12494), .ZN(n12462) );
  AOI22D1BWP30P140LVT U13025 ( .A1(i_data_bus[546]), .A2(n12479), .B1(
        i_data_bus[386]), .B2(n12506), .ZN(n12461) );
  ND4D1BWP30P140LVT U13026 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(n12475) );
  AOI22D1BWP30P140LVT U13027 ( .A1(i_data_bus[34]), .A2(n12483), .B1(
        i_data_bus[322]), .B2(n12508), .ZN(n12468) );
  AOI22D1BWP30P140LVT U13028 ( .A1(i_data_bus[2]), .A2(n12490), .B1(
        i_data_bus[514]), .B2(n12477), .ZN(n12467) );
  AOI22D1BWP30P140LVT U13029 ( .A1(i_data_bus[610]), .A2(n12504), .B1(
        i_data_bus[226]), .B2(n12493), .ZN(n12466) );
  AOI22D1BWP30P140LVT U13030 ( .A1(i_data_bus[898]), .A2(n12484), .B1(
        i_data_bus[98]), .B2(n12489), .ZN(n12465) );
  ND4D1BWP30P140LVT U13031 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n12465), .ZN(n12474) );
  AOI22D1BWP30P140LVT U13032 ( .A1(i_data_bus[674]), .A2(n12515), .B1(
        i_data_bus[834]), .B2(n12514), .ZN(n12472) );
  AOI22D1BWP30P140LVT U13033 ( .A1(i_data_bus[738]), .A2(n12518), .B1(
        i_data_bus[642]), .B2(n12520), .ZN(n12471) );
  AOI22D1BWP30P140LVT U13034 ( .A1(i_data_bus[866]), .A2(n12513), .B1(
        i_data_bus[706]), .B2(n12519), .ZN(n12470) );
  AOI22D1BWP30P140LVT U13035 ( .A1(i_data_bus[802]), .A2(n12517), .B1(
        i_data_bus[770]), .B2(n12516), .ZN(n12469) );
  ND4D1BWP30P140LVT U13036 ( .A1(n12472), .A2(n12471), .A3(n12470), .A4(n12469), .ZN(n12473) );
  OR4D1BWP30P140LVT U13037 ( .A1(n12476), .A2(n12475), .A3(n12474), .A4(n12473), .Z(o_data_bus[130]) );
  AOI22D1BWP30P140LVT U13038 ( .A1(i_data_bus[67]), .A2(n12478), .B1(
        i_data_bus[515]), .B2(n12477), .ZN(n12488) );
  AOI22D1BWP30P140LVT U13039 ( .A1(i_data_bus[579]), .A2(n12480), .B1(
        i_data_bus[547]), .B2(n12479), .ZN(n12487) );
  AOI22D1BWP30P140LVT U13040 ( .A1(i_data_bus[963]), .A2(n12482), .B1(
        i_data_bus[419]), .B2(n12481), .ZN(n12486) );
  AOI22D1BWP30P140LVT U13041 ( .A1(i_data_bus[899]), .A2(n12484), .B1(
        i_data_bus[35]), .B2(n12483), .ZN(n12485) );
  ND4D1BWP30P140LVT U13042 ( .A1(n12488), .A2(n12487), .A3(n12486), .A4(n12485), .ZN(n12528) );
  AOI22D1BWP30P140LVT U13043 ( .A1(i_data_bus[3]), .A2(n12490), .B1(
        i_data_bus[99]), .B2(n12489), .ZN(n12500) );
  AOI22D1BWP30P140LVT U13044 ( .A1(i_data_bus[931]), .A2(n12492), .B1(
        i_data_bus[355]), .B2(n12491), .ZN(n12499) );
  AOI22D1BWP30P140LVT U13045 ( .A1(i_data_bus[483]), .A2(n12494), .B1(
        i_data_bus[227]), .B2(n12493), .ZN(n12498) );
  AOI22D1BWP30P140LVT U13046 ( .A1(i_data_bus[995]), .A2(n12496), .B1(
        i_data_bus[195]), .B2(n12495), .ZN(n12497) );
  ND4D1BWP30P140LVT U13047 ( .A1(n12500), .A2(n12499), .A3(n12498), .A4(n12497), .ZN(n12527) );
  AOI22D1BWP30P140LVT U13048 ( .A1(i_data_bus[131]), .A2(n12502), .B1(
        i_data_bus[163]), .B2(n12501), .ZN(n12512) );
  AOI22D1BWP30P140LVT U13049 ( .A1(i_data_bus[611]), .A2(n12504), .B1(
        i_data_bus[259]), .B2(n12503), .ZN(n12511) );
  AOI22D1BWP30P140LVT U13050 ( .A1(i_data_bus[387]), .A2(n12506), .B1(
        i_data_bus[291]), .B2(n12505), .ZN(n12510) );
  AOI22D1BWP30P140LVT U13051 ( .A1(i_data_bus[323]), .A2(n12508), .B1(
        i_data_bus[451]), .B2(n12507), .ZN(n12509) );
  ND4D1BWP30P140LVT U13052 ( .A1(n12512), .A2(n12511), .A3(n12510), .A4(n12509), .ZN(n12526) );
  AOI22D1BWP30P140LVT U13053 ( .A1(i_data_bus[835]), .A2(n12514), .B1(
        i_data_bus[867]), .B2(n12513), .ZN(n12524) );
  AOI22D1BWP30P140LVT U13054 ( .A1(i_data_bus[771]), .A2(n12516), .B1(
        i_data_bus[675]), .B2(n12515), .ZN(n12523) );
  AOI22D1BWP30P140LVT U13055 ( .A1(i_data_bus[739]), .A2(n12518), .B1(
        i_data_bus[803]), .B2(n12517), .ZN(n12522) );
  AOI22D1BWP30P140LVT U13056 ( .A1(i_data_bus[643]), .A2(n12520), .B1(
        i_data_bus[707]), .B2(n12519), .ZN(n12521) );
  ND4D1BWP30P140LVT U13057 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12521), .ZN(n12525) );
  OR4D1BWP30P140LVT U13058 ( .A1(n12528), .A2(n12527), .A3(n12526), .A4(n12525), .Z(o_data_bus[131]) );
endmodule

