`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module controller_full(CLK, reset, from_glob_controller_delay,  input_boundary_flag, prev_dest_address, from_glob_dest_addr, packet_out, boundary_next, dest_address, from_glob_controller_valid, D, write_flag, from_glob_prefetch_valid, from_glob_prefetch_start, from_glob_prefetch_stop, from_glob_prefetch_dest, prefetch_packet_out, write_boundary_next, input_write_boundary, prefetch_next_dest_addr, prefetch_next_stop_address, prefetch_boundary_prev, input_prefetch_boundary_flag, prefetch_stop_address, prefetch_dest_addr, scenario_update);

    // parameter
    	parameter N_sample = 256;
	parameter datawidth = 16;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 4; // 16 local controllers in subscaled system
	parameter sample_address_width = 8; /// assuming 1024 rows and 64 columns: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	

//=== IO Ports ===//

     // Normal Mode Input
        input [31:0] D;



    // input
    	input CLK; // system clock, generated by VCO
	input reset;

	input from_glob_controller_valid;
	input input_boundary_flag;
	input input_prefetch_boundary_flag;
	input input_write_boundary;
	input [address_vector_width - 1:0] prev_dest_address;
	input [address_vector_width - 1:0] prefetch_next_dest_addr;
        input [address_vector_width - 1:0] prefetch_next_stop_address;
	input [address_vector_width - 1:0] from_glob_dest_addr;
	input [address_vector_width - 1:0] from_glob_prefetch_dest;
	input [sample_address_width - 1:0] from_glob_controller_delay;
	
        //input [sample_address_width-1:0] ext_sample_address_M;
	input write_flag;

	input from_glob_prefetch_valid;
	input [sample_address_width - 1:0] from_glob_prefetch_start;
	input [sample_address_width - 1:0] from_glob_prefetch_stop;
	input scenario_update;

    // output
        output [packet_width-1:0] packet_out;  
        output [packet_width-1:0] prefetch_packet_out;  
        output boundary_next;
        output write_boundary_next;
        output [address_vector_width - 1:0] dest_address;
        output prefetch_boundary_prev;
	output [address_vector_width - 1:0] prefetch_dest_addr;
    	output [sample_address_width - 1:0] prefetch_stop_address;


//////////// internal status regs/signals //////////////////////////////////
    //reg [packet_width-1:0] packet_out_internal;

    wire [2*datawidth - 1:0] data_from_sram;
    wire [2*datawidth - 1:0] sram_D;


    wire BIST;
    wire AWT;
    wire SLP;
    wire SD;
    wire CEB;
    wire WEB;
    wire CEBM;
    wire [sample_address_width-1:0] A;		
    wire [sample_address_width-1:0] AM;		
    wire sram_CEB;
    wire sram_WEB;
    wire [2*datawidth - 1:0] sram_BWEB;

    	wire [31:0] DM;
    	wire [31:0] BWEBM;
    	wire WEBM;



///////////////////////////////////////////////////////////////////////////////    

////////// logic part ///////////////////////////////////////////////////////  
    assign AM = 0;
    assign DM = 0;
    assign BWEBM = 32'hffffffff;
    assign WEBM = 1;
    assign CEBM = 1;
    assign SLP = 0;
    assign SD = 0;
    assign AWT = 0;
    assign BIST = 0;


////////////sequential logic
//
//

   only_controller_prefetch_full DUT_controller(.CLK(CLK), .reset(reset),   .from_glob_controller_delay(from_glob_controller_delay),  .input_boundary_flag(input_boundary_flag), .prev_dest_address(prev_dest_address), .from_glob_dest_addr(from_glob_dest_addr), .packet_out(packet_out), .boundary_next(boundary_next), .dest_address(dest_address), .from_glob_controller_valid(from_glob_controller_valid), .D(D), .write_flag(write_flag), .from_glob_prefetch_valid(from_glob_prefetch_valid), .from_glob_prefetch_start(from_glob_prefetch_start), .from_glob_prefetch_stop(from_glob_prefetch_stop), .from_glob_prefetch_dest(from_glob_prefetch_dest), .prefetch_packet_out(prefetch_packet_out), .write_boundary_next(write_boundary_next), .input_write_boundary(input_write_boundary), .prefetch_next_dest_addr(prefetch_next_dest_addr), .prefetch_next_stop_address(prefetch_next_stop_address), .prefetch_boundary_prev(prefetch_boundary_prev), .input_prefetch_boundary_flag(input_prefetch_boundary_flag), .prefetch_stop_address(prefetch_stop_address), .prefetch_dest_addr(prefetch_dest_addr),  .scenario_update(scenario_update), .data_from_sram(data_from_sram), .A(A), .sram_CEB(sram_CEB), .sram_WEB(sram_WEB), .sram_D(sram_D), .sram_BWEB(sram_BWEB) );

   TS1N28HPCPLVTB256X32M4SWBASO UI_dut_mem (.SLP(SLP), .SD(SD), .CLK(CLK), .CEB(sram_CEB), .WEB(sram_WEB), .CEBM(CEBM), .WEBM(WEBM), .AWT(AWT), .A(A), .D(sram_D), .BWEB(sram_BWEB), .AM(AM), .DM(DM), .BWEBM(BWEBM), .BIST(BIST), .Q(data_from_sram));



	 
	 


   
endmodule
    
