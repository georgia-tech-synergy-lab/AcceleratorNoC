
module linear_network_unicast_seq ( clk, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [31:0] i_data_bus;
  output [3:0] o_valid;
  output [127:0] o_data_bus;
  input [1:0] i_cmd;
  input clk, rst, i_valid, i_en;
  wire   N147, N148, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N284, N285, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N420, N421, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110;
  wire   [95:0] o_data_forward_reg;
  wire   [0:2] o_valid_forward_reg;
  wire   [5:0] o_cmd_forward_reg;

  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__1_ ( .D(N148), .CP(clk), .Q(
        o_cmd_forward_reg[5]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__0_ ( .D(N147), .CP(clk), .Q(
        o_cmd_forward_reg[4]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__31_ ( .D(n39), .CP(clk), .Q(
        o_data_forward_reg[95]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__30_ ( .D(n38), .CP(clk), .Q(
        o_data_forward_reg[94]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__29_ ( .D(n37), .CP(clk), .Q(
        o_data_forward_reg[93]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__28_ ( .D(n36), .CP(clk), .Q(
        o_data_forward_reg[92]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__27_ ( .D(n35), .CP(clk), .Q(
        o_data_forward_reg[91]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__26_ ( .D(n34), .CP(clk), .Q(
        o_data_forward_reg[90]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__25_ ( .D(n33), .CP(clk), .Q(
        o_data_forward_reg[89]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__24_ ( .D(n32), .CP(clk), .Q(
        o_data_forward_reg[88]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__23_ ( .D(n31), .CP(clk), .Q(
        o_data_forward_reg[87]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__22_ ( .D(n30), .CP(clk), .Q(
        o_data_forward_reg[86]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__21_ ( .D(n29), .CP(clk), .Q(
        o_data_forward_reg[85]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__20_ ( .D(n28), .CP(clk), .Q(
        o_data_forward_reg[84]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__19_ ( .D(n27), .CP(clk), .Q(
        o_data_forward_reg[83]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__18_ ( .D(n26), .CP(clk), .Q(
        o_data_forward_reg[82]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__17_ ( .D(n25), .CP(clk), .Q(
        o_data_forward_reg[81]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__16_ ( .D(n24), .CP(clk), .Q(
        o_data_forward_reg[80]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__15_ ( .D(n23), .CP(clk), .Q(
        o_data_forward_reg[79]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__14_ ( .D(n22), .CP(clk), .Q(
        o_data_forward_reg[78]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__13_ ( .D(n21), .CP(clk), .Q(
        o_data_forward_reg[77]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__12_ ( .D(n20), .CP(clk), .Q(
        o_data_forward_reg[76]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__11_ ( .D(n19), .CP(clk), .Q(
        o_data_forward_reg[75]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__10_ ( .D(n18), .CP(clk), .Q(
        o_data_forward_reg[74]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__9_ ( .D(n17), .CP(clk), .Q(
        o_data_forward_reg[73]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__8_ ( .D(n16), .CP(clk), .Q(
        o_data_forward_reg[72]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__7_ ( .D(n15), .CP(clk), .Q(
        o_data_forward_reg[71]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__6_ ( .D(n14), .CP(clk), .Q(
        o_data_forward_reg[70]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__5_ ( .D(n8), .CP(clk), .Q(
        o_data_forward_reg[69]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__4_ ( .D(n13), .CP(clk), .Q(
        o_data_forward_reg[68]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__3_ ( .D(n12), .CP(clk), .Q(
        o_data_forward_reg[67]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__2_ ( .D(n11), .CP(clk), .Q(
        o_data_forward_reg[66]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__1_ ( .D(n10), .CP(clk), .Q(
        o_data_forward_reg[65]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__0_ ( .D(n9), .CP(clk), .Q(
        o_data_forward_reg[64]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_0_ ( .D(n110), .CP(clk), .Q(
        o_valid_forward_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__1_ ( .D(N285), .CP(clk), .Q(
        o_cmd_forward_reg[3]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__0_ ( .D(N284), .CP(clk), .Q(
        o_cmd_forward_reg[2]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__31_ ( .D(N282), .CP(clk), .Q(
        o_data_forward_reg[63]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__30_ ( .D(N281), .CP(clk), .Q(
        o_data_forward_reg[62]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__29_ ( .D(N280), .CP(clk), .Q(
        o_data_forward_reg[61]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__28_ ( .D(N279), .CP(clk), .Q(
        o_data_forward_reg[60]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__27_ ( .D(N278), .CP(clk), .Q(
        o_data_forward_reg[59]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__26_ ( .D(N277), .CP(clk), .Q(
        o_data_forward_reg[58]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__25_ ( .D(N276), .CP(clk), .Q(
        o_data_forward_reg[57]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__24_ ( .D(N275), .CP(clk), .Q(
        o_data_forward_reg[56]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__23_ ( .D(N274), .CP(clk), .Q(
        o_data_forward_reg[55]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__22_ ( .D(N273), .CP(clk), .Q(
        o_data_forward_reg[54]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__21_ ( .D(N272), .CP(clk), .Q(
        o_data_forward_reg[53]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__20_ ( .D(N271), .CP(clk), .Q(
        o_data_forward_reg[52]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__19_ ( .D(N270), .CP(clk), .Q(
        o_data_forward_reg[51]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__18_ ( .D(N269), .CP(clk), .Q(
        o_data_forward_reg[50]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__17_ ( .D(N268), .CP(clk), .Q(
        o_data_forward_reg[49]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__16_ ( .D(N267), .CP(clk), .Q(
        o_data_forward_reg[48]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__15_ ( .D(N266), .CP(clk), .Q(
        o_data_forward_reg[47]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__14_ ( .D(N265), .CP(clk), .Q(
        o_data_forward_reg[46]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__13_ ( .D(N264), .CP(clk), .Q(
        o_data_forward_reg[45]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__12_ ( .D(N263), .CP(clk), .Q(
        o_data_forward_reg[44]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__11_ ( .D(N262), .CP(clk), .Q(
        o_data_forward_reg[43]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__10_ ( .D(N261), .CP(clk), .Q(
        o_data_forward_reg[42]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__9_ ( .D(N260), .CP(clk), .Q(
        o_data_forward_reg[41]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__8_ ( .D(N259), .CP(clk), .Q(
        o_data_forward_reg[40]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__7_ ( .D(N258), .CP(clk), .Q(
        o_data_forward_reg[39]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__6_ ( .D(N257), .CP(clk), .Q(
        o_data_forward_reg[38]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__5_ ( .D(N256), .CP(clk), .Q(
        o_data_forward_reg[37]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__4_ ( .D(N255), .CP(clk), .Q(
        o_data_forward_reg[36]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__3_ ( .D(N254), .CP(clk), .Q(
        o_data_forward_reg[35]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__2_ ( .D(N253), .CP(clk), .Q(
        o_data_forward_reg[34]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__1_ ( .D(N252), .CP(clk), .Q(
        o_data_forward_reg[33]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__0_ ( .D(N251), .CP(clk), .Q(
        o_data_forward_reg[32]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_1_ ( .D(n109), .CP(clk), .Q(
        o_valid_forward_reg[1]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__1_ ( .D(N421), .CP(clk), .Q(
        o_cmd_forward_reg[1]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__0_ ( .D(N420), .CP(clk), .Q(
        o_cmd_forward_reg[0]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__31_ ( .D(N418), .CP(clk), .Q(
        o_data_forward_reg[31]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__30_ ( .D(N417), .CP(clk), .Q(
        o_data_forward_reg[30]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__29_ ( .D(N416), .CP(clk), .Q(
        o_data_forward_reg[29]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__28_ ( .D(N415), .CP(clk), .Q(
        o_data_forward_reg[28]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__27_ ( .D(N414), .CP(clk), .Q(
        o_data_forward_reg[27]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__26_ ( .D(N413), .CP(clk), .Q(
        o_data_forward_reg[26]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__25_ ( .D(N412), .CP(clk), .Q(
        o_data_forward_reg[25]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__24_ ( .D(N411), .CP(clk), .Q(
        o_data_forward_reg[24]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__23_ ( .D(N410), .CP(clk), .Q(
        o_data_forward_reg[23]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__22_ ( .D(N409), .CP(clk), .Q(
        o_data_forward_reg[22]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__21_ ( .D(N408), .CP(clk), .Q(
        o_data_forward_reg[21]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__20_ ( .D(N407), .CP(clk), .Q(
        o_data_forward_reg[20]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__19_ ( .D(N406), .CP(clk), .Q(
        o_data_forward_reg[19]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__18_ ( .D(N405), .CP(clk), .Q(
        o_data_forward_reg[18]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__17_ ( .D(N404), .CP(clk), .Q(
        o_data_forward_reg[17]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__16_ ( .D(N403), .CP(clk), .Q(
        o_data_forward_reg[16]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__15_ ( .D(N402), .CP(clk), .Q(
        o_data_forward_reg[15]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__14_ ( .D(N401), .CP(clk), .Q(
        o_data_forward_reg[14]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__13_ ( .D(N400), .CP(clk), .Q(
        o_data_forward_reg[13]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__12_ ( .D(N399), .CP(clk), .Q(
        o_data_forward_reg[12]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__11_ ( .D(N398), .CP(clk), .Q(
        o_data_forward_reg[11]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__10_ ( .D(N397), .CP(clk), .Q(
        o_data_forward_reg[10]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__9_ ( .D(N396), .CP(clk), .Q(
        o_data_forward_reg[9]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__8_ ( .D(N395), .CP(clk), .Q(
        o_data_forward_reg[8]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__7_ ( .D(N394), .CP(clk), .Q(
        o_data_forward_reg[7]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__6_ ( .D(N393), .CP(clk), .Q(
        o_data_forward_reg[6]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__5_ ( .D(N392), .CP(clk), .Q(
        o_data_forward_reg[5]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__4_ ( .D(N391), .CP(clk), .Q(
        o_data_forward_reg[4]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__3_ ( .D(N390), .CP(clk), .Q(
        o_data_forward_reg[3]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__2_ ( .D(N389), .CP(clk), .Q(
        o_data_forward_reg[2]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__1_ ( .D(N388), .CP(clk), .Q(
        o_data_forward_reg[1]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__0_ ( .D(N387), .CP(clk), .Q(
        o_data_forward_reg[0]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_2_ ( .D(n107), .CP(clk), .Q(
        o_valid_forward_reg[2]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_3_ ( .D(n105), .CP(clk), .Q(o_valid[3]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_2_ ( .D(n106), .CP(clk), .Q(o_valid[2]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_1_ ( .D(n108), .CP(clk), .Q(o_valid[1]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_0_ ( .D(n104), .CP(clk), .Q(o_valid[0]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(n97), .CP(clk), .Q(
        o_data_bus[127]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(n96), .CP(clk), .Q(
        o_data_bus[126]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(n95), .CP(clk), .Q(
        o_data_bus[125]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(n94), .CP(clk), .Q(
        o_data_bus[124]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(n93), .CP(clk), .Q(
        o_data_bus[123]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(n92), .CP(clk), .Q(
        o_data_bus[122]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(n65), .CP(clk), .Q(
        o_data_bus[121]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(n64), .CP(clk), .Q(
        o_data_bus[120]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(n63), .CP(clk), .Q(
        o_data_bus[119]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(n62), .CP(clk), .Q(
        o_data_bus[118]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(n61), .CP(clk), .Q(
        o_data_bus[117]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(n60), .CP(clk), .Q(
        o_data_bus[116]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(n59), .CP(clk), .Q(
        o_data_bus[115]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(n58), .CP(clk), .Q(
        o_data_bus[114]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(n57), .CP(clk), .Q(
        o_data_bus[113]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(n56), .CP(clk), .Q(
        o_data_bus[112]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(n55), .CP(clk), .Q(
        o_data_bus[111]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(n54), .CP(clk), .Q(
        o_data_bus[110]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(n53), .CP(clk), .Q(
        o_data_bus[109]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(n52), .CP(clk), .Q(
        o_data_bus[108]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(n51), .CP(clk), .Q(
        o_data_bus[107]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(n50), .CP(clk), .Q(
        o_data_bus[106]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(n49), .CP(clk), .Q(
        o_data_bus[105]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(n48), .CP(clk), .Q(
        o_data_bus[104]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(n47), .CP(clk), .Q(
        o_data_bus[103]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(n46), .CP(clk), .Q(
        o_data_bus[102]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(n45), .CP(clk), .Q(
        o_data_bus[101]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(n44), .CP(clk), .Q(
        o_data_bus[100]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(n43), .CP(clk), .Q(
        o_data_bus[99]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(n42), .CP(clk), .Q(
        o_data_bus[98]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(n41), .CP(clk), .Q(
        o_data_bus[97]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(n40), .CP(clk), .Q(
        o_data_bus[96]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(N386), .CP(clk), .Q(
        o_data_bus[95]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(N385), .CP(clk), .Q(
        o_data_bus[94]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(N384), .CP(clk), .Q(
        o_data_bus[93]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(N383), .CP(clk), .Q(
        o_data_bus[92]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(N382), .CP(clk), .Q(
        o_data_bus[91]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(N381), .CP(clk), .Q(
        o_data_bus[90]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(N380), .CP(clk), .Q(
        o_data_bus[89]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(N379), .CP(clk), .Q(
        o_data_bus[88]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(N378), .CP(clk), .Q(
        o_data_bus[87]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(N377), .CP(clk), .Q(
        o_data_bus[86]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(N376), .CP(clk), .Q(
        o_data_bus[85]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(N375), .CP(clk), .Q(
        o_data_bus[84]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(N374), .CP(clk), .Q(
        o_data_bus[83]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(N373), .CP(clk), .Q(
        o_data_bus[82]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(N372), .CP(clk), .Q(
        o_data_bus[81]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(N371), .CP(clk), .Q(
        o_data_bus[80]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(N370), .CP(clk), .Q(
        o_data_bus[79]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(N369), .CP(clk), .Q(
        o_data_bus[78]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(N368), .CP(clk), .Q(
        o_data_bus[77]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(N367), .CP(clk), .Q(
        o_data_bus[76]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(N366), .CP(clk), .Q(
        o_data_bus[75]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N365), .CP(clk), .Q(
        o_data_bus[74]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N364), .CP(clk), .Q(
        o_data_bus[73]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N363), .CP(clk), .Q(
        o_data_bus[72]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N362), .CP(clk), .Q(
        o_data_bus[71]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N361), .CP(clk), .Q(
        o_data_bus[70]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N360), .CP(clk), .Q(
        o_data_bus[69]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N359), .CP(clk), .Q(
        o_data_bus[68]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N358), .CP(clk), .Q(
        o_data_bus[67]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N357), .CP(clk), .Q(
        o_data_bus[66]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N356), .CP(clk), .Q(
        o_data_bus[65]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N355), .CP(clk), .Q(
        o_data_bus[64]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N250), .CP(clk), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N249), .CP(clk), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N248), .CP(clk), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N247), .CP(clk), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N246), .CP(clk), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N245), .CP(clk), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N244), .CP(clk), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N243), .CP(clk), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N242), .CP(clk), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N241), .CP(clk), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N240), .CP(clk), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N239), .CP(clk), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N238), .CP(clk), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N237), .CP(clk), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N236), .CP(clk), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N235), .CP(clk), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N234), .CP(clk), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N233), .CP(clk), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N232), .CP(clk), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N231), .CP(clk), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N230), .CP(clk), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N229), .CP(clk), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N228), .CP(clk), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N227), .CP(clk), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N226), .CP(clk), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N225), .CP(clk), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N224), .CP(clk), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N223), .CP(clk), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N222), .CP(clk), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N221), .CP(clk), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N220), .CP(clk), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N219), .CP(clk), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(n103), .CP(clk), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(n102), .CP(clk), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(n101), .CP(clk), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(n100), .CP(clk), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(n99), .CP(clk), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(n98), .CP(clk), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(n91), .CP(clk), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(n90), .CP(clk), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(n89), .CP(clk), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(n88), .CP(clk), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(n87), .CP(clk), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(n86), .CP(clk), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(n85), .CP(clk), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(n84), .CP(clk), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(n83), .CP(clk), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(n82), .CP(clk), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(n81), .CP(clk), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(n80), .CP(clk), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(n79), .CP(clk), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(n78), .CP(clk), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(n77), .CP(clk), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(n76), .CP(clk), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(n75), .CP(clk), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(n74), .CP(clk), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(n73), .CP(clk), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(n72), .CP(clk), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(n71), .CP(clk), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(n70), .CP(clk), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(n69), .CP(clk), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(n68), .CP(clk), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(n67), .CP(clk), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(n66), .CP(clk), .Q(
        o_data_bus[0]) );
  INR2D4BWP30P140LVT U242 ( .A1(n110), .B1(n5), .ZN(n104) );
  NR2D1BWP30P140LVT U243 ( .A1(o_cmd_forward_reg[1]), .A2(o_cmd_forward_reg[0]), .ZN(n4) );
  OR2D1BWP30P140LVT U244 ( .A1(i_cmd[1]), .A2(i_cmd[0]), .Z(n5) );
  CKAN2D1BWP30P140LVT U245 ( .A1(n109), .A2(n4), .Z(n108) );
  CKAN2D1BWP30P140LVT U246 ( .A1(n107), .A2(n4), .Z(n106) );
  ND2D1BWP30P140LVT U247 ( .A1(o_valid_forward_reg[2]), .A2(n7), .ZN(n3) );
  INR2D1BWP30P140LVT U248 ( .A1(o_valid_forward_reg[1]), .B1(n6), .ZN(n107) );
  INR2D1BWP30P140LVT U249 ( .A1(o_valid_forward_reg[0]), .B1(n6), .ZN(n109) );
  INR2D1BWP30P140LVT U250 ( .A1(i_valid), .B1(n6), .ZN(n110) );
  INVD1BWP30P140LVT U251 ( .I(n7), .ZN(n6) );
  INR2D1BWP30P140LVT U252 ( .A1(i_en), .B1(rst), .ZN(n7) );
  CKAN2D1BWP30P140LVT U253 ( .A1(n108), .A2(o_data_forward_reg[64]), .Z(N219)
         );
  CKAN2D1BWP30P140LVT U254 ( .A1(n108), .A2(o_data_forward_reg[65]), .Z(N220)
         );
  CKAN2D1BWP30P140LVT U255 ( .A1(n108), .A2(o_data_forward_reg[66]), .Z(N221)
         );
  CKAN2D1BWP30P140LVT U256 ( .A1(n108), .A2(o_data_forward_reg[67]), .Z(N222)
         );
  CKAN2D1BWP30P140LVT U257 ( .A1(n108), .A2(o_data_forward_reg[68]), .Z(N223)
         );
  CKAN2D1BWP30P140LVT U258 ( .A1(n108), .A2(o_data_forward_reg[69]), .Z(N224)
         );
  CKAN2D1BWP30P140LVT U259 ( .A1(n108), .A2(o_data_forward_reg[70]), .Z(N225)
         );
  CKAN2D1BWP30P140LVT U260 ( .A1(n108), .A2(o_data_forward_reg[71]), .Z(N226)
         );
  CKAN2D1BWP30P140LVT U261 ( .A1(n108), .A2(o_data_forward_reg[72]), .Z(N227)
         );
  CKAN2D1BWP30P140LVT U262 ( .A1(n108), .A2(o_data_forward_reg[73]), .Z(N228)
         );
  CKAN2D1BWP30P140LVT U263 ( .A1(n108), .A2(o_data_forward_reg[74]), .Z(N229)
         );
  CKAN2D1BWP30P140LVT U264 ( .A1(n108), .A2(o_data_forward_reg[75]), .Z(N230)
         );
  CKAN2D1BWP30P140LVT U265 ( .A1(n108), .A2(o_data_forward_reg[76]), .Z(N231)
         );
  CKAN2D1BWP30P140LVT U266 ( .A1(n108), .A2(o_data_forward_reg[77]), .Z(N232)
         );
  CKAN2D1BWP30P140LVT U267 ( .A1(n108), .A2(o_data_forward_reg[78]), .Z(N233)
         );
  CKAN2D1BWP30P140LVT U268 ( .A1(n108), .A2(o_data_forward_reg[79]), .Z(N234)
         );
  CKAN2D1BWP30P140LVT U269 ( .A1(n108), .A2(o_data_forward_reg[80]), .Z(N235)
         );
  CKAN2D1BWP30P140LVT U270 ( .A1(n108), .A2(o_data_forward_reg[81]), .Z(N236)
         );
  CKAN2D1BWP30P140LVT U271 ( .A1(n108), .A2(o_data_forward_reg[82]), .Z(N237)
         );
  CKAN2D1BWP30P140LVT U272 ( .A1(n108), .A2(o_data_forward_reg[83]), .Z(N238)
         );
  CKAN2D1BWP30P140LVT U273 ( .A1(n108), .A2(o_data_forward_reg[84]), .Z(N239)
         );
  CKAN2D1BWP30P140LVT U274 ( .A1(n108), .A2(o_data_forward_reg[85]), .Z(N240)
         );
  CKAN2D1BWP30P140LVT U275 ( .A1(n108), .A2(o_data_forward_reg[86]), .Z(N241)
         );
  CKAN2D1BWP30P140LVT U276 ( .A1(n108), .A2(o_data_forward_reg[87]), .Z(N242)
         );
  CKAN2D1BWP30P140LVT U277 ( .A1(n108), .A2(o_data_forward_reg[88]), .Z(N243)
         );
  CKAN2D1BWP30P140LVT U278 ( .A1(n108), .A2(o_data_forward_reg[89]), .Z(N244)
         );
  CKAN2D1BWP30P140LVT U279 ( .A1(n108), .A2(o_data_forward_reg[90]), .Z(N245)
         );
  CKAN2D1BWP30P140LVT U280 ( .A1(n108), .A2(o_data_forward_reg[91]), .Z(N246)
         );
  CKAN2D1BWP30P140LVT U281 ( .A1(n108), .A2(o_data_forward_reg[92]), .Z(N247)
         );
  CKAN2D1BWP30P140LVT U282 ( .A1(n108), .A2(o_data_forward_reg[93]), .Z(N248)
         );
  CKAN2D1BWP30P140LVT U283 ( .A1(n108), .A2(o_data_forward_reg[94]), .Z(N249)
         );
  CKAN2D1BWP30P140LVT U284 ( .A1(n108), .A2(o_data_forward_reg[95]), .Z(N250)
         );
  CKAN2D1BWP30P140LVT U285 ( .A1(n106), .A2(o_data_forward_reg[32]), .Z(N355)
         );
  CKAN2D1BWP30P140LVT U286 ( .A1(n106), .A2(o_data_forward_reg[33]), .Z(N356)
         );
  CKAN2D1BWP30P140LVT U287 ( .A1(n106), .A2(o_data_forward_reg[34]), .Z(N357)
         );
  CKAN2D1BWP30P140LVT U288 ( .A1(n106), .A2(o_data_forward_reg[35]), .Z(N358)
         );
  CKAN2D1BWP30P140LVT U289 ( .A1(n106), .A2(o_data_forward_reg[36]), .Z(N359)
         );
  CKAN2D1BWP30P140LVT U290 ( .A1(n106), .A2(o_data_forward_reg[37]), .Z(N360)
         );
  CKAN2D1BWP30P140LVT U291 ( .A1(n106), .A2(o_data_forward_reg[38]), .Z(N361)
         );
  CKAN2D1BWP30P140LVT U292 ( .A1(n106), .A2(o_data_forward_reg[39]), .Z(N362)
         );
  CKAN2D1BWP30P140LVT U293 ( .A1(n106), .A2(o_data_forward_reg[40]), .Z(N363)
         );
  CKAN2D1BWP30P140LVT U294 ( .A1(n106), .A2(o_data_forward_reg[41]), .Z(N364)
         );
  CKAN2D1BWP30P140LVT U295 ( .A1(n106), .A2(o_data_forward_reg[42]), .Z(N365)
         );
  CKAN2D1BWP30P140LVT U296 ( .A1(n106), .A2(o_data_forward_reg[43]), .Z(N366)
         );
  CKAN2D1BWP30P140LVT U297 ( .A1(n106), .A2(o_data_forward_reg[44]), .Z(N367)
         );
  CKAN2D1BWP30P140LVT U298 ( .A1(n106), .A2(o_data_forward_reg[45]), .Z(N368)
         );
  CKAN2D1BWP30P140LVT U299 ( .A1(n106), .A2(o_data_forward_reg[46]), .Z(N369)
         );
  CKAN2D1BWP30P140LVT U300 ( .A1(n106), .A2(o_data_forward_reg[47]), .Z(N370)
         );
  CKAN2D1BWP30P140LVT U301 ( .A1(n106), .A2(o_data_forward_reg[48]), .Z(N371)
         );
  CKAN2D1BWP30P140LVT U302 ( .A1(n106), .A2(o_data_forward_reg[49]), .Z(N372)
         );
  CKAN2D1BWP30P140LVT U303 ( .A1(n106), .A2(o_data_forward_reg[50]), .Z(N373)
         );
  CKAN2D1BWP30P140LVT U304 ( .A1(n106), .A2(o_data_forward_reg[51]), .Z(N374)
         );
  CKAN2D1BWP30P140LVT U305 ( .A1(n106), .A2(o_data_forward_reg[52]), .Z(N375)
         );
  CKAN2D1BWP30P140LVT U306 ( .A1(n106), .A2(o_data_forward_reg[53]), .Z(N376)
         );
  CKAN2D1BWP30P140LVT U307 ( .A1(n106), .A2(o_data_forward_reg[54]), .Z(N377)
         );
  CKAN2D1BWP30P140LVT U308 ( .A1(n106), .A2(o_data_forward_reg[55]), .Z(N378)
         );
  CKAN2D1BWP30P140LVT U309 ( .A1(n106), .A2(o_data_forward_reg[56]), .Z(N379)
         );
  CKAN2D1BWP30P140LVT U310 ( .A1(n106), .A2(o_data_forward_reg[57]), .Z(N380)
         );
  CKAN2D1BWP30P140LVT U311 ( .A1(n106), .A2(o_data_forward_reg[58]), .Z(N381)
         );
  CKAN2D1BWP30P140LVT U312 ( .A1(n106), .A2(o_data_forward_reg[59]), .Z(N382)
         );
  CKAN2D1BWP30P140LVT U313 ( .A1(n106), .A2(o_data_forward_reg[60]), .Z(N383)
         );
  CKAN2D1BWP30P140LVT U314 ( .A1(n106), .A2(o_data_forward_reg[61]), .Z(N384)
         );
  CKAN2D1BWP30P140LVT U315 ( .A1(n106), .A2(o_data_forward_reg[62]), .Z(N385)
         );
  CKAN2D1BWP30P140LVT U316 ( .A1(n106), .A2(o_data_forward_reg[63]), .Z(N386)
         );
  CKAN2D1BWP30P140LVT U317 ( .A1(n7), .A2(o_cmd_forward_reg[4]), .Z(N284) );
  CKAN2D1BWP30P140LVT U318 ( .A1(n7), .A2(o_cmd_forward_reg[5]), .Z(N285) );
  CKAN2D1BWP30P140LVT U319 ( .A1(i_data_bus[4]), .A2(n7), .Z(n13) );
  CKAN2D1BWP30P140LVT U320 ( .A1(i_data_bus[11]), .A2(n7), .Z(n19) );
  CKAN2D1BWP30P140LVT U321 ( .A1(i_data_bus[14]), .A2(n7), .Z(n22) );
  CKAN2D1BWP30P140LVT U322 ( .A1(i_data_bus[7]), .A2(n7), .Z(n15) );
  CKAN2D1BWP30P140LVT U323 ( .A1(i_data_bus[22]), .A2(n7), .Z(n30) );
  CKAN2D1BWP30P140LVT U324 ( .A1(i_data_bus[3]), .A2(n7), .Z(n12) );
  CKAN2D1BWP30P140LVT U325 ( .A1(i_data_bus[18]), .A2(n7), .Z(n26) );
  CKAN2D1BWP30P140LVT U326 ( .A1(i_data_bus[21]), .A2(n7), .Z(n29) );
  CKAN2D1BWP30P140LVT U327 ( .A1(i_data_bus[25]), .A2(n7), .Z(n33) );
  CKAN2D1BWP30P140LVT U328 ( .A1(i_data_bus[9]), .A2(n7), .Z(n17) );
  CKAN2D1BWP30P140LVT U329 ( .A1(i_data_bus[16]), .A2(n7), .Z(n24) );
  CKAN2D1BWP30P140LVT U330 ( .A1(i_data_bus[2]), .A2(n7), .Z(n11) );
  INR2D2BWP30P140LVT U331 ( .A1(n4), .B1(n3), .ZN(n105) );
  CKAN2D1BWP30P140LVT U332 ( .A1(i_data_bus[0]), .A2(n7), .Z(n9) );
  CKAN2D1BWP30P140LVT U333 ( .A1(i_data_bus[28]), .A2(n7), .Z(n36) );
  CKAN2D1BWP30P140LVT U334 ( .A1(i_data_bus[29]), .A2(n7), .Z(n37) );
  CKAN2D1BWP30P140LVT U335 ( .A1(i_data_bus[1]), .A2(n7), .Z(n10) );
  CKAN2D1BWP30P140LVT U336 ( .A1(i_data_bus[31]), .A2(n7), .Z(n39) );
  CKAN2D1BWP30P140LVT U337 ( .A1(i_data_bus[17]), .A2(n7), .Z(n25) );
  CKAN2D1BWP30P140LVT U338 ( .A1(i_data_bus[10]), .A2(n7), .Z(n18) );
  CKAN2D1BWP30P140LVT U339 ( .A1(i_data_bus[5]), .A2(n7), .Z(n8) );
  CKAN2D1BWP30P140LVT U340 ( .A1(i_data_bus[6]), .A2(n7), .Z(n14) );
  CKAN2D1BWP30P140LVT U341 ( .A1(i_data_bus[13]), .A2(n7), .Z(n21) );
  CKAN2D1BWP30P140LVT U342 ( .A1(i_data_bus[8]), .A2(n7), .Z(n16) );
  CKAN2D1BWP30P140LVT U343 ( .A1(i_data_bus[23]), .A2(n7), .Z(n31) );
  CKAN2D1BWP30P140LVT U344 ( .A1(i_data_bus[27]), .A2(n7), .Z(n35) );
  CKAN2D1BWP30P140LVT U345 ( .A1(i_data_bus[26]), .A2(n7), .Z(n34) );
  CKAN2D1BWP30P140LVT U346 ( .A1(i_data_bus[12]), .A2(n7), .Z(n20) );
  CKAN2D1BWP30P140LVT U347 ( .A1(i_data_bus[19]), .A2(n7), .Z(n27) );
  CKAN2D1BWP30P140LVT U348 ( .A1(i_data_bus[20]), .A2(n7), .Z(n28) );
  CKAN2D1BWP30P140LVT U349 ( .A1(i_data_bus[15]), .A2(n7), .Z(n23) );
  CKAN2D1BWP30P140LVT U350 ( .A1(i_data_bus[24]), .A2(n7), .Z(n32) );
  CKAN2D1BWP30P140LVT U351 ( .A1(i_data_bus[30]), .A2(n7), .Z(n38) );
  INR2D1BWP30P140LVT U352 ( .A1(o_data_forward_reg[62]), .B1(n6), .ZN(N417) );
  INR2D1BWP30P140LVT U353 ( .A1(o_data_forward_reg[63]), .B1(n6), .ZN(N418) );
  INR2D1BWP30P140LVT U354 ( .A1(o_data_forward_reg[33]), .B1(n6), .ZN(N388) );
  INR2D1BWP30P140LVT U355 ( .A1(o_data_forward_reg[32]), .B1(n6), .ZN(N387) );
  INR2D1BWP30P140LVT U356 ( .A1(o_data_forward_reg[94]), .B1(n6), .ZN(N281) );
  INR2D1BWP30P140LVT U357 ( .A1(o_data_forward_reg[95]), .B1(n6), .ZN(N282) );
  INR2D1BWP30P140LVT U358 ( .A1(o_data_forward_reg[92]), .B1(n6), .ZN(N279) );
  INR2D1BWP30P140LVT U359 ( .A1(o_data_forward_reg[93]), .B1(n6), .ZN(N280) );
  INR2D1BWP30P140LVT U360 ( .A1(o_data_forward_reg[90]), .B1(n6), .ZN(N277) );
  INR2D1BWP30P140LVT U361 ( .A1(o_data_forward_reg[91]), .B1(n6), .ZN(N278) );
  INR2D1BWP30P140LVT U362 ( .A1(o_data_forward_reg[87]), .B1(n6), .ZN(N274) );
  INR2D1BWP30P140LVT U363 ( .A1(o_data_forward_reg[88]), .B1(n6), .ZN(N275) );
  INR2D1BWP30P140LVT U364 ( .A1(o_data_forward_reg[89]), .B1(n6), .ZN(N276) );
  INR2D1BWP30P140LVT U365 ( .A1(o_data_forward_reg[35]), .B1(n6), .ZN(N390) );
  INR2D1BWP30P140LVT U366 ( .A1(o_data_forward_reg[34]), .B1(n6), .ZN(N389) );
  INR2D1BWP30P140LVT U367 ( .A1(o_data_forward_reg[44]), .B1(n6), .ZN(N399) );
  INR2D1BWP30P140LVT U368 ( .A1(o_data_forward_reg[40]), .B1(n6), .ZN(N395) );
  INR2D1BWP30P140LVT U369 ( .A1(o_data_forward_reg[41]), .B1(n6), .ZN(N396) );
  INR2D1BWP30P140LVT U370 ( .A1(o_data_forward_reg[45]), .B1(n6), .ZN(N400) );
  INR2D1BWP30P140LVT U371 ( .A1(o_data_forward_reg[43]), .B1(n6), .ZN(N398) );
  INR2D1BWP30P140LVT U372 ( .A1(o_data_forward_reg[57]), .B1(n6), .ZN(N412) );
  INR2D1BWP30P140LVT U373 ( .A1(o_data_forward_reg[58]), .B1(n6), .ZN(N413) );
  INR2D1BWP30P140LVT U374 ( .A1(o_data_forward_reg[46]), .B1(n6), .ZN(N401) );
  INR2D1BWP30P140LVT U375 ( .A1(o_data_forward_reg[47]), .B1(n6), .ZN(N402) );
  INR2D1BWP30P140LVT U376 ( .A1(o_data_forward_reg[48]), .B1(n6), .ZN(N403) );
  INR2D1BWP30P140LVT U377 ( .A1(o_data_forward_reg[49]), .B1(n6), .ZN(N404) );
  INR2D1BWP30P140LVT U378 ( .A1(o_data_forward_reg[50]), .B1(n6), .ZN(N405) );
  INR2D1BWP30P140LVT U379 ( .A1(o_data_forward_reg[51]), .B1(n6), .ZN(N406) );
  INR2D1BWP30P140LVT U380 ( .A1(o_data_forward_reg[52]), .B1(n6), .ZN(N407) );
  INR2D1BWP30P140LVT U381 ( .A1(o_data_forward_reg[53]), .B1(n6), .ZN(N408) );
  INR2D1BWP30P140LVT U382 ( .A1(o_data_forward_reg[54]), .B1(n6), .ZN(N409) );
  INR2D1BWP30P140LVT U383 ( .A1(o_data_forward_reg[42]), .B1(n6), .ZN(N397) );
  INR2D1BWP30P140LVT U384 ( .A1(o_data_forward_reg[56]), .B1(n6), .ZN(N411) );
  INR2D1BWP30P140LVT U385 ( .A1(o_data_forward_reg[68]), .B1(n6), .ZN(N255) );
  INR2D1BWP30P140LVT U386 ( .A1(o_data_forward_reg[69]), .B1(n6), .ZN(N256) );
  INR2D1BWP30P140LVT U387 ( .A1(o_data_forward_reg[70]), .B1(n6), .ZN(N257) );
  INR2D1BWP30P140LVT U388 ( .A1(o_data_forward_reg[71]), .B1(n6), .ZN(N258) );
  INR2D1BWP30P140LVT U389 ( .A1(o_data_forward_reg[72]), .B1(n6), .ZN(N259) );
  INR2D1BWP30P140LVT U390 ( .A1(o_data_forward_reg[73]), .B1(n6), .ZN(N260) );
  INR2D1BWP30P140LVT U391 ( .A1(o_data_forward_reg[74]), .B1(n6), .ZN(N261) );
  INR2D1BWP30P140LVT U392 ( .A1(o_data_forward_reg[75]), .B1(n6), .ZN(N262) );
  INR2D1BWP30P140LVT U393 ( .A1(o_data_forward_reg[76]), .B1(n6), .ZN(N263) );
  INR2D1BWP30P140LVT U394 ( .A1(o_data_forward_reg[38]), .B1(n6), .ZN(N393) );
  INR2D1BWP30P140LVT U395 ( .A1(o_data_forward_reg[78]), .B1(n6), .ZN(N265) );
  INR2D1BWP30P140LVT U396 ( .A1(o_data_forward_reg[55]), .B1(n6), .ZN(N410) );
  INR2D1BWP30P140LVT U397 ( .A1(o_data_forward_reg[39]), .B1(n6), .ZN(N394) );
  INR2D1BWP30P140LVT U398 ( .A1(o_data_forward_reg[81]), .B1(n6), .ZN(N268) );
  INR2D1BWP30P140LVT U399 ( .A1(o_data_forward_reg[82]), .B1(n6), .ZN(N269) );
  INR2D1BWP30P140LVT U400 ( .A1(o_data_forward_reg[83]), .B1(n6), .ZN(N270) );
  INR2D1BWP30P140LVT U401 ( .A1(o_data_forward_reg[84]), .B1(n6), .ZN(N271) );
  INR2D1BWP30P140LVT U402 ( .A1(o_data_forward_reg[85]), .B1(n6), .ZN(N272) );
  INR2D1BWP30P140LVT U403 ( .A1(o_data_forward_reg[86]), .B1(n6), .ZN(N273) );
  INR2D1BWP30P140LVT U404 ( .A1(o_data_forward_reg[59]), .B1(n6), .ZN(N414) );
  INR2D1BWP30P140LVT U405 ( .A1(o_data_forward_reg[60]), .B1(n6), .ZN(N415) );
  INR2D1BWP30P140LVT U406 ( .A1(o_data_forward_reg[61]), .B1(n6), .ZN(N416) );
  INR2D1BWP30P140LVT U407 ( .A1(o_data_forward_reg[37]), .B1(n6), .ZN(N392) );
  INR2D1BWP30P140LVT U408 ( .A1(o_data_forward_reg[36]), .B1(n6), .ZN(N391) );
  INR2D1BWP30P140LVT U409 ( .A1(o_data_forward_reg[79]), .B1(n6), .ZN(N266) );
  INR2D1BWP30P140LVT U410 ( .A1(o_data_forward_reg[80]), .B1(n6), .ZN(N267) );
  INR2D1BWP30P140LVT U411 ( .A1(o_data_forward_reg[64]), .B1(n6), .ZN(N251) );
  INR2D1BWP30P140LVT U412 ( .A1(o_data_forward_reg[65]), .B1(n6), .ZN(N252) );
  INR2D1BWP30P140LVT U413 ( .A1(o_data_forward_reg[66]), .B1(n6), .ZN(N253) );
  INR2D1BWP30P140LVT U414 ( .A1(o_data_forward_reg[67]), .B1(n6), .ZN(N254) );
  INR2D1BWP30P140LVT U415 ( .A1(o_data_forward_reg[77]), .B1(n6), .ZN(N264) );
  CKAN2D1BWP30P140LVT U416 ( .A1(n105), .A2(o_data_forward_reg[0]), .Z(n40) );
  CKAN2D1BWP30P140LVT U417 ( .A1(n105), .A2(o_data_forward_reg[1]), .Z(n41) );
  CKAN2D1BWP30P140LVT U418 ( .A1(n105), .A2(o_data_forward_reg[2]), .Z(n42) );
  CKAN2D1BWP30P140LVT U419 ( .A1(n105), .A2(o_data_forward_reg[3]), .Z(n43) );
  CKAN2D1BWP30P140LVT U420 ( .A1(n105), .A2(o_data_forward_reg[4]), .Z(n44) );
  CKAN2D1BWP30P140LVT U421 ( .A1(n105), .A2(o_data_forward_reg[5]), .Z(n45) );
  CKAN2D1BWP30P140LVT U422 ( .A1(n105), .A2(o_data_forward_reg[6]), .Z(n46) );
  CKAN2D1BWP30P140LVT U423 ( .A1(n105), .A2(o_data_forward_reg[7]), .Z(n47) );
  CKAN2D1BWP30P140LVT U424 ( .A1(n105), .A2(o_data_forward_reg[8]), .Z(n48) );
  CKAN2D1BWP30P140LVT U425 ( .A1(n105), .A2(o_data_forward_reg[9]), .Z(n49) );
  CKAN2D1BWP30P140LVT U426 ( .A1(n105), .A2(o_data_forward_reg[10]), .Z(n50)
         );
  CKAN2D1BWP30P140LVT U427 ( .A1(n105), .A2(o_data_forward_reg[11]), .Z(n51)
         );
  CKAN2D1BWP30P140LVT U428 ( .A1(n105), .A2(o_data_forward_reg[12]), .Z(n52)
         );
  CKAN2D1BWP30P140LVT U429 ( .A1(n105), .A2(o_data_forward_reg[13]), .Z(n53)
         );
  CKAN2D1BWP30P140LVT U430 ( .A1(n105), .A2(o_data_forward_reg[14]), .Z(n54)
         );
  CKAN2D1BWP30P140LVT U431 ( .A1(n105), .A2(o_data_forward_reg[15]), .Z(n55)
         );
  CKAN2D1BWP30P140LVT U432 ( .A1(n105), .A2(o_data_forward_reg[16]), .Z(n56)
         );
  CKAN2D1BWP30P140LVT U433 ( .A1(n105), .A2(o_data_forward_reg[17]), .Z(n57)
         );
  CKAN2D1BWP30P140LVT U434 ( .A1(n105), .A2(o_data_forward_reg[18]), .Z(n58)
         );
  CKAN2D1BWP30P140LVT U435 ( .A1(n105), .A2(o_data_forward_reg[19]), .Z(n59)
         );
  CKAN2D1BWP30P140LVT U436 ( .A1(n105), .A2(o_data_forward_reg[20]), .Z(n60)
         );
  CKAN2D1BWP30P140LVT U437 ( .A1(n105), .A2(o_data_forward_reg[21]), .Z(n61)
         );
  CKAN2D1BWP30P140LVT U438 ( .A1(n105), .A2(o_data_forward_reg[22]), .Z(n62)
         );
  CKAN2D1BWP30P140LVT U439 ( .A1(n105), .A2(o_data_forward_reg[23]), .Z(n63)
         );
  CKAN2D1BWP30P140LVT U440 ( .A1(n105), .A2(o_data_forward_reg[24]), .Z(n64)
         );
  CKAN2D1BWP30P140LVT U441 ( .A1(n105), .A2(o_data_forward_reg[25]), .Z(n65)
         );
  CKAN2D1BWP30P140LVT U442 ( .A1(n104), .A2(i_data_bus[0]), .Z(n66) );
  CKAN2D1BWP30P140LVT U443 ( .A1(n104), .A2(i_data_bus[1]), .Z(n67) );
  CKAN2D1BWP30P140LVT U444 ( .A1(n104), .A2(i_data_bus[2]), .Z(n68) );
  CKAN2D1BWP30P140LVT U445 ( .A1(n104), .A2(i_data_bus[3]), .Z(n69) );
  CKAN2D1BWP30P140LVT U446 ( .A1(n104), .A2(i_data_bus[4]), .Z(n70) );
  CKAN2D1BWP30P140LVT U447 ( .A1(n104), .A2(i_data_bus[5]), .Z(n71) );
  CKAN2D1BWP30P140LVT U448 ( .A1(n104), .A2(i_data_bus[6]), .Z(n72) );
  CKAN2D1BWP30P140LVT U449 ( .A1(n104), .A2(i_data_bus[7]), .Z(n73) );
  CKAN2D1BWP30P140LVT U450 ( .A1(n104), .A2(i_data_bus[8]), .Z(n74) );
  CKAN2D1BWP30P140LVT U451 ( .A1(n104), .A2(i_data_bus[9]), .Z(n75) );
  CKAN2D1BWP30P140LVT U452 ( .A1(n104), .A2(i_data_bus[10]), .Z(n76) );
  CKAN2D1BWP30P140LVT U453 ( .A1(n104), .A2(i_data_bus[11]), .Z(n77) );
  CKAN2D1BWP30P140LVT U454 ( .A1(n104), .A2(i_data_bus[12]), .Z(n78) );
  CKAN2D1BWP30P140LVT U455 ( .A1(n104), .A2(i_data_bus[13]), .Z(n79) );
  CKAN2D1BWP30P140LVT U456 ( .A1(n104), .A2(i_data_bus[14]), .Z(n80) );
  CKAN2D1BWP30P140LVT U457 ( .A1(n104), .A2(i_data_bus[15]), .Z(n81) );
  CKAN2D1BWP30P140LVT U458 ( .A1(n104), .A2(i_data_bus[16]), .Z(n82) );
  CKAN2D1BWP30P140LVT U459 ( .A1(n104), .A2(i_data_bus[17]), .Z(n83) );
  CKAN2D1BWP30P140LVT U460 ( .A1(n104), .A2(i_data_bus[18]), .Z(n84) );
  CKAN2D1BWP30P140LVT U461 ( .A1(n104), .A2(i_data_bus[19]), .Z(n85) );
  CKAN2D1BWP30P140LVT U462 ( .A1(n104), .A2(i_data_bus[20]), .Z(n86) );
  CKAN2D1BWP30P140LVT U463 ( .A1(n104), .A2(i_data_bus[21]), .Z(n87) );
  CKAN2D1BWP30P140LVT U464 ( .A1(n104), .A2(i_data_bus[22]), .Z(n88) );
  CKAN2D1BWP30P140LVT U465 ( .A1(n104), .A2(i_data_bus[23]), .Z(n89) );
  CKAN2D1BWP30P140LVT U466 ( .A1(n104), .A2(i_data_bus[24]), .Z(n90) );
  CKAN2D1BWP30P140LVT U467 ( .A1(n104), .A2(i_data_bus[25]), .Z(n91) );
  CKAN2D1BWP30P140LVT U468 ( .A1(n105), .A2(o_data_forward_reg[26]), .Z(n92)
         );
  CKAN2D1BWP30P140LVT U469 ( .A1(n105), .A2(o_data_forward_reg[27]), .Z(n93)
         );
  CKAN2D1BWP30P140LVT U470 ( .A1(n105), .A2(o_data_forward_reg[28]), .Z(n94)
         );
  CKAN2D1BWP30P140LVT U471 ( .A1(n105), .A2(o_data_forward_reg[29]), .Z(n95)
         );
  CKAN2D1BWP30P140LVT U472 ( .A1(n105), .A2(o_data_forward_reg[30]), .Z(n96)
         );
  CKAN2D1BWP30P140LVT U473 ( .A1(n105), .A2(o_data_forward_reg[31]), .Z(n97)
         );
  CKAN2D1BWP30P140LVT U474 ( .A1(n104), .A2(i_data_bus[26]), .Z(n98) );
  CKAN2D1BWP30P140LVT U475 ( .A1(n104), .A2(i_data_bus[27]), .Z(n99) );
  CKAN2D1BWP30P140LVT U476 ( .A1(n104), .A2(i_data_bus[28]), .Z(n100) );
  CKAN2D1BWP30P140LVT U477 ( .A1(n104), .A2(i_data_bus[29]), .Z(n101) );
  CKAN2D1BWP30P140LVT U478 ( .A1(n104), .A2(i_data_bus[30]), .Z(n102) );
  CKAN2D1BWP30P140LVT U479 ( .A1(n104), .A2(i_data_bus[31]), .Z(n103) );
  CKAN2D1BWP30P140LVT U480 ( .A1(n7), .A2(o_cmd_forward_reg[2]), .Z(N420) );
  CKAN2D1BWP30P140LVT U481 ( .A1(n7), .A2(o_cmd_forward_reg[3]), .Z(N421) );
  CKAN2D1BWP30P140LVT U482 ( .A1(n7), .A2(i_cmd[0]), .Z(N147) );
  CKAN2D1BWP30P140LVT U483 ( .A1(n7), .A2(i_cmd[1]), .Z(N148) );
endmodule

