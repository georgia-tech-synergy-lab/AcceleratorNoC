

    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;
  tri   CLK;
  tri   rst;
  tri   i_en;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_0 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD4BWP30P140LVT U3 ( .I(n42), .ZN(n174) );
  NR2D3BWP30P140LVT U4 ( .A1(n32), .A2(n7), .ZN(n173) );
  INVD4BWP30P140LVT U5 ( .I(n16), .ZN(n170) );
  BUFFD4BWP30P140LVT U6 ( .I(n9), .Z(n172) );
  INVD4BWP30P140LVT U7 ( .I(n42), .ZN(n91) );
  INVD4BWP30P140LVT U8 ( .I(n2), .ZN(n3) );
  NR2D1BWP30P140LVT U9 ( .A1(n32), .A2(n8), .ZN(n9) );
  INVD1BWP30P140LVT U10 ( .I(n12), .ZN(n40) );
  INVD2BWP30P140LVT U11 ( .I(n33), .ZN(n2) );
  NR4D1BWP30P140LVT U12 ( .A1(n32), .A2(i_cmd[1]), .A3(n31), .A4(n30), .ZN(n33) );
  INVD0P7BWP30P140LVT U13 ( .I(i_cmd[0]), .ZN(n14) );
  CKND2D2BWP30P140LVT U14 ( .A1(n1), .A2(n22), .ZN(n32) );
  NR2D1BWP30P140LVT U15 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n10) );
  INVD1BWP30P140LVT U16 ( .I(i_cmd[6]), .ZN(n27) );
  INVD0P7BWP30P140LVT U17 ( .I(i_cmd[3]), .ZN(n18) );
  AOI22D1BWP30P140LVT U18 ( .A1(n175), .A2(i_data_bus[205]), .B1(n174), .B2(
        i_data_bus[173]), .ZN(n106) );
  CKAN2D1BWP30P140LVT U19 ( .A1(n27), .A2(n6), .Z(n1) );
  INVD1BWP30P140LVT U20 ( .I(i_cmd[4]), .ZN(n11) );
  NR3OPTPAD2BWP30P140LVT U21 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .A3(n5), .ZN(n6)
         );
  INVD2BWP30P140LVT U22 ( .I(n15), .ZN(n16) );
  INVD1BWP30P140LVT U23 ( .I(n29), .ZN(n41) );
  INVD2BWP30P140LVT U24 ( .I(n37), .ZN(n42) );
  NR4D1BWP30P140LVT U25 ( .A1(n36), .A2(i_cmd[6]), .A3(n35), .A4(n34), .ZN(n37) );
  INVD1BWP30P140LVT U26 ( .I(i_cmd[5]), .ZN(n35) );
  INVD1BWP30P140LVT U27 ( .I(i_cmd[2]), .ZN(n31) );
  NR2D3BWP30P140LVT U28 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n22) );
  IND3D2BWP30P140LVT U29 ( .A1(i_cmd[1]), .B1(n10), .B2(n1), .ZN(n13) );
  ND2D1BWP30P140LVT U30 ( .A1(n39), .A2(n38), .ZN(N402) );
  AN2D2BWP30P140LVT U31 ( .A1(n26), .A2(n25), .Z(n4) );
  INR2D1BWP30P140LVT U32 ( .A1(i_en), .B1(rst), .ZN(n17) );
  INVD1BWP30P140LVT U33 ( .I(n17), .ZN(n5) );
  ND3D1BWP30P140LVT U34 ( .A1(n10), .A2(i_valid[1]), .A3(i_cmd[1]), .ZN(n7) );
  NR2OPTPAD1BWP30P140LVT U35 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n19) );
  ND3D1BWP30P140LVT U36 ( .A1(n19), .A2(i_valid[3]), .A3(i_cmd[3]), .ZN(n8) );
  INR4D1BWP30P140LVT U37 ( .A1(i_valid[4]), .B1(i_cmd[0]), .B2(n11), .B3(n13), 
        .ZN(n12) );
  INVD2BWP30P140LVT U38 ( .I(n40), .ZN(n171) );
  INR4D1BWP30P140LVT U39 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n14), .B3(n13), 
        .ZN(n15) );
  NR4D0BWP30P140LVT U40 ( .A1(n173), .A2(n172), .A3(n171), .A4(n170), .ZN(n39)
         );
  CKAN2D1BWP30P140LVT U41 ( .A1(n18), .A2(n17), .Z(n20) );
  ND2OPTIBD1BWP30P140LVT U42 ( .A1(n20), .A2(n19), .ZN(n21) );
  INR2D2BWP30P140LVT U43 ( .A1(n22), .B1(n21), .ZN(n26) );
  INVD1BWP30P140LVT U44 ( .I(i_cmd[7]), .ZN(n24) );
  INVD1BWP30P140LVT U45 ( .I(i_valid[7]), .ZN(n23) );
  NR4D0BWP30P140LVT U46 ( .A1(i_cmd[6]), .A2(n24), .A3(i_cmd[5]), .A4(n23), 
        .ZN(n25) );
  INVD2BWP30P140LVT U47 ( .I(n26), .ZN(n36) );
  IND2D1BWP30P140LVT U48 ( .A1(i_cmd[7]), .B1(i_valid[6]), .ZN(n28) );
  NR4D1BWP30P140LVT U49 ( .A1(n36), .A2(i_cmd[5]), .A3(n28), .A4(n27), .ZN(n29) );
  INVD2BWP30P140LVT U50 ( .I(n41), .ZN(n165) );
  IND2D1BWP30P140LVT U51 ( .A1(i_cmd[3]), .B1(i_valid[2]), .ZN(n30) );
  IND2D1BWP30P140LVT U52 ( .A1(i_cmd[7]), .B1(i_valid[5]), .ZN(n34) );
  NR4D0BWP30P140LVT U53 ( .A1(n4), .A2(n165), .A3(n3), .A4(n174), .ZN(n38) );
  INVD2BWP30P140LVT U54 ( .I(n40), .ZN(n104) );
  AOI22D1BWP30P140LVT U55 ( .A1(n104), .A2(i_data_bus[140]), .B1(n170), .B2(
        i_data_bus[12]), .ZN(n46) );
  AOI22D1BWP30P140LVT U56 ( .A1(n173), .A2(i_data_bus[44]), .B1(n172), .B2(
        i_data_bus[108]), .ZN(n45) );
  INVD2BWP30P140LVT U57 ( .I(n41), .ZN(n175) );
  AOI22D1BWP30P140LVT U58 ( .A1(n175), .A2(i_data_bus[204]), .B1(n91), .B2(
        i_data_bus[172]), .ZN(n44) );
  AOI22D1BWP30P140LVT U59 ( .A1(n4), .A2(i_data_bus[236]), .B1(n3), .B2(
        i_data_bus[76]), .ZN(n43) );
  ND4D1BWP30P140LVT U60 ( .A1(n46), .A2(n45), .A3(n44), .A4(n43), .ZN(N381) );
  AOI22D1BWP30P140LVT U61 ( .A1(n104), .A2(i_data_bus[138]), .B1(n170), .B2(
        i_data_bus[10]), .ZN(n50) );
  AOI22D1BWP30P140LVT U62 ( .A1(n173), .A2(i_data_bus[42]), .B1(n172), .B2(
        i_data_bus[106]), .ZN(n49) );
  AOI22D1BWP30P140LVT U63 ( .A1(n175), .A2(i_data_bus[202]), .B1(n91), .B2(
        i_data_bus[170]), .ZN(n48) );
  AOI22D1BWP30P140LVT U64 ( .A1(n4), .A2(i_data_bus[234]), .B1(n3), .B2(
        i_data_bus[74]), .ZN(n47) );
  ND4D1BWP30P140LVT U65 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(N379) );
  AOI22D1BWP30P140LVT U66 ( .A1(n104), .A2(i_data_bus[137]), .B1(n170), .B2(
        i_data_bus[9]), .ZN(n54) );
  AOI22D1BWP30P140LVT U67 ( .A1(n173), .A2(i_data_bus[41]), .B1(n172), .B2(
        i_data_bus[105]), .ZN(n53) );
  AOI22D1BWP30P140LVT U68 ( .A1(n175), .A2(i_data_bus[201]), .B1(n91), .B2(
        i_data_bus[169]), .ZN(n52) );
  AOI22D1BWP30P140LVT U69 ( .A1(n4), .A2(i_data_bus[233]), .B1(n3), .B2(
        i_data_bus[73]), .ZN(n51) );
  ND4D1BWP30P140LVT U70 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(N378) );
  AOI22D1BWP30P140LVT U71 ( .A1(n104), .A2(i_data_bus[135]), .B1(n170), .B2(
        i_data_bus[7]), .ZN(n58) );
  AOI22D1BWP30P140LVT U72 ( .A1(n173), .A2(i_data_bus[39]), .B1(n172), .B2(
        i_data_bus[103]), .ZN(n57) );
  AOI22D1BWP30P140LVT U73 ( .A1(n175), .A2(i_data_bus[199]), .B1(n91), .B2(
        i_data_bus[167]), .ZN(n56) );
  AOI22D1BWP30P140LVT U74 ( .A1(n4), .A2(i_data_bus[231]), .B1(n3), .B2(
        i_data_bus[71]), .ZN(n55) );
  ND4D1BWP30P140LVT U75 ( .A1(n58), .A2(n57), .A3(n56), .A4(n55), .ZN(N376) );
  AOI22D1BWP30P140LVT U76 ( .A1(n104), .A2(i_data_bus[134]), .B1(n170), .B2(
        i_data_bus[6]), .ZN(n62) );
  AOI22D1BWP30P140LVT U77 ( .A1(n173), .A2(i_data_bus[38]), .B1(n172), .B2(
        i_data_bus[102]), .ZN(n61) );
  AOI22D1BWP30P140LVT U78 ( .A1(n175), .A2(i_data_bus[198]), .B1(n91), .B2(
        i_data_bus[166]), .ZN(n60) );
  AOI22D1BWP30P140LVT U79 ( .A1(n4), .A2(i_data_bus[230]), .B1(n3), .B2(
        i_data_bus[70]), .ZN(n59) );
  ND4D1BWP30P140LVT U80 ( .A1(n62), .A2(n61), .A3(n60), .A4(n59), .ZN(N375) );
  AOI22D1BWP30P140LVT U81 ( .A1(n104), .A2(i_data_bus[132]), .B1(n170), .B2(
        i_data_bus[4]), .ZN(n66) );
  AOI22D1BWP30P140LVT U82 ( .A1(n173), .A2(i_data_bus[36]), .B1(n172), .B2(
        i_data_bus[100]), .ZN(n65) );
  AOI22D1BWP30P140LVT U83 ( .A1(n175), .A2(i_data_bus[196]), .B1(n91), .B2(
        i_data_bus[164]), .ZN(n64) );
  AOI22D1BWP30P140LVT U84 ( .A1(n4), .A2(i_data_bus[228]), .B1(n3), .B2(
        i_data_bus[68]), .ZN(n63) );
  ND4D1BWP30P140LVT U85 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(N373) );
  AOI22D1BWP30P140LVT U86 ( .A1(n104), .A2(i_data_bus[131]), .B1(n170), .B2(
        i_data_bus[3]), .ZN(n70) );
  AOI22D1BWP30P140LVT U87 ( .A1(n173), .A2(i_data_bus[35]), .B1(n172), .B2(
        i_data_bus[99]), .ZN(n69) );
  AOI22D1BWP30P140LVT U88 ( .A1(n175), .A2(i_data_bus[195]), .B1(n91), .B2(
        i_data_bus[163]), .ZN(n68) );
  AOI22D1BWP30P140LVT U89 ( .A1(n4), .A2(i_data_bus[227]), .B1(n3), .B2(
        i_data_bus[67]), .ZN(n67) );
  ND4D1BWP30P140LVT U90 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(N372) );
  AOI22D1BWP30P140LVT U91 ( .A1(n104), .A2(i_data_bus[129]), .B1(n170), .B2(
        i_data_bus[1]), .ZN(n74) );
  AOI22D1BWP30P140LVT U92 ( .A1(n173), .A2(i_data_bus[33]), .B1(n172), .B2(
        i_data_bus[97]), .ZN(n73) );
  AOI22D1BWP30P140LVT U93 ( .A1(n175), .A2(i_data_bus[193]), .B1(n91), .B2(
        i_data_bus[161]), .ZN(n72) );
  AOI22D1BWP30P140LVT U94 ( .A1(n4), .A2(i_data_bus[225]), .B1(n3), .B2(
        i_data_bus[65]), .ZN(n71) );
  ND4D1BWP30P140LVT U95 ( .A1(n74), .A2(n73), .A3(n72), .A4(n71), .ZN(N370) );
  AOI22D1BWP30P140LVT U96 ( .A1(n104), .A2(i_data_bus[139]), .B1(n170), .B2(
        i_data_bus[11]), .ZN(n78) );
  AOI22D1BWP30P140LVT U97 ( .A1(n173), .A2(i_data_bus[43]), .B1(n172), .B2(
        i_data_bus[107]), .ZN(n77) );
  AOI22D1BWP30P140LVT U98 ( .A1(n175), .A2(i_data_bus[203]), .B1(n91), .B2(
        i_data_bus[171]), .ZN(n76) );
  AOI22D1BWP30P140LVT U99 ( .A1(n4), .A2(i_data_bus[235]), .B1(n3), .B2(
        i_data_bus[75]), .ZN(n75) );
  ND4D1BWP30P140LVT U100 ( .A1(n78), .A2(n77), .A3(n76), .A4(n75), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U101 ( .A1(n104), .A2(i_data_bus[136]), .B1(n170), .B2(
        i_data_bus[8]), .ZN(n82) );
  AOI22D1BWP30P140LVT U102 ( .A1(n173), .A2(i_data_bus[40]), .B1(n172), .B2(
        i_data_bus[104]), .ZN(n81) );
  AOI22D1BWP30P140LVT U103 ( .A1(n175), .A2(i_data_bus[200]), .B1(n91), .B2(
        i_data_bus[168]), .ZN(n80) );
  AOI22D1BWP30P140LVT U104 ( .A1(n4), .A2(i_data_bus[232]), .B1(n3), .B2(
        i_data_bus[72]), .ZN(n79) );
  ND4D1BWP30P140LVT U105 ( .A1(n82), .A2(n81), .A3(n80), .A4(n79), .ZN(N377)
         );
  AOI22D1BWP30P140LVT U106 ( .A1(n104), .A2(i_data_bus[133]), .B1(n170), .B2(
        i_data_bus[5]), .ZN(n86) );
  AOI22D1BWP30P140LVT U107 ( .A1(n173), .A2(i_data_bus[37]), .B1(n172), .B2(
        i_data_bus[101]), .ZN(n85) );
  AOI22D1BWP30P140LVT U108 ( .A1(n175), .A2(i_data_bus[197]), .B1(n91), .B2(
        i_data_bus[165]), .ZN(n84) );
  AOI22D1BWP30P140LVT U109 ( .A1(n4), .A2(i_data_bus[229]), .B1(n3), .B2(
        i_data_bus[69]), .ZN(n83) );
  ND4D1BWP30P140LVT U110 ( .A1(n86), .A2(n85), .A3(n84), .A4(n83), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U111 ( .A1(n104), .A2(i_data_bus[130]), .B1(n170), .B2(
        i_data_bus[2]), .ZN(n90) );
  AOI22D1BWP30P140LVT U112 ( .A1(n173), .A2(i_data_bus[34]), .B1(n172), .B2(
        i_data_bus[98]), .ZN(n89) );
  AOI22D1BWP30P140LVT U113 ( .A1(n175), .A2(i_data_bus[194]), .B1(n91), .B2(
        i_data_bus[162]), .ZN(n88) );
  AOI22D1BWP30P140LVT U114 ( .A1(n4), .A2(i_data_bus[226]), .B1(n3), .B2(
        i_data_bus[66]), .ZN(n87) );
  ND4D1BWP30P140LVT U115 ( .A1(n90), .A2(n89), .A3(n88), .A4(n87), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U116 ( .A1(n104), .A2(i_data_bus[128]), .B1(n170), .B2(
        i_data_bus[0]), .ZN(n95) );
  AOI22D1BWP30P140LVT U117 ( .A1(n173), .A2(i_data_bus[32]), .B1(n172), .B2(
        i_data_bus[96]), .ZN(n94) );
  AOI22D1BWP30P140LVT U118 ( .A1(n165), .A2(i_data_bus[192]), .B1(n91), .B2(
        i_data_bus[160]), .ZN(n93) );
  AOI22D1BWP30P140LVT U119 ( .A1(n4), .A2(i_data_bus[224]), .B1(n3), .B2(
        i_data_bus[64]), .ZN(n92) );
  ND4D1BWP30P140LVT U120 ( .A1(n95), .A2(n94), .A3(n93), .A4(n92), .ZN(N369)
         );
  AOI22D1BWP30P140LVT U121 ( .A1(n104), .A2(i_data_bus[143]), .B1(n170), .B2(
        i_data_bus[15]), .ZN(n99) );
  AOI22D1BWP30P140LVT U122 ( .A1(n173), .A2(i_data_bus[47]), .B1(n172), .B2(
        i_data_bus[111]), .ZN(n98) );
  AOI22D1BWP30P140LVT U123 ( .A1(n175), .A2(i_data_bus[207]), .B1(n174), .B2(
        i_data_bus[175]), .ZN(n97) );
  AOI22D1BWP30P140LVT U124 ( .A1(n4), .A2(i_data_bus[239]), .B1(n3), .B2(
        i_data_bus[79]), .ZN(n96) );
  ND4D1BWP30P140LVT U125 ( .A1(n99), .A2(n98), .A3(n97), .A4(n96), .ZN(N384)
         );
  AOI22D1BWP30P140LVT U126 ( .A1(n104), .A2(i_data_bus[142]), .B1(n170), .B2(
        i_data_bus[14]), .ZN(n103) );
  AOI22D1BWP30P140LVT U127 ( .A1(n173), .A2(i_data_bus[46]), .B1(n172), .B2(
        i_data_bus[110]), .ZN(n102) );
  AOI22D1BWP30P140LVT U128 ( .A1(n175), .A2(i_data_bus[206]), .B1(n174), .B2(
        i_data_bus[174]), .ZN(n101) );
  AOI22D1BWP30P140LVT U129 ( .A1(n4), .A2(i_data_bus[238]), .B1(n3), .B2(
        i_data_bus[78]), .ZN(n100) );
  ND4D1BWP30P140LVT U130 ( .A1(n103), .A2(n102), .A3(n101), .A4(n100), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U131 ( .A1(n104), .A2(i_data_bus[141]), .B1(n170), .B2(
        i_data_bus[13]), .ZN(n108) );
  AOI22D1BWP30P140LVT U132 ( .A1(n173), .A2(i_data_bus[45]), .B1(n172), .B2(
        i_data_bus[109]), .ZN(n107) );
  AOI22D1BWP30P140LVT U133 ( .A1(n4), .A2(i_data_bus[237]), .B1(n3), .B2(
        i_data_bus[77]), .ZN(n105) );
  ND4D1BWP30P140LVT U134 ( .A1(n108), .A2(n107), .A3(n106), .A4(n105), .ZN(
        N382) );
  AOI22D1BWP30P140LVT U135 ( .A1(n171), .A2(i_data_bus[159]), .B1(n170), .B2(
        i_data_bus[31]), .ZN(n112) );
  AOI22D1BWP30P140LVT U136 ( .A1(n173), .A2(i_data_bus[63]), .B1(n172), .B2(
        i_data_bus[127]), .ZN(n111) );
  AOI22D1BWP30P140LVT U137 ( .A1(n165), .A2(i_data_bus[223]), .B1(n174), .B2(
        i_data_bus[191]), .ZN(n110) );
  AOI22D1BWP30P140LVT U138 ( .A1(n4), .A2(i_data_bus[255]), .B1(n3), .B2(
        i_data_bus[95]), .ZN(n109) );
  ND4D1BWP30P140LVT U139 ( .A1(n112), .A2(n111), .A3(n110), .A4(n109), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U140 ( .A1(n171), .A2(i_data_bus[158]), .B1(n170), .B2(
        i_data_bus[30]), .ZN(n116) );
  AOI22D1BWP30P140LVT U141 ( .A1(n173), .A2(i_data_bus[62]), .B1(n172), .B2(
        i_data_bus[126]), .ZN(n115) );
  AOI22D1BWP30P140LVT U142 ( .A1(n165), .A2(i_data_bus[222]), .B1(n174), .B2(
        i_data_bus[190]), .ZN(n114) );
  AOI22D1BWP30P140LVT U143 ( .A1(n4), .A2(i_data_bus[254]), .B1(n3), .B2(
        i_data_bus[94]), .ZN(n113) );
  ND4D1BWP30P140LVT U144 ( .A1(n116), .A2(n115), .A3(n114), .A4(n113), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U145 ( .A1(n171), .A2(i_data_bus[157]), .B1(n170), .B2(
        i_data_bus[29]), .ZN(n120) );
  AOI22D1BWP30P140LVT U146 ( .A1(n173), .A2(i_data_bus[61]), .B1(n172), .B2(
        i_data_bus[125]), .ZN(n119) );
  AOI22D1BWP30P140LVT U147 ( .A1(n165), .A2(i_data_bus[221]), .B1(n174), .B2(
        i_data_bus[189]), .ZN(n118) );
  AOI22D1BWP30P140LVT U148 ( .A1(n4), .A2(i_data_bus[253]), .B1(n3), .B2(
        i_data_bus[93]), .ZN(n117) );
  ND4D1BWP30P140LVT U149 ( .A1(n120), .A2(n119), .A3(n118), .A4(n117), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U150 ( .A1(n171), .A2(i_data_bus[156]), .B1(n170), .B2(
        i_data_bus[28]), .ZN(n124) );
  AOI22D1BWP30P140LVT U151 ( .A1(n173), .A2(i_data_bus[60]), .B1(n172), .B2(
        i_data_bus[124]), .ZN(n123) );
  AOI22D1BWP30P140LVT U152 ( .A1(n165), .A2(i_data_bus[220]), .B1(n174), .B2(
        i_data_bus[188]), .ZN(n122) );
  AOI22D1BWP30P140LVT U153 ( .A1(n4), .A2(i_data_bus[252]), .B1(n3), .B2(
        i_data_bus[92]), .ZN(n121) );
  ND4D1BWP30P140LVT U154 ( .A1(n124), .A2(n123), .A3(n122), .A4(n121), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U155 ( .A1(n171), .A2(i_data_bus[155]), .B1(n170), .B2(
        i_data_bus[27]), .ZN(n128) );
  AOI22D1BWP30P140LVT U156 ( .A1(n173), .A2(i_data_bus[59]), .B1(n172), .B2(
        i_data_bus[123]), .ZN(n127) );
  AOI22D1BWP30P140LVT U157 ( .A1(n165), .A2(i_data_bus[219]), .B1(n174), .B2(
        i_data_bus[187]), .ZN(n126) );
  AOI22D1BWP30P140LVT U158 ( .A1(n4), .A2(i_data_bus[251]), .B1(n3), .B2(
        i_data_bus[91]), .ZN(n125) );
  ND4D1BWP30P140LVT U159 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U160 ( .A1(n171), .A2(i_data_bus[154]), .B1(n170), .B2(
        i_data_bus[26]), .ZN(n132) );
  AOI22D1BWP30P140LVT U161 ( .A1(n173), .A2(i_data_bus[58]), .B1(n172), .B2(
        i_data_bus[122]), .ZN(n131) );
  AOI22D1BWP30P140LVT U162 ( .A1(n165), .A2(i_data_bus[218]), .B1(n174), .B2(
        i_data_bus[186]), .ZN(n130) );
  AOI22D1BWP30P140LVT U163 ( .A1(n4), .A2(i_data_bus[250]), .B1(n3), .B2(
        i_data_bus[90]), .ZN(n129) );
  ND4D1BWP30P140LVT U164 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U165 ( .A1(n171), .A2(i_data_bus[153]), .B1(n170), .B2(
        i_data_bus[25]), .ZN(n136) );
  AOI22D1BWP30P140LVT U166 ( .A1(n173), .A2(i_data_bus[57]), .B1(n172), .B2(
        i_data_bus[121]), .ZN(n135) );
  AOI22D1BWP30P140LVT U167 ( .A1(n165), .A2(i_data_bus[217]), .B1(n174), .B2(
        i_data_bus[185]), .ZN(n134) );
  AOI22D1BWP30P140LVT U168 ( .A1(n4), .A2(i_data_bus[249]), .B1(n3), .B2(
        i_data_bus[89]), .ZN(n133) );
  ND4D1BWP30P140LVT U169 ( .A1(n136), .A2(n135), .A3(n134), .A4(n133), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U170 ( .A1(n171), .A2(i_data_bus[152]), .B1(n170), .B2(
        i_data_bus[24]), .ZN(n140) );
  AOI22D1BWP30P140LVT U171 ( .A1(n173), .A2(i_data_bus[56]), .B1(n172), .B2(
        i_data_bus[120]), .ZN(n139) );
  AOI22D1BWP30P140LVT U172 ( .A1(n165), .A2(i_data_bus[216]), .B1(n174), .B2(
        i_data_bus[184]), .ZN(n138) );
  AOI22D1BWP30P140LVT U173 ( .A1(n4), .A2(i_data_bus[248]), .B1(n3), .B2(
        i_data_bus[88]), .ZN(n137) );
  ND4D1BWP30P140LVT U174 ( .A1(n140), .A2(n139), .A3(n138), .A4(n137), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U175 ( .A1(n171), .A2(i_data_bus[151]), .B1(n170), .B2(
        i_data_bus[23]), .ZN(n144) );
  AOI22D1BWP30P140LVT U176 ( .A1(n173), .A2(i_data_bus[55]), .B1(n172), .B2(
        i_data_bus[119]), .ZN(n143) );
  AOI22D1BWP30P140LVT U177 ( .A1(n165), .A2(i_data_bus[215]), .B1(n174), .B2(
        i_data_bus[183]), .ZN(n142) );
  AOI22D1BWP30P140LVT U178 ( .A1(n4), .A2(i_data_bus[247]), .B1(n3), .B2(
        i_data_bus[87]), .ZN(n141) );
  ND4D1BWP30P140LVT U179 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U180 ( .A1(n171), .A2(i_data_bus[150]), .B1(n170), .B2(
        i_data_bus[22]), .ZN(n148) );
  AOI22D1BWP30P140LVT U181 ( .A1(n173), .A2(i_data_bus[54]), .B1(n172), .B2(
        i_data_bus[118]), .ZN(n147) );
  AOI22D1BWP30P140LVT U182 ( .A1(n165), .A2(i_data_bus[214]), .B1(n174), .B2(
        i_data_bus[182]), .ZN(n146) );
  AOI22D1BWP30P140LVT U183 ( .A1(n4), .A2(i_data_bus[246]), .B1(n3), .B2(
        i_data_bus[86]), .ZN(n145) );
  ND4D1BWP30P140LVT U184 ( .A1(n148), .A2(n147), .A3(n146), .A4(n145), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U185 ( .A1(n171), .A2(i_data_bus[149]), .B1(n170), .B2(
        i_data_bus[21]), .ZN(n152) );
  AOI22D1BWP30P140LVT U186 ( .A1(n173), .A2(i_data_bus[53]), .B1(n172), .B2(
        i_data_bus[117]), .ZN(n151) );
  AOI22D1BWP30P140LVT U187 ( .A1(n165), .A2(i_data_bus[213]), .B1(n174), .B2(
        i_data_bus[181]), .ZN(n150) );
  AOI22D1BWP30P140LVT U188 ( .A1(n4), .A2(i_data_bus[245]), .B1(n3), .B2(
        i_data_bus[85]), .ZN(n149) );
  ND4D1BWP30P140LVT U189 ( .A1(n152), .A2(n151), .A3(n150), .A4(n149), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U190 ( .A1(n171), .A2(i_data_bus[148]), .B1(n170), .B2(
        i_data_bus[20]), .ZN(n156) );
  AOI22D1BWP30P140LVT U191 ( .A1(n173), .A2(i_data_bus[52]), .B1(n172), .B2(
        i_data_bus[116]), .ZN(n155) );
  AOI22D1BWP30P140LVT U192 ( .A1(n165), .A2(i_data_bus[212]), .B1(n174), .B2(
        i_data_bus[180]), .ZN(n154) );
  AOI22D1BWP30P140LVT U193 ( .A1(n4), .A2(i_data_bus[244]), .B1(n3), .B2(
        i_data_bus[84]), .ZN(n153) );
  ND4D1BWP30P140LVT U194 ( .A1(n156), .A2(n155), .A3(n154), .A4(n153), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U195 ( .A1(n171), .A2(i_data_bus[147]), .B1(n170), .B2(
        i_data_bus[19]), .ZN(n160) );
  AOI22D1BWP30P140LVT U196 ( .A1(n173), .A2(i_data_bus[51]), .B1(n172), .B2(
        i_data_bus[115]), .ZN(n159) );
  AOI22D1BWP30P140LVT U197 ( .A1(n165), .A2(i_data_bus[211]), .B1(n174), .B2(
        i_data_bus[179]), .ZN(n158) );
  AOI22D1BWP30P140LVT U198 ( .A1(n4), .A2(i_data_bus[243]), .B1(n3), .B2(
        i_data_bus[83]), .ZN(n157) );
  ND4D1BWP30P140LVT U199 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U200 ( .A1(n171), .A2(i_data_bus[146]), .B1(n170), .B2(
        i_data_bus[18]), .ZN(n164) );
  AOI22D1BWP30P140LVT U201 ( .A1(n173), .A2(i_data_bus[50]), .B1(n172), .B2(
        i_data_bus[114]), .ZN(n163) );
  AOI22D1BWP30P140LVT U202 ( .A1(n165), .A2(i_data_bus[210]), .B1(n174), .B2(
        i_data_bus[178]), .ZN(n162) );
  AOI22D1BWP30P140LVT U203 ( .A1(n4), .A2(i_data_bus[242]), .B1(n3), .B2(
        i_data_bus[82]), .ZN(n161) );
  ND4D1BWP30P140LVT U204 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U205 ( .A1(n171), .A2(i_data_bus[145]), .B1(n170), .B2(
        i_data_bus[17]), .ZN(n169) );
  AOI22D1BWP30P140LVT U206 ( .A1(n173), .A2(i_data_bus[49]), .B1(n172), .B2(
        i_data_bus[113]), .ZN(n168) );
  AOI22D1BWP30P140LVT U207 ( .A1(n165), .A2(i_data_bus[209]), .B1(n174), .B2(
        i_data_bus[177]), .ZN(n167) );
  AOI22D1BWP30P140LVT U208 ( .A1(n4), .A2(i_data_bus[241]), .B1(n3), .B2(
        i_data_bus[81]), .ZN(n166) );
  ND4D1BWP30P140LVT U209 ( .A1(n169), .A2(n168), .A3(n167), .A4(n166), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U210 ( .A1(n171), .A2(i_data_bus[144]), .B1(n170), .B2(
        i_data_bus[16]), .ZN(n179) );
  AOI22D1BWP30P140LVT U211 ( .A1(n173), .A2(i_data_bus[48]), .B1(n172), .B2(
        i_data_bus[112]), .ZN(n178) );
  AOI22D1BWP30P140LVT U212 ( .A1(n175), .A2(i_data_bus[208]), .B1(n174), .B2(
        i_data_bus[176]), .ZN(n177) );
  AOI22D1BWP30P140LVT U213 ( .A1(n4), .A2(i_data_bus[240]), .B1(n3), .B2(
        i_data_bus[80]), .ZN(n176) );
  ND4D1BWP30P140LVT U214 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(
        N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_1 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  DFQD2BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  INVD3BWP30P140LVT U3 ( .I(n12), .ZN(n173) );
  INVD1BWP30P140LVT U4 ( .I(n4), .ZN(n5) );
  INVD1BWP30P140LVT U5 ( .I(n23), .ZN(n24) );
  INR2D1BWP30P140LVT U6 ( .A1(n29), .B1(n3), .ZN(n4) );
  INR2D1BWP30P140LVT U7 ( .A1(n25), .B1(n22), .ZN(n23) );
  NR2D1BWP30P140LVT U8 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n18) );
  NR2D2BWP30P140LVT U9 ( .A1(i_cmd[6]), .A2(i_cmd[5]), .ZN(n21) );
  INR2D1BWP30P140LVT U10 ( .A1(n16), .B1(i_cmd[7]), .ZN(n2) );
  ND2OPTIBD2BWP30P140LVT U11 ( .A1(n21), .A2(n2), .ZN(n7) );
  INVD1BWP30P140LVT U12 ( .I(n11), .ZN(n12) );
  INVD6BWP30P140LVT U13 ( .I(n24), .ZN(n178) );
  INVD8BWP30P140LVT U14 ( .I(n42), .ZN(n1) );
  INVD6BWP30P140LVT U15 ( .I(n5), .ZN(n175) );
  INVD1BWP30P140LVT U16 ( .I(i_cmd[2]), .ZN(n31) );
  INVD1BWP30P140LVT U17 ( .I(i_cmd[6]), .ZN(n26) );
  INVD1BWP30P140LVT U18 ( .I(i_cmd[4]), .ZN(n10) );
  INVD3BWP30P140LVT U19 ( .I(n40), .ZN(n172) );
  INVD1BWP30P140LVT U20 ( .I(i_cmd[5]), .ZN(n35) );
  INVD1BWP30P140LVT U21 ( .I(n15), .ZN(n40) );
  INVD1BWP30P140LVT U22 ( .I(i_cmd[0]), .ZN(n14) );
  INVD1BWP30P140LVT U23 ( .I(n29), .ZN(n32) );
  INR2D4BWP30P140LVT U24 ( .A1(n29), .B1(n6), .ZN(n174) );
  ND2D1BWP30P140LVT U25 ( .A1(n39), .A2(n38), .ZN(N402) );
  INR2D1BWP30P140LVT U26 ( .A1(i_en), .B1(rst), .ZN(n16) );
  INR2D2BWP30P140LVT U27 ( .A1(n18), .B1(n7), .ZN(n29) );
  NR2OPTPAD1BWP30P140LVT U28 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n9) );
  ND3D1BWP30P140LVT U29 ( .A1(n9), .A2(i_cmd[1]), .A3(i_valid[1]), .ZN(n3) );
  NR2OPTPAD1BWP30P140LVT U30 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n20) );
  ND3D1BWP30P140LVT U31 ( .A1(n20), .A2(i_valid[3]), .A3(i_cmd[3]), .ZN(n6) );
  INVD2BWP30P140LVT U32 ( .I(n7), .ZN(n8) );
  IND3D2BWP30P140LVT U33 ( .A1(i_cmd[1]), .B1(n9), .B2(n8), .ZN(n13) );
  INR4D1BWP30P140LVT U34 ( .A1(i_valid[4]), .B1(i_cmd[0]), .B2(n10), .B3(n13), 
        .ZN(n11) );
  INR4D1BWP30P140LVT U35 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n14), .B3(n13), 
        .ZN(n15) );
  NR4D0BWP30P140LVT U36 ( .A1(n175), .A2(n174), .A3(n173), .A4(n172), .ZN(n39)
         );
  INR2D1BWP30P140LVT U37 ( .A1(n16), .B1(i_cmd[3]), .ZN(n17) );
  ND2OPTIBD1BWP30P140LVT U38 ( .A1(n18), .A2(n17), .ZN(n19) );
  INR2D2BWP30P140LVT U39 ( .A1(n20), .B1(n19), .ZN(n25) );
  ND3D1BWP30P140LVT U40 ( .A1(n21), .A2(i_valid[7]), .A3(i_cmd[7]), .ZN(n22)
         );
  INVD2BWP30P140LVT U41 ( .I(n25), .ZN(n36) );
  IND2D1BWP30P140LVT U42 ( .A1(i_cmd[7]), .B1(i_valid[6]), .ZN(n27) );
  NR4D1BWP30P140LVT U43 ( .A1(n36), .A2(i_cmd[5]), .A3(n27), .A4(n26), .ZN(n28) );
  INVD2BWP30P140LVT U44 ( .I(n28), .ZN(n71) );
  INVD2BWP30P140LVT U45 ( .I(n71), .ZN(n167) );
  IND2D1BWP30P140LVT U46 ( .A1(i_cmd[3]), .B1(i_valid[2]), .ZN(n30) );
  NR4D2BWP30P140LVT U47 ( .A1(n32), .A2(i_cmd[1]), .A3(n31), .A4(n30), .ZN(n33) );
  INVD3BWP30P140LVT U48 ( .I(n33), .ZN(n42) );
  IND2D1BWP30P140LVT U49 ( .A1(i_cmd[7]), .B1(i_valid[5]), .ZN(n34) );
  NR4D1BWP30P140LVT U50 ( .A1(n36), .A2(i_cmd[6]), .A3(n35), .A4(n34), .ZN(n37) );
  INVD2BWP30P140LVT U51 ( .I(n37), .ZN(n41) );
  INVD6BWP30P140LVT U52 ( .I(n41), .ZN(n176) );
  NR4D0BWP30P140LVT U53 ( .A1(n178), .A2(n167), .A3(n1), .A4(n176), .ZN(n38)
         );
  INVD2BWP30P140LVT U54 ( .I(n40), .ZN(n93) );
  AOI22D1BWP30P140LVT U55 ( .A1(n173), .A2(i_data_bus[140]), .B1(n93), .B2(
        i_data_bus[12]), .ZN(n46) );
  AOI22D1BWP30P140LVT U56 ( .A1(n175), .A2(i_data_bus[44]), .B1(n174), .B2(
        i_data_bus[108]), .ZN(n45) );
  INVD2BWP30P140LVT U57 ( .I(n71), .ZN(n177) );
  INVD4BWP30P140LVT U58 ( .I(n41), .ZN(n94) );
  AOI22D1BWP30P140LVT U59 ( .A1(n177), .A2(i_data_bus[204]), .B1(n94), .B2(
        i_data_bus[172]), .ZN(n44) );
  AOI22D1BWP30P140LVT U60 ( .A1(n178), .A2(i_data_bus[236]), .B1(n1), .B2(
        i_data_bus[76]), .ZN(n43) );
  ND4D1BWP30P140LVT U61 ( .A1(n46), .A2(n45), .A3(n44), .A4(n43), .ZN(N381) );
  AOI22D1BWP30P140LVT U62 ( .A1(n173), .A2(i_data_bus[138]), .B1(n93), .B2(
        i_data_bus[10]), .ZN(n50) );
  AOI22D1BWP30P140LVT U63 ( .A1(n175), .A2(i_data_bus[42]), .B1(n174), .B2(
        i_data_bus[106]), .ZN(n49) );
  AOI22D1BWP30P140LVT U64 ( .A1(n177), .A2(i_data_bus[202]), .B1(n94), .B2(
        i_data_bus[170]), .ZN(n48) );
  AOI22D1BWP30P140LVT U65 ( .A1(n178), .A2(i_data_bus[234]), .B1(n1), .B2(
        i_data_bus[74]), .ZN(n47) );
  ND4D1BWP30P140LVT U66 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(N379) );
  AOI22D1BWP30P140LVT U67 ( .A1(n173), .A2(i_data_bus[137]), .B1(n93), .B2(
        i_data_bus[9]), .ZN(n54) );
  AOI22D1BWP30P140LVT U68 ( .A1(n175), .A2(i_data_bus[41]), .B1(n174), .B2(
        i_data_bus[105]), .ZN(n53) );
  AOI22D1BWP30P140LVT U69 ( .A1(n177), .A2(i_data_bus[201]), .B1(n94), .B2(
        i_data_bus[169]), .ZN(n52) );
  AOI22D1BWP30P140LVT U70 ( .A1(n178), .A2(i_data_bus[233]), .B1(n1), .B2(
        i_data_bus[73]), .ZN(n51) );
  ND4D1BWP30P140LVT U71 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(N378) );
  AOI22D1BWP30P140LVT U72 ( .A1(n173), .A2(i_data_bus[135]), .B1(n93), .B2(
        i_data_bus[7]), .ZN(n58) );
  AOI22D1BWP30P140LVT U73 ( .A1(n175), .A2(i_data_bus[39]), .B1(n174), .B2(
        i_data_bus[103]), .ZN(n57) );
  AOI22D1BWP30P140LVT U74 ( .A1(n177), .A2(i_data_bus[199]), .B1(n94), .B2(
        i_data_bus[167]), .ZN(n56) );
  AOI22D1BWP30P140LVT U75 ( .A1(n178), .A2(i_data_bus[231]), .B1(n1), .B2(
        i_data_bus[71]), .ZN(n55) );
  ND4D1BWP30P140LVT U76 ( .A1(n58), .A2(n57), .A3(n56), .A4(n55), .ZN(N376) );
  AOI22D1BWP30P140LVT U77 ( .A1(n173), .A2(i_data_bus[134]), .B1(n93), .B2(
        i_data_bus[6]), .ZN(n62) );
  AOI22D1BWP30P140LVT U78 ( .A1(n175), .A2(i_data_bus[38]), .B1(n174), .B2(
        i_data_bus[102]), .ZN(n61) );
  AOI22D1BWP30P140LVT U79 ( .A1(n177), .A2(i_data_bus[198]), .B1(n94), .B2(
        i_data_bus[166]), .ZN(n60) );
  AOI22D1BWP30P140LVT U80 ( .A1(n178), .A2(i_data_bus[230]), .B1(n1), .B2(
        i_data_bus[70]), .ZN(n59) );
  ND4D1BWP30P140LVT U81 ( .A1(n62), .A2(n61), .A3(n60), .A4(n59), .ZN(N375) );
  AOI22D1BWP30P140LVT U82 ( .A1(n173), .A2(i_data_bus[132]), .B1(n93), .B2(
        i_data_bus[4]), .ZN(n66) );
  AOI22D1BWP30P140LVT U83 ( .A1(n175), .A2(i_data_bus[36]), .B1(n174), .B2(
        i_data_bus[100]), .ZN(n65) );
  AOI22D1BWP30P140LVT U84 ( .A1(n177), .A2(i_data_bus[196]), .B1(n94), .B2(
        i_data_bus[164]), .ZN(n64) );
  AOI22D1BWP30P140LVT U85 ( .A1(n178), .A2(i_data_bus[228]), .B1(n1), .B2(
        i_data_bus[68]), .ZN(n63) );
  ND4D1BWP30P140LVT U86 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(N373) );
  AOI22D1BWP30P140LVT U87 ( .A1(n173), .A2(i_data_bus[131]), .B1(n93), .B2(
        i_data_bus[3]), .ZN(n70) );
  AOI22D1BWP30P140LVT U88 ( .A1(n175), .A2(i_data_bus[35]), .B1(n174), .B2(
        i_data_bus[99]), .ZN(n69) );
  AOI22D1BWP30P140LVT U89 ( .A1(n177), .A2(i_data_bus[195]), .B1(n94), .B2(
        i_data_bus[163]), .ZN(n68) );
  AOI22D1BWP30P140LVT U90 ( .A1(n178), .A2(i_data_bus[227]), .B1(n1), .B2(
        i_data_bus[67]), .ZN(n67) );
  ND4D1BWP30P140LVT U91 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(N372) );
  AOI22D1BWP30P140LVT U92 ( .A1(n173), .A2(i_data_bus[128]), .B1(n93), .B2(
        i_data_bus[0]), .ZN(n76) );
  AOI22D1BWP30P140LVT U93 ( .A1(n175), .A2(i_data_bus[32]), .B1(n174), .B2(
        i_data_bus[96]), .ZN(n75) );
  INVD1BWP30P140LVT U94 ( .I(n71), .ZN(n72) );
  AOI22D1BWP30P140LVT U95 ( .A1(n72), .A2(i_data_bus[192]), .B1(n94), .B2(
        i_data_bus[160]), .ZN(n74) );
  AOI22D1BWP30P140LVT U96 ( .A1(n178), .A2(i_data_bus[224]), .B1(n1), .B2(
        i_data_bus[64]), .ZN(n73) );
  ND4D1BWP30P140LVT U97 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(N369) );
  AOI22D1BWP30P140LVT U98 ( .A1(n173), .A2(i_data_bus[139]), .B1(n93), .B2(
        i_data_bus[11]), .ZN(n80) );
  AOI22D1BWP30P140LVT U99 ( .A1(n175), .A2(i_data_bus[43]), .B1(n174), .B2(
        i_data_bus[107]), .ZN(n79) );
  AOI22D1BWP30P140LVT U100 ( .A1(n177), .A2(i_data_bus[203]), .B1(n94), .B2(
        i_data_bus[171]), .ZN(n78) );
  AOI22D1BWP30P140LVT U101 ( .A1(n178), .A2(i_data_bus[235]), .B1(n1), .B2(
        i_data_bus[75]), .ZN(n77) );
  ND4D1BWP30P140LVT U102 ( .A1(n80), .A2(n79), .A3(n78), .A4(n77), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U103 ( .A1(n173), .A2(i_data_bus[136]), .B1(n93), .B2(
        i_data_bus[8]), .ZN(n84) );
  AOI22D1BWP30P140LVT U104 ( .A1(n175), .A2(i_data_bus[40]), .B1(n174), .B2(
        i_data_bus[104]), .ZN(n83) );
  AOI22D1BWP30P140LVT U105 ( .A1(n177), .A2(i_data_bus[200]), .B1(n94), .B2(
        i_data_bus[168]), .ZN(n82) );
  AOI22D1BWP30P140LVT U106 ( .A1(n178), .A2(i_data_bus[232]), .B1(n1), .B2(
        i_data_bus[72]), .ZN(n81) );
  ND4D1BWP30P140LVT U107 ( .A1(n84), .A2(n83), .A3(n82), .A4(n81), .ZN(N377)
         );
  AOI22D1BWP30P140LVT U108 ( .A1(n173), .A2(i_data_bus[133]), .B1(n93), .B2(
        i_data_bus[5]), .ZN(n88) );
  AOI22D1BWP30P140LVT U109 ( .A1(n175), .A2(i_data_bus[37]), .B1(n174), .B2(
        i_data_bus[101]), .ZN(n87) );
  AOI22D1BWP30P140LVT U110 ( .A1(n177), .A2(i_data_bus[197]), .B1(n94), .B2(
        i_data_bus[165]), .ZN(n86) );
  AOI22D1BWP30P140LVT U111 ( .A1(n178), .A2(i_data_bus[229]), .B1(n1), .B2(
        i_data_bus[69]), .ZN(n85) );
  ND4D1BWP30P140LVT U112 ( .A1(n88), .A2(n87), .A3(n86), .A4(n85), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U113 ( .A1(n173), .A2(i_data_bus[130]), .B1(n93), .B2(
        i_data_bus[2]), .ZN(n92) );
  AOI22D1BWP30P140LVT U114 ( .A1(n175), .A2(i_data_bus[34]), .B1(n174), .B2(
        i_data_bus[98]), .ZN(n91) );
  AOI22D1BWP30P140LVT U115 ( .A1(n177), .A2(i_data_bus[194]), .B1(n94), .B2(
        i_data_bus[162]), .ZN(n90) );
  AOI22D1BWP30P140LVT U116 ( .A1(n178), .A2(i_data_bus[226]), .B1(n1), .B2(
        i_data_bus[66]), .ZN(n89) );
  ND4D1BWP30P140LVT U117 ( .A1(n92), .A2(n91), .A3(n90), .A4(n89), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U118 ( .A1(n173), .A2(i_data_bus[129]), .B1(n93), .B2(
        i_data_bus[1]), .ZN(n98) );
  AOI22D1BWP30P140LVT U119 ( .A1(n175), .A2(i_data_bus[33]), .B1(n174), .B2(
        i_data_bus[97]), .ZN(n97) );
  AOI22D1BWP30P140LVT U120 ( .A1(n177), .A2(i_data_bus[193]), .B1(n94), .B2(
        i_data_bus[161]), .ZN(n96) );
  AOI22D1BWP30P140LVT U121 ( .A1(n178), .A2(i_data_bus[225]), .B1(n1), .B2(
        i_data_bus[65]), .ZN(n95) );
  ND4D1BWP30P140LVT U122 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .ZN(N370)
         );
  AOI22D1BWP30P140LVT U123 ( .A1(n173), .A2(i_data_bus[143]), .B1(n172), .B2(
        i_data_bus[15]), .ZN(n102) );
  AOI22D1BWP30P140LVT U124 ( .A1(n175), .A2(i_data_bus[47]), .B1(n174), .B2(
        i_data_bus[111]), .ZN(n101) );
  AOI22D1BWP30P140LVT U125 ( .A1(n177), .A2(i_data_bus[207]), .B1(n176), .B2(
        i_data_bus[175]), .ZN(n100) );
  AOI22D1BWP30P140LVT U126 ( .A1(n178), .A2(i_data_bus[239]), .B1(n1), .B2(
        i_data_bus[79]), .ZN(n99) );
  ND4D1BWP30P140LVT U127 ( .A1(n102), .A2(n101), .A3(n100), .A4(n99), .ZN(N384) );
  AOI22D1BWP30P140LVT U128 ( .A1(n173), .A2(i_data_bus[142]), .B1(n172), .B2(
        i_data_bus[14]), .ZN(n106) );
  AOI22D1BWP30P140LVT U129 ( .A1(n175), .A2(i_data_bus[46]), .B1(n174), .B2(
        i_data_bus[110]), .ZN(n105) );
  AOI22D1BWP30P140LVT U130 ( .A1(n177), .A2(i_data_bus[206]), .B1(n176), .B2(
        i_data_bus[174]), .ZN(n104) );
  AOI22D1BWP30P140LVT U131 ( .A1(n178), .A2(i_data_bus[238]), .B1(n1), .B2(
        i_data_bus[78]), .ZN(n103) );
  ND4D1BWP30P140LVT U132 ( .A1(n106), .A2(n105), .A3(n104), .A4(n103), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U133 ( .A1(n173), .A2(i_data_bus[141]), .B1(n172), .B2(
        i_data_bus[13]), .ZN(n110) );
  AOI22D1BWP30P140LVT U134 ( .A1(n175), .A2(i_data_bus[45]), .B1(n174), .B2(
        i_data_bus[109]), .ZN(n109) );
  AOI22D1BWP30P140LVT U135 ( .A1(n177), .A2(i_data_bus[205]), .B1(n176), .B2(
        i_data_bus[173]), .ZN(n108) );
  AOI22D1BWP30P140LVT U136 ( .A1(n178), .A2(i_data_bus[237]), .B1(n1), .B2(
        i_data_bus[77]), .ZN(n107) );
  ND4D1BWP30P140LVT U137 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .ZN(
        N382) );
  AOI22D1BWP30P140LVT U138 ( .A1(n173), .A2(i_data_bus[159]), .B1(n172), .B2(
        i_data_bus[31]), .ZN(n114) );
  AOI22D1BWP30P140LVT U139 ( .A1(n175), .A2(i_data_bus[63]), .B1(n174), .B2(
        i_data_bus[127]), .ZN(n113) );
  AOI22D1BWP30P140LVT U140 ( .A1(n167), .A2(i_data_bus[223]), .B1(n176), .B2(
        i_data_bus[191]), .ZN(n112) );
  AOI22D1BWP30P140LVT U141 ( .A1(n178), .A2(i_data_bus[255]), .B1(n1), .B2(
        i_data_bus[95]), .ZN(n111) );
  ND4D1BWP30P140LVT U142 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U143 ( .A1(n173), .A2(i_data_bus[158]), .B1(n172), .B2(
        i_data_bus[30]), .ZN(n118) );
  AOI22D1BWP30P140LVT U144 ( .A1(n175), .A2(i_data_bus[62]), .B1(n174), .B2(
        i_data_bus[126]), .ZN(n117) );
  AOI22D1BWP30P140LVT U145 ( .A1(n167), .A2(i_data_bus[222]), .B1(n176), .B2(
        i_data_bus[190]), .ZN(n116) );
  AOI22D1BWP30P140LVT U146 ( .A1(n178), .A2(i_data_bus[254]), .B1(n1), .B2(
        i_data_bus[94]), .ZN(n115) );
  ND4D1BWP30P140LVT U147 ( .A1(n118), .A2(n117), .A3(n116), .A4(n115), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U148 ( .A1(n173), .A2(i_data_bus[157]), .B1(n172), .B2(
        i_data_bus[29]), .ZN(n122) );
  AOI22D1BWP30P140LVT U149 ( .A1(n175), .A2(i_data_bus[61]), .B1(n174), .B2(
        i_data_bus[125]), .ZN(n121) );
  AOI22D1BWP30P140LVT U150 ( .A1(n167), .A2(i_data_bus[221]), .B1(n176), .B2(
        i_data_bus[189]), .ZN(n120) );
  AOI22D1BWP30P140LVT U151 ( .A1(n178), .A2(i_data_bus[253]), .B1(n1), .B2(
        i_data_bus[93]), .ZN(n119) );
  ND4D1BWP30P140LVT U152 ( .A1(n122), .A2(n121), .A3(n120), .A4(n119), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U153 ( .A1(n173), .A2(i_data_bus[156]), .B1(n172), .B2(
        i_data_bus[28]), .ZN(n126) );
  AOI22D1BWP30P140LVT U154 ( .A1(n175), .A2(i_data_bus[60]), .B1(n174), .B2(
        i_data_bus[124]), .ZN(n125) );
  AOI22D1BWP30P140LVT U155 ( .A1(n167), .A2(i_data_bus[220]), .B1(n176), .B2(
        i_data_bus[188]), .ZN(n124) );
  AOI22D1BWP30P140LVT U156 ( .A1(n178), .A2(i_data_bus[252]), .B1(n1), .B2(
        i_data_bus[92]), .ZN(n123) );
  ND4D1BWP30P140LVT U157 ( .A1(n126), .A2(n125), .A3(n124), .A4(n123), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U158 ( .A1(n173), .A2(i_data_bus[155]), .B1(n172), .B2(
        i_data_bus[27]), .ZN(n130) );
  AOI22D1BWP30P140LVT U159 ( .A1(n175), .A2(i_data_bus[59]), .B1(n174), .B2(
        i_data_bus[123]), .ZN(n129) );
  AOI22D1BWP30P140LVT U160 ( .A1(n167), .A2(i_data_bus[219]), .B1(n176), .B2(
        i_data_bus[187]), .ZN(n128) );
  AOI22D1BWP30P140LVT U161 ( .A1(n178), .A2(i_data_bus[251]), .B1(n1), .B2(
        i_data_bus[91]), .ZN(n127) );
  ND4D1BWP30P140LVT U162 ( .A1(n130), .A2(n129), .A3(n128), .A4(n127), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U163 ( .A1(n173), .A2(i_data_bus[154]), .B1(n172), .B2(
        i_data_bus[26]), .ZN(n134) );
  AOI22D1BWP30P140LVT U164 ( .A1(n175), .A2(i_data_bus[58]), .B1(n174), .B2(
        i_data_bus[122]), .ZN(n133) );
  AOI22D1BWP30P140LVT U165 ( .A1(n167), .A2(i_data_bus[218]), .B1(n176), .B2(
        i_data_bus[186]), .ZN(n132) );
  AOI22D1BWP30P140LVT U166 ( .A1(n178), .A2(i_data_bus[250]), .B1(n1), .B2(
        i_data_bus[90]), .ZN(n131) );
  ND4D1BWP30P140LVT U167 ( .A1(n134), .A2(n133), .A3(n132), .A4(n131), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U168 ( .A1(n173), .A2(i_data_bus[153]), .B1(n172), .B2(
        i_data_bus[25]), .ZN(n138) );
  AOI22D1BWP30P140LVT U169 ( .A1(n175), .A2(i_data_bus[57]), .B1(n174), .B2(
        i_data_bus[121]), .ZN(n137) );
  AOI22D1BWP30P140LVT U170 ( .A1(n167), .A2(i_data_bus[217]), .B1(n176), .B2(
        i_data_bus[185]), .ZN(n136) );
  AOI22D1BWP30P140LVT U171 ( .A1(n178), .A2(i_data_bus[249]), .B1(n1), .B2(
        i_data_bus[89]), .ZN(n135) );
  ND4D1BWP30P140LVT U172 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U173 ( .A1(n173), .A2(i_data_bus[152]), .B1(n172), .B2(
        i_data_bus[24]), .ZN(n142) );
  AOI22D1BWP30P140LVT U174 ( .A1(n175), .A2(i_data_bus[56]), .B1(n174), .B2(
        i_data_bus[120]), .ZN(n141) );
  AOI22D1BWP30P140LVT U175 ( .A1(n167), .A2(i_data_bus[216]), .B1(n176), .B2(
        i_data_bus[184]), .ZN(n140) );
  AOI22D1BWP30P140LVT U176 ( .A1(n178), .A2(i_data_bus[248]), .B1(n1), .B2(
        i_data_bus[88]), .ZN(n139) );
  ND4D1BWP30P140LVT U177 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U178 ( .A1(n173), .A2(i_data_bus[151]), .B1(n172), .B2(
        i_data_bus[23]), .ZN(n146) );
  AOI22D1BWP30P140LVT U179 ( .A1(n175), .A2(i_data_bus[55]), .B1(n174), .B2(
        i_data_bus[119]), .ZN(n145) );
  AOI22D1BWP30P140LVT U180 ( .A1(n167), .A2(i_data_bus[215]), .B1(n176), .B2(
        i_data_bus[183]), .ZN(n144) );
  AOI22D1BWP30P140LVT U181 ( .A1(n178), .A2(i_data_bus[247]), .B1(n1), .B2(
        i_data_bus[87]), .ZN(n143) );
  ND4D1BWP30P140LVT U182 ( .A1(n146), .A2(n145), .A3(n144), .A4(n143), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U183 ( .A1(n173), .A2(i_data_bus[150]), .B1(n172), .B2(
        i_data_bus[22]), .ZN(n150) );
  AOI22D1BWP30P140LVT U184 ( .A1(n175), .A2(i_data_bus[54]), .B1(n174), .B2(
        i_data_bus[118]), .ZN(n149) );
  AOI22D1BWP30P140LVT U185 ( .A1(n167), .A2(i_data_bus[214]), .B1(n176), .B2(
        i_data_bus[182]), .ZN(n148) );
  AOI22D1BWP30P140LVT U186 ( .A1(n178), .A2(i_data_bus[246]), .B1(n1), .B2(
        i_data_bus[86]), .ZN(n147) );
  ND4D1BWP30P140LVT U187 ( .A1(n150), .A2(n149), .A3(n148), .A4(n147), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U188 ( .A1(n173), .A2(i_data_bus[149]), .B1(n172), .B2(
        i_data_bus[21]), .ZN(n154) );
  AOI22D1BWP30P140LVT U189 ( .A1(n175), .A2(i_data_bus[53]), .B1(n174), .B2(
        i_data_bus[117]), .ZN(n153) );
  AOI22D1BWP30P140LVT U190 ( .A1(n167), .A2(i_data_bus[213]), .B1(n176), .B2(
        i_data_bus[181]), .ZN(n152) );
  AOI22D1BWP30P140LVT U191 ( .A1(n178), .A2(i_data_bus[245]), .B1(n1), .B2(
        i_data_bus[85]), .ZN(n151) );
  ND4D1BWP30P140LVT U192 ( .A1(n154), .A2(n153), .A3(n152), .A4(n151), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U193 ( .A1(n173), .A2(i_data_bus[148]), .B1(n172), .B2(
        i_data_bus[20]), .ZN(n158) );
  AOI22D1BWP30P140LVT U194 ( .A1(n175), .A2(i_data_bus[52]), .B1(n174), .B2(
        i_data_bus[116]), .ZN(n157) );
  AOI22D1BWP30P140LVT U195 ( .A1(n167), .A2(i_data_bus[212]), .B1(n176), .B2(
        i_data_bus[180]), .ZN(n156) );
  AOI22D1BWP30P140LVT U196 ( .A1(n178), .A2(i_data_bus[244]), .B1(n1), .B2(
        i_data_bus[84]), .ZN(n155) );
  ND4D1BWP30P140LVT U197 ( .A1(n158), .A2(n157), .A3(n156), .A4(n155), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U198 ( .A1(n173), .A2(i_data_bus[147]), .B1(n172), .B2(
        i_data_bus[19]), .ZN(n162) );
  AOI22D1BWP30P140LVT U199 ( .A1(n175), .A2(i_data_bus[51]), .B1(n174), .B2(
        i_data_bus[115]), .ZN(n161) );
  AOI22D1BWP30P140LVT U200 ( .A1(n167), .A2(i_data_bus[211]), .B1(n176), .B2(
        i_data_bus[179]), .ZN(n160) );
  AOI22D1BWP30P140LVT U201 ( .A1(n178), .A2(i_data_bus[243]), .B1(n1), .B2(
        i_data_bus[83]), .ZN(n159) );
  ND4D1BWP30P140LVT U202 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U203 ( .A1(n173), .A2(i_data_bus[146]), .B1(n172), .B2(
        i_data_bus[18]), .ZN(n166) );
  AOI22D1BWP30P140LVT U204 ( .A1(n175), .A2(i_data_bus[50]), .B1(n174), .B2(
        i_data_bus[114]), .ZN(n165) );
  AOI22D1BWP30P140LVT U205 ( .A1(n167), .A2(i_data_bus[210]), .B1(n176), .B2(
        i_data_bus[178]), .ZN(n164) );
  AOI22D1BWP30P140LVT U206 ( .A1(n178), .A2(i_data_bus[242]), .B1(n1), .B2(
        i_data_bus[82]), .ZN(n163) );
  ND4D1BWP30P140LVT U207 ( .A1(n166), .A2(n165), .A3(n164), .A4(n163), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U208 ( .A1(n173), .A2(i_data_bus[145]), .B1(n172), .B2(
        i_data_bus[17]), .ZN(n171) );
  AOI22D1BWP30P140LVT U209 ( .A1(n175), .A2(i_data_bus[49]), .B1(n174), .B2(
        i_data_bus[113]), .ZN(n170) );
  AOI22D1BWP30P140LVT U210 ( .A1(n167), .A2(i_data_bus[209]), .B1(n176), .B2(
        i_data_bus[177]), .ZN(n169) );
  AOI22D1BWP30P140LVT U211 ( .A1(n178), .A2(i_data_bus[241]), .B1(n1), .B2(
        i_data_bus[81]), .ZN(n168) );
  ND4D1BWP30P140LVT U212 ( .A1(n171), .A2(n170), .A3(n169), .A4(n168), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U213 ( .A1(n173), .A2(i_data_bus[144]), .B1(n172), .B2(
        i_data_bus[16]), .ZN(n182) );
  AOI22D1BWP30P140LVT U214 ( .A1(n175), .A2(i_data_bus[48]), .B1(n174), .B2(
        i_data_bus[112]), .ZN(n181) );
  AOI22D1BWP30P140LVT U215 ( .A1(n177), .A2(i_data_bus[208]), .B1(n176), .B2(
        i_data_bus[176]), .ZN(n180) );
  AOI22D1BWP30P140LVT U216 ( .A1(n178), .A2(i_data_bus[240]), .B1(n1), .B2(
        i_data_bus[80]), .ZN(n179) );
  ND4D1BWP30P140LVT U217 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(
        N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_2 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n24), .Z(n178) );
  INVD3BWP30P140LVT U4 ( .I(n12), .ZN(n173) );
  INVD1BWP30P140LVT U5 ( .I(n11), .ZN(n12) );
  NR2D1BWP30P140LVT U6 ( .A1(i_cmd[2]), .A2(i_cmd[1]), .ZN(n20) );
  CKND2D2BWP30P140LVT U7 ( .A1(n3), .A2(n2), .ZN(n10) );
  INVD1BWP30P140LVT U8 ( .I(i_cmd[3]), .ZN(n18) );
  INVD1BWP30P140LVT U9 ( .I(i_cmd[7]), .ZN(n2) );
  INR2D2BWP30P140LVT U10 ( .A1(n17), .B1(i_cmd[5]), .ZN(n3) );
  IND3D4BWP30P140LVT U11 ( .A1(n10), .B1(n9), .B2(n8), .ZN(n14) );
  BUFFD4BWP30P140LVT U12 ( .I(n36), .Z(n1) );
  INVD1BWP30P140LVT U13 ( .I(n27), .ZN(n73) );
  NR4D0BWP30P140LVT U14 ( .A1(n35), .A2(i_cmd[5]), .A3(n26), .A4(n25), .ZN(n27) );
  INVD1BWP30P140LVT U15 ( .I(i_cmd[6]), .ZN(n25) );
  INVD1BWP30P140LVT U16 ( .I(i_cmd[2]), .ZN(n30) );
  NR2D1BWP30P140LVT U17 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n9) );
  NR2D1BWP30P140LVT U18 ( .A1(i_cmd[6]), .A2(i_cmd[1]), .ZN(n8) );
  INR2D4BWP30P140LVT U19 ( .A1(n28), .B1(n7), .ZN(n174) );
  ND2D1BWP30P140LVT U20 ( .A1(n20), .A2(n6), .ZN(n7) );
  NR2D1BWP30P140LVT U21 ( .A1(n18), .A2(n5), .ZN(n6) );
  NR4D1BWP30P140LVT U22 ( .A1(n35), .A2(i_cmd[6]), .A3(n34), .A4(n33), .ZN(n36) );
  NR2D1BWP30P140LVT U23 ( .A1(n35), .A2(n23), .ZN(n24) );
  NR2D1BWP30P140LVT U24 ( .A1(i_cmd[6]), .A2(i_cmd[5]), .ZN(n22) );
  ND2D1BWP30P140LVT U25 ( .A1(n38), .A2(n37), .ZN(N402) );
  INVD1BWP30P140LVT U26 ( .I(i_cmd[4]), .ZN(n13) );
  INR2D1BWP30P140LVT U27 ( .A1(i_en), .B1(rst), .ZN(n17) );
  NR4D3BWP30P140LVT U28 ( .A1(n10), .A2(i_cmd[0]), .A3(i_cmd[6]), .A4(i_cmd[4]), .ZN(n28) );
  ND3D1BWP30P140LVT U29 ( .A1(n9), .A2(i_valid[1]), .A3(i_cmd[1]), .ZN(n4) );
  INR2D4BWP30P140LVT U30 ( .A1(n28), .B1(n4), .ZN(n175) );
  INVD1BWP30P140LVT U31 ( .I(i_valid[3]), .ZN(n5) );
  INR4D1BWP30P140LVT U32 ( .A1(i_valid[4]), .B1(i_cmd[0]), .B2(n13), .B3(n14), 
        .ZN(n11) );
  INVD1BWP30P140LVT U33 ( .I(i_cmd[0]), .ZN(n15) );
  INR4D1BWP30P140LVT U34 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n15), .B3(n14), 
        .ZN(n16) );
  INVD2BWP30P140LVT U35 ( .I(n16), .ZN(n87) );
  INVD6BWP30P140LVT U36 ( .I(n87), .ZN(n172) );
  NR4D0BWP30P140LVT U37 ( .A1(n175), .A2(n174), .A3(n173), .A4(n172), .ZN(n38)
         );
  NR2OPTPAD1BWP30P140LVT U38 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n21) );
  CKAN2D1BWP30P140LVT U39 ( .A1(n18), .A2(n17), .Z(n19) );
  ND3OPTPAD2BWP30P140LVT U40 ( .A1(n21), .A2(n20), .A3(n19), .ZN(n35) );
  ND3D1BWP30P140LVT U41 ( .A1(n22), .A2(i_valid[7]), .A3(i_cmd[7]), .ZN(n23)
         );
  IND2D1BWP30P140LVT U42 ( .A1(i_cmd[7]), .B1(i_valid[6]), .ZN(n26) );
  INVD2BWP30P140LVT U43 ( .I(n73), .ZN(n167) );
  INVD2BWP30P140LVT U44 ( .I(n28), .ZN(n31) );
  IND2D1BWP30P140LVT U45 ( .A1(i_cmd[3]), .B1(i_valid[2]), .ZN(n29) );
  NR4D1BWP30P140LVT U46 ( .A1(n31), .A2(i_cmd[1]), .A3(n30), .A4(n29), .ZN(n32) );
  INVD2BWP30P140LVT U47 ( .I(n32), .ZN(n93) );
  INVD2BWP30P140LVT U48 ( .I(n93), .ZN(n177) );
  INVD1BWP30P140LVT U49 ( .I(i_cmd[5]), .ZN(n34) );
  IND2D1BWP30P140LVT U50 ( .A1(i_cmd[7]), .B1(i_valid[5]), .ZN(n33) );
  NR4D0BWP30P140LVT U51 ( .A1(n178), .A2(n167), .A3(n177), .A4(n1), .ZN(n37)
         );
  AOI22D1BWP30P140LVT U52 ( .A1(n173), .A2(i_data_bus[140]), .B1(n172), .B2(
        i_data_bus[12]), .ZN(n42) );
  AOI22D1BWP30P140LVT U53 ( .A1(n175), .A2(i_data_bus[44]), .B1(n174), .B2(
        i_data_bus[108]), .ZN(n41) );
  INVD2BWP30P140LVT U54 ( .I(n73), .ZN(n176) );
  AOI22D1BWP30P140LVT U55 ( .A1(n176), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n40) );
  INVD2BWP30P140LVT U56 ( .I(n93), .ZN(n158) );
  AOI22D1BWP30P140LVT U57 ( .A1(n178), .A2(i_data_bus[236]), .B1(n158), .B2(
        i_data_bus[76]), .ZN(n39) );
  ND4D1BWP30P140LVT U58 ( .A1(n42), .A2(n41), .A3(n40), .A4(n39), .ZN(N381) );
  AOI22D1BWP30P140LVT U59 ( .A1(n173), .A2(i_data_bus[138]), .B1(n172), .B2(
        i_data_bus[10]), .ZN(n46) );
  AOI22D1BWP30P140LVT U60 ( .A1(n175), .A2(i_data_bus[42]), .B1(n174), .B2(
        i_data_bus[106]), .ZN(n45) );
  AOI22D1BWP30P140LVT U61 ( .A1(n176), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n44) );
  AOI22D1BWP30P140LVT U62 ( .A1(n178), .A2(i_data_bus[234]), .B1(n158), .B2(
        i_data_bus[74]), .ZN(n43) );
  ND4D1BWP30P140LVT U63 ( .A1(n46), .A2(n45), .A3(n44), .A4(n43), .ZN(N379) );
  AOI22D1BWP30P140LVT U64 ( .A1(n173), .A2(i_data_bus[137]), .B1(n172), .B2(
        i_data_bus[9]), .ZN(n50) );
  AOI22D1BWP30P140LVT U65 ( .A1(n175), .A2(i_data_bus[41]), .B1(n174), .B2(
        i_data_bus[105]), .ZN(n49) );
  AOI22D1BWP30P140LVT U66 ( .A1(n176), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n48) );
  AOI22D1BWP30P140LVT U67 ( .A1(n178), .A2(i_data_bus[233]), .B1(n158), .B2(
        i_data_bus[73]), .ZN(n47) );
  ND4D1BWP30P140LVT U68 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(N378) );
  AOI22D1BWP30P140LVT U69 ( .A1(n173), .A2(i_data_bus[135]), .B1(n172), .B2(
        i_data_bus[7]), .ZN(n54) );
  AOI22D1BWP30P140LVT U70 ( .A1(n175), .A2(i_data_bus[39]), .B1(n174), .B2(
        i_data_bus[103]), .ZN(n53) );
  AOI22D1BWP30P140LVT U71 ( .A1(n176), .A2(i_data_bus[199]), .B1(n1), .B2(
        i_data_bus[167]), .ZN(n52) );
  AOI22D1BWP30P140LVT U72 ( .A1(n178), .A2(i_data_bus[231]), .B1(n158), .B2(
        i_data_bus[71]), .ZN(n51) );
  ND4D1BWP30P140LVT U73 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(N376) );
  INVD1BWP30P140LVT U74 ( .I(i_data_bus[6]), .ZN(n55) );
  MAOI22D1BWP30P140LVT U75 ( .A1(n173), .A2(i_data_bus[134]), .B1(n87), .B2(
        n55), .ZN(n59) );
  AOI22D1BWP30P140LVT U76 ( .A1(n175), .A2(i_data_bus[38]), .B1(n174), .B2(
        i_data_bus[102]), .ZN(n58) );
  AOI22D1BWP30P140LVT U77 ( .A1(n176), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n57) );
  AOI22D1BWP30P140LVT U78 ( .A1(n178), .A2(i_data_bus[230]), .B1(n158), .B2(
        i_data_bus[70]), .ZN(n56) );
  ND4D1BWP30P140LVT U79 ( .A1(n59), .A2(n58), .A3(n57), .A4(n56), .ZN(N375) );
  AOI22D1BWP30P140LVT U80 ( .A1(n173), .A2(i_data_bus[132]), .B1(n172), .B2(
        i_data_bus[4]), .ZN(n63) );
  AOI22D1BWP30P140LVT U81 ( .A1(n175), .A2(i_data_bus[36]), .B1(n174), .B2(
        i_data_bus[100]), .ZN(n62) );
  AOI22D1BWP30P140LVT U82 ( .A1(n176), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n61) );
  AOI22D1BWP30P140LVT U83 ( .A1(n178), .A2(i_data_bus[228]), .B1(n158), .B2(
        i_data_bus[68]), .ZN(n60) );
  ND4D1BWP30P140LVT U84 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(N373) );
  AOI22D1BWP30P140LVT U85 ( .A1(n173), .A2(i_data_bus[131]), .B1(n172), .B2(
        i_data_bus[3]), .ZN(n67) );
  AOI22D1BWP30P140LVT U86 ( .A1(n175), .A2(i_data_bus[35]), .B1(n174), .B2(
        i_data_bus[99]), .ZN(n66) );
  AOI22D1BWP30P140LVT U87 ( .A1(n176), .A2(i_data_bus[195]), .B1(n1), .B2(
        i_data_bus[163]), .ZN(n65) );
  AOI22D1BWP30P140LVT U88 ( .A1(n178), .A2(i_data_bus[227]), .B1(n158), .B2(
        i_data_bus[67]), .ZN(n64) );
  ND4D1BWP30P140LVT U89 ( .A1(n67), .A2(n66), .A3(n65), .A4(n64), .ZN(N372) );
  AOI22D1BWP30P140LVT U90 ( .A1(n173), .A2(i_data_bus[129]), .B1(n172), .B2(
        i_data_bus[1]), .ZN(n71) );
  AOI22D1BWP30P140LVT U91 ( .A1(n175), .A2(i_data_bus[33]), .B1(n174), .B2(
        i_data_bus[97]), .ZN(n70) );
  AOI22D1BWP30P140LVT U92 ( .A1(n176), .A2(i_data_bus[193]), .B1(n1), .B2(
        i_data_bus[161]), .ZN(n69) );
  AOI22D1BWP30P140LVT U93 ( .A1(n178), .A2(i_data_bus[225]), .B1(n158), .B2(
        i_data_bus[65]), .ZN(n68) );
  ND4D1BWP30P140LVT U94 ( .A1(n71), .A2(n70), .A3(n69), .A4(n68), .ZN(N370) );
  INVD1BWP30P140LVT U95 ( .I(i_data_bus[0]), .ZN(n72) );
  MAOI22D1BWP30P140LVT U96 ( .A1(n173), .A2(i_data_bus[128]), .B1(n87), .B2(
        n72), .ZN(n77) );
  AOI22D1BWP30P140LVT U97 ( .A1(n175), .A2(i_data_bus[32]), .B1(n174), .B2(
        i_data_bus[96]), .ZN(n76) );
  AOI22D1BWP30P140LVT U98 ( .A1(n167), .A2(i_data_bus[192]), .B1(n1), .B2(
        i_data_bus[160]), .ZN(n75) );
  AOI22D1BWP30P140LVT U99 ( .A1(n178), .A2(i_data_bus[224]), .B1(n158), .B2(
        i_data_bus[64]), .ZN(n74) );
  ND4D1BWP30P140LVT U100 ( .A1(n77), .A2(n76), .A3(n75), .A4(n74), .ZN(N369)
         );
  AOI22D1BWP30P140LVT U101 ( .A1(n173), .A2(i_data_bus[139]), .B1(n172), .B2(
        i_data_bus[11]), .ZN(n81) );
  AOI22D1BWP30P140LVT U102 ( .A1(n175), .A2(i_data_bus[43]), .B1(n174), .B2(
        i_data_bus[107]), .ZN(n80) );
  AOI22D1BWP30P140LVT U103 ( .A1(n176), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n79) );
  AOI22D1BWP30P140LVT U104 ( .A1(n178), .A2(i_data_bus[235]), .B1(n158), .B2(
        i_data_bus[75]), .ZN(n78) );
  ND4D1BWP30P140LVT U105 ( .A1(n81), .A2(n80), .A3(n79), .A4(n78), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U106 ( .A1(n173), .A2(i_data_bus[136]), .B1(n172), .B2(
        i_data_bus[8]), .ZN(n85) );
  AOI22D1BWP30P140LVT U107 ( .A1(n175), .A2(i_data_bus[40]), .B1(n174), .B2(
        i_data_bus[104]), .ZN(n84) );
  AOI22D1BWP30P140LVT U108 ( .A1(n176), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n83) );
  AOI22D1BWP30P140LVT U109 ( .A1(n178), .A2(i_data_bus[232]), .B1(n158), .B2(
        i_data_bus[72]), .ZN(n82) );
  ND4D1BWP30P140LVT U110 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(N377)
         );
  INVD1BWP30P140LVT U111 ( .I(i_data_bus[5]), .ZN(n86) );
  MAOI22D1BWP30P140LVT U112 ( .A1(n173), .A2(i_data_bus[133]), .B1(n87), .B2(
        n86), .ZN(n91) );
  AOI22D1BWP30P140LVT U113 ( .A1(n175), .A2(i_data_bus[37]), .B1(n174), .B2(
        i_data_bus[101]), .ZN(n90) );
  AOI22D1BWP30P140LVT U114 ( .A1(n176), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n89) );
  AOI22D1BWP30P140LVT U115 ( .A1(n178), .A2(i_data_bus[229]), .B1(n158), .B2(
        i_data_bus[69]), .ZN(n88) );
  ND4D1BWP30P140LVT U116 ( .A1(n91), .A2(n90), .A3(n89), .A4(n88), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U117 ( .A1(n173), .A2(i_data_bus[130]), .B1(n172), .B2(
        i_data_bus[2]), .ZN(n97) );
  AOI22D1BWP30P140LVT U118 ( .A1(n175), .A2(i_data_bus[34]), .B1(n174), .B2(
        i_data_bus[98]), .ZN(n96) );
  AOI22D1BWP30P140LVT U119 ( .A1(n176), .A2(i_data_bus[194]), .B1(n1), .B2(
        i_data_bus[162]), .ZN(n95) );
  INVD1BWP30P140LVT U120 ( .I(i_data_bus[66]), .ZN(n92) );
  MAOI22D1BWP30P140LVT U121 ( .A1(n178), .A2(i_data_bus[226]), .B1(n93), .B2(
        n92), .ZN(n94) );
  ND4D1BWP30P140LVT U122 ( .A1(n97), .A2(n96), .A3(n95), .A4(n94), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U123 ( .A1(n173), .A2(i_data_bus[159]), .B1(n172), .B2(
        i_data_bus[31]), .ZN(n101) );
  AOI22D1BWP30P140LVT U124 ( .A1(n175), .A2(i_data_bus[63]), .B1(n174), .B2(
        i_data_bus[127]), .ZN(n100) );
  AOI22D1BWP30P140LVT U125 ( .A1(n167), .A2(i_data_bus[223]), .B1(n1), .B2(
        i_data_bus[191]), .ZN(n99) );
  AOI22D1BWP30P140LVT U126 ( .A1(n178), .A2(i_data_bus[255]), .B1(n177), .B2(
        i_data_bus[95]), .ZN(n98) );
  ND4D1BWP30P140LVT U127 ( .A1(n101), .A2(n100), .A3(n99), .A4(n98), .ZN(N400)
         );
  AOI22D1BWP30P140LVT U128 ( .A1(n173), .A2(i_data_bus[158]), .B1(n172), .B2(
        i_data_bus[30]), .ZN(n105) );
  AOI22D1BWP30P140LVT U129 ( .A1(n175), .A2(i_data_bus[62]), .B1(n174), .B2(
        i_data_bus[126]), .ZN(n104) );
  AOI22D1BWP30P140LVT U130 ( .A1(n167), .A2(i_data_bus[222]), .B1(n1), .B2(
        i_data_bus[190]), .ZN(n103) );
  AOI22D1BWP30P140LVT U131 ( .A1(n178), .A2(i_data_bus[254]), .B1(n177), .B2(
        i_data_bus[94]), .ZN(n102) );
  ND4D1BWP30P140LVT U132 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U133 ( .A1(n173), .A2(i_data_bus[156]), .B1(n172), .B2(
        i_data_bus[28]), .ZN(n109) );
  AOI22D1BWP30P140LVT U134 ( .A1(n175), .A2(i_data_bus[60]), .B1(n174), .B2(
        i_data_bus[124]), .ZN(n108) );
  AOI22D1BWP30P140LVT U135 ( .A1(n167), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n107) );
  AOI22D1BWP30P140LVT U136 ( .A1(n178), .A2(i_data_bus[252]), .B1(n177), .B2(
        i_data_bus[92]), .ZN(n106) );
  ND4D1BWP30P140LVT U137 ( .A1(n109), .A2(n108), .A3(n107), .A4(n106), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U138 ( .A1(n173), .A2(i_data_bus[155]), .B1(n172), .B2(
        i_data_bus[27]), .ZN(n113) );
  AOI22D1BWP30P140LVT U139 ( .A1(n175), .A2(i_data_bus[59]), .B1(n174), .B2(
        i_data_bus[123]), .ZN(n112) );
  AOI22D1BWP30P140LVT U140 ( .A1(n167), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n111) );
  AOI22D1BWP30P140LVT U141 ( .A1(n178), .A2(i_data_bus[251]), .B1(n177), .B2(
        i_data_bus[91]), .ZN(n110) );
  ND4D1BWP30P140LVT U142 ( .A1(n113), .A2(n112), .A3(n111), .A4(n110), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U143 ( .A1(n173), .A2(i_data_bus[153]), .B1(n172), .B2(
        i_data_bus[25]), .ZN(n117) );
  AOI22D1BWP30P140LVT U144 ( .A1(n175), .A2(i_data_bus[57]), .B1(n174), .B2(
        i_data_bus[121]), .ZN(n116) );
  AOI22D1BWP30P140LVT U145 ( .A1(n167), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n115) );
  AOI22D1BWP30P140LVT U146 ( .A1(n178), .A2(i_data_bus[249]), .B1(n177), .B2(
        i_data_bus[89]), .ZN(n114) );
  ND4D1BWP30P140LVT U147 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U148 ( .A1(n173), .A2(i_data_bus[152]), .B1(n172), .B2(
        i_data_bus[24]), .ZN(n121) );
  AOI22D1BWP30P140LVT U149 ( .A1(n175), .A2(i_data_bus[56]), .B1(n174), .B2(
        i_data_bus[120]), .ZN(n120) );
  AOI22D1BWP30P140LVT U150 ( .A1(n167), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n119) );
  AOI22D1BWP30P140LVT U151 ( .A1(n178), .A2(i_data_bus[248]), .B1(n177), .B2(
        i_data_bus[88]), .ZN(n118) );
  ND4D1BWP30P140LVT U152 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U153 ( .A1(n173), .A2(i_data_bus[150]), .B1(n172), .B2(
        i_data_bus[22]), .ZN(n125) );
  AOI22D1BWP30P140LVT U154 ( .A1(n175), .A2(i_data_bus[54]), .B1(n174), .B2(
        i_data_bus[118]), .ZN(n124) );
  AOI22D1BWP30P140LVT U155 ( .A1(n167), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n123) );
  AOI22D1BWP30P140LVT U156 ( .A1(n178), .A2(i_data_bus[246]), .B1(n177), .B2(
        i_data_bus[86]), .ZN(n122) );
  ND4D1BWP30P140LVT U157 ( .A1(n125), .A2(n124), .A3(n123), .A4(n122), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U158 ( .A1(n173), .A2(i_data_bus[149]), .B1(n172), .B2(
        i_data_bus[21]), .ZN(n129) );
  AOI22D1BWP30P140LVT U159 ( .A1(n175), .A2(i_data_bus[53]), .B1(n174), .B2(
        i_data_bus[117]), .ZN(n128) );
  AOI22D1BWP30P140LVT U160 ( .A1(n167), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n127) );
  AOI22D1BWP30P140LVT U161 ( .A1(n178), .A2(i_data_bus[245]), .B1(n177), .B2(
        i_data_bus[85]), .ZN(n126) );
  ND4D1BWP30P140LVT U162 ( .A1(n129), .A2(n128), .A3(n127), .A4(n126), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U163 ( .A1(n173), .A2(i_data_bus[147]), .B1(n172), .B2(
        i_data_bus[19]), .ZN(n133) );
  AOI22D1BWP30P140LVT U164 ( .A1(n175), .A2(i_data_bus[51]), .B1(n174), .B2(
        i_data_bus[115]), .ZN(n132) );
  AOI22D1BWP30P140LVT U165 ( .A1(n167), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n131) );
  AOI22D1BWP30P140LVT U166 ( .A1(n178), .A2(i_data_bus[243]), .B1(n177), .B2(
        i_data_bus[83]), .ZN(n130) );
  ND4D1BWP30P140LVT U167 ( .A1(n133), .A2(n132), .A3(n131), .A4(n130), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U168 ( .A1(n173), .A2(i_data_bus[143]), .B1(n172), .B2(
        i_data_bus[15]), .ZN(n137) );
  AOI22D1BWP30P140LVT U169 ( .A1(n175), .A2(i_data_bus[47]), .B1(n174), .B2(
        i_data_bus[111]), .ZN(n136) );
  AOI22D1BWP30P140LVT U170 ( .A1(n176), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n135) );
  AOI22D1BWP30P140LVT U171 ( .A1(n178), .A2(i_data_bus[239]), .B1(n158), .B2(
        i_data_bus[79]), .ZN(n134) );
  ND4D1BWP30P140LVT U172 ( .A1(n137), .A2(n136), .A3(n135), .A4(n134), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U173 ( .A1(n173), .A2(i_data_bus[141]), .B1(n172), .B2(
        i_data_bus[13]), .ZN(n141) );
  AOI22D1BWP30P140LVT U174 ( .A1(n175), .A2(i_data_bus[45]), .B1(n174), .B2(
        i_data_bus[109]), .ZN(n140) );
  AOI22D1BWP30P140LVT U175 ( .A1(n176), .A2(i_data_bus[205]), .B1(n1), .B2(
        i_data_bus[173]), .ZN(n139) );
  AOI22D1BWP30P140LVT U176 ( .A1(n178), .A2(i_data_bus[237]), .B1(n158), .B2(
        i_data_bus[77]), .ZN(n138) );
  ND4D1BWP30P140LVT U177 ( .A1(n141), .A2(n140), .A3(n139), .A4(n138), .ZN(
        N382) );
  AOI22D1BWP30P140LVT U178 ( .A1(n173), .A2(i_data_bus[157]), .B1(n172), .B2(
        i_data_bus[29]), .ZN(n145) );
  AOI22D1BWP30P140LVT U179 ( .A1(n175), .A2(i_data_bus[61]), .B1(n174), .B2(
        i_data_bus[125]), .ZN(n144) );
  AOI22D1BWP30P140LVT U180 ( .A1(n167), .A2(i_data_bus[221]), .B1(n1), .B2(
        i_data_bus[189]), .ZN(n143) );
  AOI22D1BWP30P140LVT U181 ( .A1(n178), .A2(i_data_bus[253]), .B1(n177), .B2(
        i_data_bus[93]), .ZN(n142) );
  ND4D1BWP30P140LVT U182 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U183 ( .A1(n173), .A2(i_data_bus[154]), .B1(n172), .B2(
        i_data_bus[26]), .ZN(n149) );
  AOI22D1BWP30P140LVT U184 ( .A1(n175), .A2(i_data_bus[58]), .B1(n174), .B2(
        i_data_bus[122]), .ZN(n148) );
  AOI22D1BWP30P140LVT U185 ( .A1(n167), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n147) );
  AOI22D1BWP30P140LVT U186 ( .A1(n178), .A2(i_data_bus[250]), .B1(n177), .B2(
        i_data_bus[90]), .ZN(n146) );
  ND4D1BWP30P140LVT U187 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U188 ( .A1(n173), .A2(i_data_bus[151]), .B1(n172), .B2(
        i_data_bus[23]), .ZN(n153) );
  AOI22D1BWP30P140LVT U189 ( .A1(n175), .A2(i_data_bus[55]), .B1(n174), .B2(
        i_data_bus[119]), .ZN(n152) );
  AOI22D1BWP30P140LVT U190 ( .A1(n167), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n151) );
  AOI22D1BWP30P140LVT U191 ( .A1(n178), .A2(i_data_bus[247]), .B1(n177), .B2(
        i_data_bus[87]), .ZN(n150) );
  ND4D1BWP30P140LVT U192 ( .A1(n153), .A2(n152), .A3(n151), .A4(n150), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U193 ( .A1(n173), .A2(i_data_bus[148]), .B1(n172), .B2(
        i_data_bus[20]), .ZN(n157) );
  AOI22D1BWP30P140LVT U194 ( .A1(n175), .A2(i_data_bus[52]), .B1(n174), .B2(
        i_data_bus[116]), .ZN(n156) );
  AOI22D1BWP30P140LVT U195 ( .A1(n167), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n155) );
  AOI22D1BWP30P140LVT U196 ( .A1(n178), .A2(i_data_bus[244]), .B1(n177), .B2(
        i_data_bus[84]), .ZN(n154) );
  ND4D1BWP30P140LVT U197 ( .A1(n157), .A2(n156), .A3(n155), .A4(n154), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U198 ( .A1(n173), .A2(i_data_bus[142]), .B1(n172), .B2(
        i_data_bus[14]), .ZN(n162) );
  AOI22D1BWP30P140LVT U199 ( .A1(n175), .A2(i_data_bus[46]), .B1(n174), .B2(
        i_data_bus[110]), .ZN(n161) );
  AOI22D1BWP30P140LVT U200 ( .A1(n176), .A2(i_data_bus[206]), .B1(n1), .B2(
        i_data_bus[174]), .ZN(n160) );
  AOI22D1BWP30P140LVT U201 ( .A1(n178), .A2(i_data_bus[238]), .B1(n158), .B2(
        i_data_bus[78]), .ZN(n159) );
  ND4D1BWP30P140LVT U202 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U203 ( .A1(n173), .A2(i_data_bus[146]), .B1(n172), .B2(
        i_data_bus[18]), .ZN(n166) );
  AOI22D1BWP30P140LVT U204 ( .A1(n175), .A2(i_data_bus[50]), .B1(n174), .B2(
        i_data_bus[114]), .ZN(n165) );
  AOI22D1BWP30P140LVT U205 ( .A1(n167), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n164) );
  AOI22D1BWP30P140LVT U206 ( .A1(n178), .A2(i_data_bus[242]), .B1(n177), .B2(
        i_data_bus[82]), .ZN(n163) );
  ND4D1BWP30P140LVT U207 ( .A1(n166), .A2(n165), .A3(n164), .A4(n163), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U208 ( .A1(n173), .A2(i_data_bus[145]), .B1(n172), .B2(
        i_data_bus[17]), .ZN(n171) );
  AOI22D1BWP30P140LVT U209 ( .A1(n175), .A2(i_data_bus[49]), .B1(n174), .B2(
        i_data_bus[113]), .ZN(n170) );
  AOI22D1BWP30P140LVT U210 ( .A1(n167), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n169) );
  AOI22D1BWP30P140LVT U211 ( .A1(n178), .A2(i_data_bus[241]), .B1(n177), .B2(
        i_data_bus[81]), .ZN(n168) );
  ND4D1BWP30P140LVT U212 ( .A1(n171), .A2(n170), .A3(n169), .A4(n168), .ZN(
        N386) );
  AOI22D1BWP30P140LVT U213 ( .A1(n173), .A2(i_data_bus[144]), .B1(n172), .B2(
        i_data_bus[16]), .ZN(n182) );
  AOI22D1BWP30P140LVT U214 ( .A1(n175), .A2(i_data_bus[48]), .B1(n174), .B2(
        i_data_bus[112]), .ZN(n181) );
  AOI22D1BWP30P140LVT U215 ( .A1(n176), .A2(i_data_bus[208]), .B1(n1), .B2(
        i_data_bus[176]), .ZN(n180) );
  AOI22D1BWP30P140LVT U216 ( .A1(n178), .A2(i_data_bus[240]), .B1(n177), .B2(
        i_data_bus[80]), .ZN(n179) );
  ND4D1BWP30P140LVT U217 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(
        N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_3 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD2BWP30P140LVT U3 ( .I(n39), .ZN(n42) );
  OR2D1BWP30P140LVT U4 ( .A1(n34), .A2(n5), .Z(n2) );
  NR4D1BWP30P140LVT U5 ( .A1(n38), .A2(i_cmd[6]), .A3(n37), .A4(n36), .ZN(n39)
         );
  IND3D2BWP30P140LVT U6 ( .A1(i_cmd[1]), .B1(n11), .B2(n10), .ZN(n14) );
  NR2D1BWP30P140LVT U7 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n11) );
  INVD1BWP30P140LVT U8 ( .I(i_cmd[6]), .ZN(n28) );
  NR3D1P5BWP30P140LVT U9 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .A3(n3), .ZN(n4) );
  INVD1BWP30P140LVT U10 ( .I(n7), .ZN(n8) );
  INVD6BWP30P140LVT U11 ( .I(n42), .ZN(n1) );
  INVD6BWP30P140LVT U12 ( .I(n2), .ZN(n167) );
  INVD6BWP30P140LVT U13 ( .I(n8), .ZN(n181) );
  INR2D2BWP30P140LVT U14 ( .A1(n19), .B1(n9), .ZN(n31) );
  NR2OPTPAD1BWP30P140LVT U15 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n19) );
  ND2OPTIBD2BWP30P140LVT U16 ( .A1(n4), .A2(n28), .ZN(n9) );
  INVD4BWP30P140LVT U17 ( .I(n17), .ZN(n180) );
  INVD2BWP30P140LVT U18 ( .I(n16), .ZN(n17) );
  ND2D1BWP30P140LVT U19 ( .A1(n19), .A2(n18), .ZN(n23) );
  INVD2BWP30P140LVT U20 ( .I(n13), .ZN(n179) );
  INVD1BWP30P140LVT U21 ( .I(i_cmd[4]), .ZN(n12) );
  INVD2BWP30P140LVT U22 ( .I(n179), .ZN(n156) );
  INVD2BWP30P140LVT U23 ( .I(n179), .ZN(n106) );
  NR4D0BWP30P140LVT U24 ( .A1(i_cmd[6]), .A2(n25), .A3(i_cmd[5]), .A4(n24), 
        .ZN(n26) );
  ND2D1BWP30P140LVT U25 ( .A1(n41), .A2(n40), .ZN(N402) );
  INR2D1BWP30P140LVT U26 ( .A1(i_en), .B1(rst), .ZN(n20) );
  INVD1BWP30P140LVT U27 ( .I(n20), .ZN(n3) );
  ND3D1BWP30P140LVT U28 ( .A1(n11), .A2(i_valid[1]), .A3(i_cmd[1]), .ZN(n5) );
  NR2OPTPAD1BWP30P140LVT U29 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n21) );
  ND3D1BWP30P140LVT U30 ( .A1(i_cmd[3]), .A2(n21), .A3(i_valid[3]), .ZN(n6) );
  INR2D1BWP30P140LVT U31 ( .A1(n31), .B1(n6), .ZN(n7) );
  INVD2BWP30P140LVT U32 ( .I(n9), .ZN(n10) );
  INR4D1BWP30P140LVT U33 ( .A1(i_valid[4]), .B1(i_cmd[0]), .B2(n12), .B3(n14), 
        .ZN(n13) );
  INVD1BWP30P140LVT U34 ( .I(i_cmd[0]), .ZN(n15) );
  INR4D1BWP30P140LVT U35 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n15), .B3(n14), 
        .ZN(n16) );
  NR4D0BWP30P140LVT U36 ( .A1(n167), .A2(n181), .A3(n156), .A4(n180), .ZN(n41)
         );
  INVD1BWP30P140LVT U37 ( .I(i_cmd[3]), .ZN(n18) );
  ND2OPTIBD1BWP30P140LVT U38 ( .A1(n21), .A2(n20), .ZN(n22) );
  NR2OPTPAD1BWP30P140LVT U39 ( .A1(n23), .A2(n22), .ZN(n27) );
  INVD1BWP30P140LVT U40 ( .I(i_cmd[7]), .ZN(n25) );
  INVD1BWP30P140LVT U41 ( .I(i_valid[7]), .ZN(n24) );
  AN2D2BWP30P140LVT U42 ( .A1(n27), .A2(n26), .Z(n184) );
  INVD2BWP30P140LVT U43 ( .I(n27), .ZN(n38) );
  IND2D1BWP30P140LVT U44 ( .A1(i_cmd[7]), .B1(i_valid[6]), .ZN(n29) );
  NR4D1BWP30P140LVT U45 ( .A1(n38), .A2(i_cmd[5]), .A3(n29), .A4(n28), .ZN(n30) );
  INVD2BWP30P140LVT U46 ( .I(n30), .ZN(n76) );
  INVD2BWP30P140LVT U47 ( .I(n76), .ZN(n173) );
  INVD2BWP30P140LVT U48 ( .I(n31), .ZN(n34) );
  INVD1BWP30P140LVT U49 ( .I(i_cmd[2]), .ZN(n33) );
  IND2D1BWP30P140LVT U50 ( .A1(i_cmd[3]), .B1(i_valid[2]), .ZN(n32) );
  NR4D1BWP30P140LVT U51 ( .A1(n34), .A2(i_cmd[1]), .A3(n33), .A4(n32), .ZN(n35) );
  INVD2BWP30P140LVT U52 ( .I(n35), .ZN(n43) );
  INVD2BWP30P140LVT U53 ( .I(n43), .ZN(n183) );
  INVD1BWP30P140LVT U54 ( .I(i_cmd[5]), .ZN(n37) );
  IND2D1BWP30P140LVT U55 ( .A1(i_cmd[7]), .B1(i_valid[5]), .ZN(n36) );
  NR4D0BWP30P140LVT U56 ( .A1(n184), .A2(n173), .A3(n183), .A4(n1), .ZN(n40)
         );
  AOI22D1BWP30P140LVT U57 ( .A1(n106), .A2(i_data_bus[140]), .B1(n180), .B2(
        i_data_bus[12]), .ZN(n47) );
  AOI22D1BWP30P140LVT U58 ( .A1(n167), .A2(i_data_bus[44]), .B1(n181), .B2(
        i_data_bus[108]), .ZN(n46) );
  INVD2BWP30P140LVT U59 ( .I(n76), .ZN(n182) );
  AOI22D1BWP30P140LVT U60 ( .A1(n182), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n45) );
  INVD2BWP30P140LVT U61 ( .I(n43), .ZN(n107) );
  AOI22D1BWP30P140LVT U62 ( .A1(n184), .A2(i_data_bus[236]), .B1(n107), .B2(
        i_data_bus[76]), .ZN(n44) );
  ND4D1BWP30P140LVT U63 ( .A1(n47), .A2(n46), .A3(n45), .A4(n44), .ZN(N381) );
  AOI22D1BWP30P140LVT U64 ( .A1(n106), .A2(i_data_bus[138]), .B1(n180), .B2(
        i_data_bus[10]), .ZN(n51) );
  AOI22D1BWP30P140LVT U65 ( .A1(n167), .A2(i_data_bus[42]), .B1(n181), .B2(
        i_data_bus[106]), .ZN(n50) );
  AOI22D1BWP30P140LVT U66 ( .A1(n182), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n49) );
  AOI22D1BWP30P140LVT U67 ( .A1(n184), .A2(i_data_bus[234]), .B1(n107), .B2(
        i_data_bus[74]), .ZN(n48) );
  ND4D1BWP30P140LVT U68 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(N379) );
  AOI22D1BWP30P140LVT U69 ( .A1(n106), .A2(i_data_bus[137]), .B1(n180), .B2(
        i_data_bus[9]), .ZN(n55) );
  AOI22D1BWP30P140LVT U70 ( .A1(n167), .A2(i_data_bus[41]), .B1(n181), .B2(
        i_data_bus[105]), .ZN(n54) );
  AOI22D1BWP30P140LVT U71 ( .A1(n182), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n53) );
  AOI22D1BWP30P140LVT U72 ( .A1(n184), .A2(i_data_bus[233]), .B1(n107), .B2(
        i_data_bus[73]), .ZN(n52) );
  ND4D1BWP30P140LVT U73 ( .A1(n55), .A2(n54), .A3(n53), .A4(n52), .ZN(N378) );
  AOI22D1BWP30P140LVT U74 ( .A1(n106), .A2(i_data_bus[135]), .B1(n180), .B2(
        i_data_bus[7]), .ZN(n59) );
  AOI22D1BWP30P140LVT U75 ( .A1(n167), .A2(i_data_bus[39]), .B1(n181), .B2(
        i_data_bus[103]), .ZN(n58) );
  AOI22D1BWP30P140LVT U76 ( .A1(n182), .A2(i_data_bus[199]), .B1(n1), .B2(
        i_data_bus[167]), .ZN(n57) );
  AOI22D1BWP30P140LVT U77 ( .A1(n184), .A2(i_data_bus[231]), .B1(n107), .B2(
        i_data_bus[71]), .ZN(n56) );
  ND4D1BWP30P140LVT U78 ( .A1(n59), .A2(n58), .A3(n57), .A4(n56), .ZN(N376) );
  AOI22D1BWP30P140LVT U79 ( .A1(n106), .A2(i_data_bus[134]), .B1(n180), .B2(
        i_data_bus[6]), .ZN(n63) );
  AOI22D1BWP30P140LVT U80 ( .A1(n167), .A2(i_data_bus[38]), .B1(n181), .B2(
        i_data_bus[102]), .ZN(n62) );
  AOI22D1BWP30P140LVT U81 ( .A1(n182), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n61) );
  AOI22D1BWP30P140LVT U82 ( .A1(n184), .A2(i_data_bus[230]), .B1(n107), .B2(
        i_data_bus[70]), .ZN(n60) );
  ND4D1BWP30P140LVT U83 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(N375) );
  AOI22D1BWP30P140LVT U84 ( .A1(n106), .A2(i_data_bus[132]), .B1(n180), .B2(
        i_data_bus[4]), .ZN(n67) );
  AOI22D1BWP30P140LVT U85 ( .A1(n167), .A2(i_data_bus[36]), .B1(n181), .B2(
        i_data_bus[100]), .ZN(n66) );
  AOI22D1BWP30P140LVT U86 ( .A1(n182), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n65) );
  AOI22D1BWP30P140LVT U87 ( .A1(n184), .A2(i_data_bus[228]), .B1(n107), .B2(
        i_data_bus[68]), .ZN(n64) );
  ND4D1BWP30P140LVT U88 ( .A1(n67), .A2(n66), .A3(n65), .A4(n64), .ZN(N373) );
  AOI22D1BWP30P140LVT U89 ( .A1(n106), .A2(i_data_bus[131]), .B1(n180), .B2(
        i_data_bus[3]), .ZN(n71) );
  AOI22D1BWP30P140LVT U90 ( .A1(n167), .A2(i_data_bus[35]), .B1(n181), .B2(
        i_data_bus[99]), .ZN(n70) );
  AOI22D1BWP30P140LVT U91 ( .A1(n182), .A2(i_data_bus[195]), .B1(n1), .B2(
        i_data_bus[163]), .ZN(n69) );
  AOI22D1BWP30P140LVT U92 ( .A1(n184), .A2(i_data_bus[227]), .B1(n107), .B2(
        i_data_bus[67]), .ZN(n68) );
  ND4D1BWP30P140LVT U93 ( .A1(n71), .A2(n70), .A3(n69), .A4(n68), .ZN(N372) );
  AOI22D1BWP30P140LVT U94 ( .A1(n106), .A2(i_data_bus[129]), .B1(n180), .B2(
        i_data_bus[1]), .ZN(n75) );
  AOI22D1BWP30P140LVT U95 ( .A1(n167), .A2(i_data_bus[33]), .B1(n181), .B2(
        i_data_bus[97]), .ZN(n74) );
  AOI22D1BWP30P140LVT U96 ( .A1(n182), .A2(i_data_bus[193]), .B1(n1), .B2(
        i_data_bus[161]), .ZN(n73) );
  AOI22D1BWP30P140LVT U97 ( .A1(n184), .A2(i_data_bus[225]), .B1(n107), .B2(
        i_data_bus[65]), .ZN(n72) );
  ND4D1BWP30P140LVT U98 ( .A1(n75), .A2(n74), .A3(n73), .A4(n72), .ZN(N370) );
  AOI22D1BWP30P140LVT U99 ( .A1(n106), .A2(i_data_bus[128]), .B1(n180), .B2(
        i_data_bus[0]), .ZN(n81) );
  AOI22D1BWP30P140LVT U100 ( .A1(n167), .A2(i_data_bus[32]), .B1(n181), .B2(
        i_data_bus[96]), .ZN(n80) );
  INVD1BWP30P140LVT U101 ( .I(n76), .ZN(n77) );
  AOI22D1BWP30P140LVT U102 ( .A1(n77), .A2(i_data_bus[192]), .B1(n1), .B2(
        i_data_bus[160]), .ZN(n79) );
  AOI22D1BWP30P140LVT U103 ( .A1(n184), .A2(i_data_bus[224]), .B1(n107), .B2(
        i_data_bus[64]), .ZN(n78) );
  ND4D1BWP30P140LVT U104 ( .A1(n81), .A2(n80), .A3(n79), .A4(n78), .ZN(N369)
         );
  AOI22D1BWP30P140LVT U105 ( .A1(n106), .A2(i_data_bus[139]), .B1(n180), .B2(
        i_data_bus[11]), .ZN(n85) );
  AOI22D1BWP30P140LVT U106 ( .A1(n167), .A2(i_data_bus[43]), .B1(n181), .B2(
        i_data_bus[107]), .ZN(n84) );
  AOI22D1BWP30P140LVT U107 ( .A1(n182), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n83) );
  AOI22D1BWP30P140LVT U108 ( .A1(n184), .A2(i_data_bus[235]), .B1(n107), .B2(
        i_data_bus[75]), .ZN(n82) );
  ND4D1BWP30P140LVT U109 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(N380)
         );
  AOI22D1BWP30P140LVT U110 ( .A1(n106), .A2(i_data_bus[136]), .B1(n180), .B2(
        i_data_bus[8]), .ZN(n89) );
  AOI22D1BWP30P140LVT U111 ( .A1(n167), .A2(i_data_bus[40]), .B1(n181), .B2(
        i_data_bus[104]), .ZN(n88) );
  AOI22D1BWP30P140LVT U112 ( .A1(n182), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n87) );
  AOI22D1BWP30P140LVT U113 ( .A1(n184), .A2(i_data_bus[232]), .B1(n107), .B2(
        i_data_bus[72]), .ZN(n86) );
  ND4D1BWP30P140LVT U114 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(N377)
         );
  AOI22D1BWP30P140LVT U115 ( .A1(n106), .A2(i_data_bus[133]), .B1(n180), .B2(
        i_data_bus[5]), .ZN(n93) );
  AOI22D1BWP30P140LVT U116 ( .A1(n167), .A2(i_data_bus[37]), .B1(n181), .B2(
        i_data_bus[101]), .ZN(n92) );
  AOI22D1BWP30P140LVT U117 ( .A1(n182), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n91) );
  AOI22D1BWP30P140LVT U118 ( .A1(n184), .A2(i_data_bus[229]), .B1(n107), .B2(
        i_data_bus[69]), .ZN(n90) );
  ND4D1BWP30P140LVT U119 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U120 ( .A1(n106), .A2(i_data_bus[130]), .B1(n180), .B2(
        i_data_bus[2]), .ZN(n97) );
  AOI22D1BWP30P140LVT U121 ( .A1(n167), .A2(i_data_bus[34]), .B1(n181), .B2(
        i_data_bus[98]), .ZN(n96) );
  AOI22D1BWP30P140LVT U122 ( .A1(n182), .A2(i_data_bus[194]), .B1(n1), .B2(
        i_data_bus[162]), .ZN(n95) );
  AOI22D1BWP30P140LVT U123 ( .A1(n184), .A2(i_data_bus[226]), .B1(n107), .B2(
        i_data_bus[66]), .ZN(n94) );
  ND4D1BWP30P140LVT U124 ( .A1(n97), .A2(n96), .A3(n95), .A4(n94), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U125 ( .A1(n106), .A2(i_data_bus[143]), .B1(n180), .B2(
        i_data_bus[15]), .ZN(n101) );
  AOI22D1BWP30P140LVT U126 ( .A1(n167), .A2(i_data_bus[47]), .B1(n181), .B2(
        i_data_bus[111]), .ZN(n100) );
  AOI22D1BWP30P140LVT U127 ( .A1(n182), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n99) );
  AOI22D1BWP30P140LVT U128 ( .A1(n184), .A2(i_data_bus[239]), .B1(n107), .B2(
        i_data_bus[79]), .ZN(n98) );
  ND4D1BWP30P140LVT U129 ( .A1(n101), .A2(n100), .A3(n99), .A4(n98), .ZN(N384)
         );
  AOI22D1BWP30P140LVT U130 ( .A1(n106), .A2(i_data_bus[142]), .B1(n180), .B2(
        i_data_bus[14]), .ZN(n105) );
  AOI22D1BWP30P140LVT U131 ( .A1(n167), .A2(i_data_bus[46]), .B1(n181), .B2(
        i_data_bus[110]), .ZN(n104) );
  AOI22D1BWP30P140LVT U132 ( .A1(n182), .A2(i_data_bus[206]), .B1(n1), .B2(
        i_data_bus[174]), .ZN(n103) );
  AOI22D1BWP30P140LVT U133 ( .A1(n184), .A2(i_data_bus[238]), .B1(n107), .B2(
        i_data_bus[78]), .ZN(n102) );
  ND4D1BWP30P140LVT U134 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U135 ( .A1(n106), .A2(i_data_bus[141]), .B1(n180), .B2(
        i_data_bus[13]), .ZN(n111) );
  AOI22D1BWP30P140LVT U136 ( .A1(n167), .A2(i_data_bus[45]), .B1(n181), .B2(
        i_data_bus[109]), .ZN(n110) );
  AOI22D1BWP30P140LVT U137 ( .A1(n182), .A2(i_data_bus[205]), .B1(n1), .B2(
        i_data_bus[173]), .ZN(n109) );
  AOI22D1BWP30P140LVT U138 ( .A1(n184), .A2(i_data_bus[237]), .B1(n107), .B2(
        i_data_bus[77]), .ZN(n108) );
  ND4D1BWP30P140LVT U139 ( .A1(n111), .A2(n110), .A3(n109), .A4(n108), .ZN(
        N382) );
  AOI22D1BWP30P140LVT U140 ( .A1(n156), .A2(i_data_bus[159]), .B1(n180), .B2(
        i_data_bus[31]), .ZN(n115) );
  AOI22D1BWP30P140LVT U141 ( .A1(n167), .A2(i_data_bus[63]), .B1(n181), .B2(
        i_data_bus[127]), .ZN(n114) );
  AOI22D1BWP30P140LVT U142 ( .A1(n173), .A2(i_data_bus[223]), .B1(n1), .B2(
        i_data_bus[191]), .ZN(n113) );
  AOI22D1BWP30P140LVT U143 ( .A1(n184), .A2(i_data_bus[255]), .B1(n183), .B2(
        i_data_bus[95]), .ZN(n112) );
  ND4D1BWP30P140LVT U144 ( .A1(n115), .A2(n114), .A3(n113), .A4(n112), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U145 ( .A1(n156), .A2(i_data_bus[158]), .B1(n180), .B2(
        i_data_bus[30]), .ZN(n119) );
  AOI22D1BWP30P140LVT U146 ( .A1(n167), .A2(i_data_bus[62]), .B1(n181), .B2(
        i_data_bus[126]), .ZN(n118) );
  AOI22D1BWP30P140LVT U147 ( .A1(n173), .A2(i_data_bus[222]), .B1(n1), .B2(
        i_data_bus[190]), .ZN(n117) );
  AOI22D1BWP30P140LVT U148 ( .A1(n184), .A2(i_data_bus[254]), .B1(n183), .B2(
        i_data_bus[94]), .ZN(n116) );
  ND4D1BWP30P140LVT U149 ( .A1(n119), .A2(n118), .A3(n117), .A4(n116), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U150 ( .A1(n156), .A2(i_data_bus[157]), .B1(n180), .B2(
        i_data_bus[29]), .ZN(n123) );
  AOI22D1BWP30P140LVT U151 ( .A1(n167), .A2(i_data_bus[61]), .B1(n181), .B2(
        i_data_bus[125]), .ZN(n122) );
  AOI22D1BWP30P140LVT U152 ( .A1(n173), .A2(i_data_bus[221]), .B1(n1), .B2(
        i_data_bus[189]), .ZN(n121) );
  AOI22D1BWP30P140LVT U153 ( .A1(n184), .A2(i_data_bus[253]), .B1(n183), .B2(
        i_data_bus[93]), .ZN(n120) );
  ND4D1BWP30P140LVT U154 ( .A1(n123), .A2(n122), .A3(n121), .A4(n120), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U155 ( .A1(n156), .A2(i_data_bus[156]), .B1(n180), .B2(
        i_data_bus[28]), .ZN(n127) );
  AOI22D1BWP30P140LVT U156 ( .A1(n167), .A2(i_data_bus[60]), .B1(n181), .B2(
        i_data_bus[124]), .ZN(n126) );
  AOI22D1BWP30P140LVT U157 ( .A1(n173), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n125) );
  AOI22D1BWP30P140LVT U158 ( .A1(n184), .A2(i_data_bus[252]), .B1(n183), .B2(
        i_data_bus[92]), .ZN(n124) );
  ND4D1BWP30P140LVT U159 ( .A1(n127), .A2(n126), .A3(n125), .A4(n124), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U160 ( .A1(n156), .A2(i_data_bus[155]), .B1(n180), .B2(
        i_data_bus[27]), .ZN(n131) );
  AOI22D1BWP30P140LVT U161 ( .A1(n167), .A2(i_data_bus[59]), .B1(n181), .B2(
        i_data_bus[123]), .ZN(n130) );
  AOI22D1BWP30P140LVT U162 ( .A1(n173), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n129) );
  AOI22D1BWP30P140LVT U163 ( .A1(n184), .A2(i_data_bus[251]), .B1(n183), .B2(
        i_data_bus[91]), .ZN(n128) );
  ND4D1BWP30P140LVT U164 ( .A1(n131), .A2(n130), .A3(n129), .A4(n128), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U165 ( .A1(n156), .A2(i_data_bus[154]), .B1(n180), .B2(
        i_data_bus[26]), .ZN(n135) );
  AOI22D1BWP30P140LVT U166 ( .A1(n167), .A2(i_data_bus[58]), .B1(n181), .B2(
        i_data_bus[122]), .ZN(n134) );
  AOI22D1BWP30P140LVT U167 ( .A1(n173), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n133) );
  AOI22D1BWP30P140LVT U168 ( .A1(n184), .A2(i_data_bus[250]), .B1(n183), .B2(
        i_data_bus[90]), .ZN(n132) );
  ND4D1BWP30P140LVT U169 ( .A1(n135), .A2(n134), .A3(n133), .A4(n132), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U170 ( .A1(n156), .A2(i_data_bus[153]), .B1(n180), .B2(
        i_data_bus[25]), .ZN(n139) );
  AOI22D1BWP30P140LVT U171 ( .A1(n167), .A2(i_data_bus[57]), .B1(n181), .B2(
        i_data_bus[121]), .ZN(n138) );
  AOI22D1BWP30P140LVT U172 ( .A1(n173), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n137) );
  AOI22D1BWP30P140LVT U173 ( .A1(n184), .A2(i_data_bus[249]), .B1(n183), .B2(
        i_data_bus[89]), .ZN(n136) );
  ND4D1BWP30P140LVT U174 ( .A1(n139), .A2(n138), .A3(n137), .A4(n136), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U175 ( .A1(n156), .A2(i_data_bus[152]), .B1(n180), .B2(
        i_data_bus[24]), .ZN(n143) );
  AOI22D1BWP30P140LVT U176 ( .A1(n167), .A2(i_data_bus[56]), .B1(n181), .B2(
        i_data_bus[120]), .ZN(n142) );
  AOI22D1BWP30P140LVT U177 ( .A1(n173), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n141) );
  AOI22D1BWP30P140LVT U178 ( .A1(n184), .A2(i_data_bus[248]), .B1(n183), .B2(
        i_data_bus[88]), .ZN(n140) );
  ND4D1BWP30P140LVT U179 ( .A1(n143), .A2(n142), .A3(n141), .A4(n140), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U180 ( .A1(n156), .A2(i_data_bus[151]), .B1(n180), .B2(
        i_data_bus[23]), .ZN(n147) );
  AOI22D1BWP30P140LVT U181 ( .A1(n167), .A2(i_data_bus[55]), .B1(n181), .B2(
        i_data_bus[119]), .ZN(n146) );
  AOI22D1BWP30P140LVT U182 ( .A1(n173), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n145) );
  AOI22D1BWP30P140LVT U183 ( .A1(n184), .A2(i_data_bus[247]), .B1(n183), .B2(
        i_data_bus[87]), .ZN(n144) );
  ND4D1BWP30P140LVT U184 ( .A1(n147), .A2(n146), .A3(n145), .A4(n144), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U185 ( .A1(n156), .A2(i_data_bus[150]), .B1(n180), .B2(
        i_data_bus[22]), .ZN(n151) );
  AOI22D1BWP30P140LVT U186 ( .A1(n167), .A2(i_data_bus[54]), .B1(n181), .B2(
        i_data_bus[118]), .ZN(n150) );
  AOI22D1BWP30P140LVT U187 ( .A1(n173), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n149) );
  AOI22D1BWP30P140LVT U188 ( .A1(n184), .A2(i_data_bus[246]), .B1(n183), .B2(
        i_data_bus[86]), .ZN(n148) );
  ND4D1BWP30P140LVT U189 ( .A1(n151), .A2(n150), .A3(n149), .A4(n148), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U190 ( .A1(n156), .A2(i_data_bus[149]), .B1(n180), .B2(
        i_data_bus[21]), .ZN(n155) );
  AOI22D1BWP30P140LVT U191 ( .A1(n167), .A2(i_data_bus[53]), .B1(n181), .B2(
        i_data_bus[117]), .ZN(n154) );
  AOI22D1BWP30P140LVT U192 ( .A1(n173), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n153) );
  AOI22D1BWP30P140LVT U193 ( .A1(n184), .A2(i_data_bus[245]), .B1(n183), .B2(
        i_data_bus[85]), .ZN(n152) );
  ND4D1BWP30P140LVT U194 ( .A1(n155), .A2(n154), .A3(n153), .A4(n152), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U195 ( .A1(n156), .A2(i_data_bus[148]), .B1(n180), .B2(
        i_data_bus[20]), .ZN(n160) );
  AOI22D1BWP30P140LVT U196 ( .A1(n167), .A2(i_data_bus[52]), .B1(n181), .B2(
        i_data_bus[116]), .ZN(n159) );
  AOI22D1BWP30P140LVT U197 ( .A1(n173), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n158) );
  AOI22D1BWP30P140LVT U198 ( .A1(n184), .A2(i_data_bus[244]), .B1(n183), .B2(
        i_data_bus[84]), .ZN(n157) );
  ND4D1BWP30P140LVT U199 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(
        N389) );
  INVD1BWP30P140LVT U200 ( .I(i_data_bus[147]), .ZN(n161) );
  MAOI22D1BWP30P140LVT U201 ( .A1(n180), .A2(i_data_bus[19]), .B1(n179), .B2(
        n161), .ZN(n165) );
  AOI22D1BWP30P140LVT U202 ( .A1(n167), .A2(i_data_bus[51]), .B1(n181), .B2(
        i_data_bus[115]), .ZN(n164) );
  AOI22D1BWP30P140LVT U203 ( .A1(n173), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n163) );
  AOI22D1BWP30P140LVT U204 ( .A1(n184), .A2(i_data_bus[243]), .B1(n183), .B2(
        i_data_bus[83]), .ZN(n162) );
  ND4D1BWP30P140LVT U205 ( .A1(n165), .A2(n164), .A3(n163), .A4(n162), .ZN(
        N388) );
  INVD1BWP30P140LVT U206 ( .I(i_data_bus[146]), .ZN(n166) );
  MAOI22D1BWP30P140LVT U207 ( .A1(n180), .A2(i_data_bus[18]), .B1(n179), .B2(
        n166), .ZN(n171) );
  AOI22D1BWP30P140LVT U208 ( .A1(n167), .A2(i_data_bus[50]), .B1(n181), .B2(
        i_data_bus[114]), .ZN(n170) );
  AOI22D1BWP30P140LVT U209 ( .A1(n173), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n169) );
  AOI22D1BWP30P140LVT U210 ( .A1(n184), .A2(i_data_bus[242]), .B1(n183), .B2(
        i_data_bus[82]), .ZN(n168) );
  ND4D1BWP30P140LVT U211 ( .A1(n171), .A2(n170), .A3(n169), .A4(n168), .ZN(
        N387) );
  INVD1BWP30P140LVT U212 ( .I(i_data_bus[145]), .ZN(n172) );
  MAOI22D1BWP30P140LVT U213 ( .A1(n180), .A2(i_data_bus[17]), .B1(n179), .B2(
        n172), .ZN(n177) );
  AOI22D1BWP30P140LVT U214 ( .A1(n167), .A2(i_data_bus[49]), .B1(n181), .B2(
        i_data_bus[113]), .ZN(n176) );
  AOI22D1BWP30P140LVT U215 ( .A1(n173), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n175) );
  AOI22D1BWP30P140LVT U216 ( .A1(n184), .A2(i_data_bus[241]), .B1(n183), .B2(
        i_data_bus[81]), .ZN(n174) );
  ND4D1BWP30P140LVT U217 ( .A1(n177), .A2(n176), .A3(n175), .A4(n174), .ZN(
        N386) );
  INVD1BWP30P140LVT U218 ( .I(i_data_bus[144]), .ZN(n178) );
  MAOI22D1BWP30P140LVT U219 ( .A1(n180), .A2(i_data_bus[16]), .B1(n179), .B2(
        n178), .ZN(n188) );
  AOI22D1BWP30P140LVT U220 ( .A1(n167), .A2(i_data_bus[48]), .B1(n181), .B2(
        i_data_bus[112]), .ZN(n187) );
  AOI22D1BWP30P140LVT U221 ( .A1(n182), .A2(i_data_bus[208]), .B1(n1), .B2(
        i_data_bus[176]), .ZN(n186) );
  AOI22D1BWP30P140LVT U222 ( .A1(n184), .A2(i_data_bus[240]), .B1(n183), .B2(
        i_data_bus[80]), .ZN(n185) );
  ND4D1BWP30P140LVT U223 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .ZN(
        N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_4 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD4BWP30P140LVT U3 ( .I(n14), .ZN(n174) );
  INVD6BWP30P140LVT U4 ( .I(n50), .ZN(n1) );
  INVD2BWP30P140LVT U5 ( .I(n13), .ZN(n14) );
  INVD1BWP30P140LVT U6 ( .I(n10), .ZN(n49) );
  INVD2BWP30P140LVT U7 ( .I(n35), .ZN(n50) );
  INR2D6BWP30P140LVT U8 ( .A1(n27), .B1(n5), .ZN(n176) );
  INR2D2BWP30P140LVT U9 ( .A1(n27), .B1(n3), .ZN(n177) );
  NR4D1BWP30P140LVT U10 ( .A1(n34), .A2(i_cmd[5]), .A3(n25), .A4(n24), .ZN(n26) );
  INVD0P7BWP30P140LVT U11 ( .I(i_cmd[2]), .ZN(n29) );
  CKND2D2BWP30P140LVT U12 ( .A1(n4), .A2(i_cmd[3]), .ZN(n5) );
  NR2OPTPAD1BWP30P140LVT U13 ( .A1(i_cmd[6]), .A2(i_cmd[5]), .ZN(n21) );
  INVD1BWP30P140LVT U14 ( .I(n31), .ZN(n51) );
  INVD1BWP30P140LVT U15 ( .I(i_cmd[6]), .ZN(n24) );
  INVD1BWP30P140LVT U16 ( .I(i_cmd[0]), .ZN(n12) );
  IND3D2BWP30P140LVT U17 ( .A1(i_cmd[1]), .B1(n8), .B2(n7), .ZN(n11) );
  NR2OPTPAD1BWP30P140LVT U18 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n8) );
  NR4D1BWP30P140LVT U19 ( .A1(n30), .A2(i_cmd[1]), .A3(n29), .A4(n28), .ZN(n31) );
  ND2OPTIBD2BWP30P140LVT U20 ( .A1(n21), .A2(n2), .ZN(n6) );
  NR4D2BWP30P140LVT U21 ( .A1(n34), .A2(i_cmd[6]), .A3(n33), .A4(n32), .ZN(n35) );
  AOI22D1BWP30P140LVT U22 ( .A1(n175), .A2(i_data_bus[145]), .B1(n174), .B2(
        i_data_bus[17]), .ZN(n48) );
  INVD1BWP30P140LVT U23 ( .I(i_cmd[5]), .ZN(n33) );
  INVD1BWP30P140LVT U24 ( .I(i_cmd[4]), .ZN(n9) );
  INR2D1BWP30P140LVT U25 ( .A1(n15), .B1(i_cmd[7]), .ZN(n2) );
  NR2OPTPAD1BWP30P140LVT U26 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n18) );
  INVD1BWP30P140LVT U27 ( .I(n6), .ZN(n7) );
  ND2D1BWP30P140LVT U28 ( .A1(n37), .A2(n36), .ZN(N402) );
  NR2OPTPAD1BWP30P140LVT U29 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n20) );
  INR2D1BWP30P140LVT U30 ( .A1(i_en), .B1(rst), .ZN(n15) );
  INR2D2BWP30P140LVT U31 ( .A1(n20), .B1(n6), .ZN(n27) );
  ND3D1BWP30P140LVT U32 ( .A1(n8), .A2(i_valid[1]), .A3(i_cmd[1]), .ZN(n3) );
  BUFFD4BWP30P140LVT U33 ( .I(n177), .Z(n145) );
  CKAN2D1BWP30P140LVT U34 ( .A1(n18), .A2(i_valid[3]), .Z(n4) );
  INR4D1BWP30P140LVT U35 ( .A1(i_valid[4]), .B1(i_cmd[0]), .B2(n9), .B3(n11), 
        .ZN(n10) );
  INVD2BWP30P140LVT U36 ( .I(n49), .ZN(n175) );
  INR4D1BWP30P140LVT U37 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n12), .B3(n11), 
        .ZN(n13) );
  NR4D0BWP30P140LVT U38 ( .A1(n145), .A2(n176), .A3(n175), .A4(n174), .ZN(n37)
         );
  INVD1BWP30P140LVT U39 ( .I(n15), .ZN(n16) );
  NR2OPTPAD1BWP30P140LVT U40 ( .A1(i_cmd[3]), .A2(n16), .ZN(n17) );
  ND2OPTIBD1BWP30P140LVT U41 ( .A1(n18), .A2(n17), .ZN(n19) );
  INR2D2BWP30P140LVT U42 ( .A1(n20), .B1(n19), .ZN(n23) );
  ND3D1BWP30P140LVT U43 ( .A1(n21), .A2(i_valid[7]), .A3(i_cmd[7]), .ZN(n22)
         );
  INR2D6BWP30P140LVT U44 ( .A1(n23), .B1(n22), .ZN(n180) );
  INVD2BWP30P140LVT U45 ( .I(n23), .ZN(n34) );
  IND2D1BWP30P140LVT U46 ( .A1(i_cmd[7]), .B1(i_valid[6]), .ZN(n25) );
  INVD2BWP30P140LVT U47 ( .I(n26), .ZN(n100) );
  INVD2BWP30P140LVT U48 ( .I(n100), .ZN(n178) );
  INVD2BWP30P140LVT U49 ( .I(n27), .ZN(n30) );
  IND2D1BWP30P140LVT U50 ( .A1(i_cmd[3]), .B1(i_valid[2]), .ZN(n28) );
  INVD2BWP30P140LVT U51 ( .I(n51), .ZN(n179) );
  IND2D1BWP30P140LVT U52 ( .A1(i_cmd[7]), .B1(i_valid[5]), .ZN(n32) );
  NR4D0BWP30P140LVT U53 ( .A1(n180), .A2(n178), .A3(n179), .A4(n1), .ZN(n36)
         );
  AOI22D1BWP30P140LVT U54 ( .A1(n175), .A2(i_data_bus[144]), .B1(n174), .B2(
        i_data_bus[16]), .ZN(n44) );
  INVD2BWP30P140LVT U55 ( .I(n100), .ZN(n115) );
  AOI22D1BWP30P140LVT U56 ( .A1(n115), .A2(i_data_bus[208]), .B1(n1), .B2(
        i_data_bus[176]), .ZN(n43) );
  ND2OPTIBD1BWP30P140LVT U57 ( .A1(n180), .A2(i_data_bus[240]), .ZN(n40) );
  ND2D1BWP30P140LVT U58 ( .A1(n176), .A2(i_data_bus[112]), .ZN(n39) );
  ND2OPTIBD1BWP30P140LVT U59 ( .A1(n177), .A2(i_data_bus[48]), .ZN(n38) );
  ND3D1BWP30P140LVT U60 ( .A1(n40), .A2(n39), .A3(n38), .ZN(n41) );
  AOI21D1BWP30P140LVT U61 ( .A1(n179), .A2(i_data_bus[80]), .B(n41), .ZN(n42)
         );
  ND3D1BWP30P140LVT U62 ( .A1(n44), .A2(n43), .A3(n42), .ZN(N385) );
  AOI22D1BWP30P140LVT U63 ( .A1(n145), .A2(i_data_bus[49]), .B1(n176), .B2(
        i_data_bus[113]), .ZN(n47) );
  AOI22D1BWP30P140LVT U64 ( .A1(n178), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n46) );
  AOI22D1BWP30P140LVT U65 ( .A1(n180), .A2(i_data_bus[241]), .B1(n179), .B2(
        i_data_bus[81]), .ZN(n45) );
  ND4D1BWP30P140LVT U66 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(N386) );
  INVD2BWP30P140LVT U67 ( .I(n49), .ZN(n114) );
  AOI22D1BWP30P140LVT U68 ( .A1(n114), .A2(i_data_bus[140]), .B1(n174), .B2(
        i_data_bus[12]), .ZN(n55) );
  AOI22D1BWP30P140LVT U69 ( .A1(n145), .A2(i_data_bus[44]), .B1(n176), .B2(
        i_data_bus[108]), .ZN(n54) );
  AOI22D1BWP30P140LVT U70 ( .A1(n115), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n53) );
  INVD2BWP30P140LVT U71 ( .I(n51), .ZN(n116) );
  AOI22D1BWP30P140LVT U72 ( .A1(n180), .A2(i_data_bus[236]), .B1(n116), .B2(
        i_data_bus[76]), .ZN(n52) );
  ND4D1BWP30P140LVT U73 ( .A1(n55), .A2(n54), .A3(n53), .A4(n52), .ZN(N381) );
  AOI22D1BWP30P140LVT U74 ( .A1(n114), .A2(i_data_bus[139]), .B1(n174), .B2(
        i_data_bus[11]), .ZN(n59) );
  AOI22D1BWP30P140LVT U75 ( .A1(n145), .A2(i_data_bus[43]), .B1(n176), .B2(
        i_data_bus[107]), .ZN(n58) );
  AOI22D1BWP30P140LVT U76 ( .A1(n115), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n57) );
  AOI22D1BWP30P140LVT U77 ( .A1(n180), .A2(i_data_bus[235]), .B1(n116), .B2(
        i_data_bus[75]), .ZN(n56) );
  ND4D1BWP30P140LVT U78 ( .A1(n59), .A2(n58), .A3(n57), .A4(n56), .ZN(N380) );
  AOI22D1BWP30P140LVT U79 ( .A1(n114), .A2(i_data_bus[138]), .B1(n174), .B2(
        i_data_bus[10]), .ZN(n63) );
  AOI22D1BWP30P140LVT U80 ( .A1(n145), .A2(i_data_bus[42]), .B1(n176), .B2(
        i_data_bus[106]), .ZN(n62) );
  AOI22D1BWP30P140LVT U81 ( .A1(n115), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n61) );
  AOI22D1BWP30P140LVT U82 ( .A1(n180), .A2(i_data_bus[234]), .B1(n116), .B2(
        i_data_bus[74]), .ZN(n60) );
  ND4D1BWP30P140LVT U83 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(N379) );
  AOI22D1BWP30P140LVT U84 ( .A1(n114), .A2(i_data_bus[137]), .B1(n174), .B2(
        i_data_bus[9]), .ZN(n67) );
  AOI22D1BWP30P140LVT U85 ( .A1(n145), .A2(i_data_bus[41]), .B1(n176), .B2(
        i_data_bus[105]), .ZN(n66) );
  AOI22D1BWP30P140LVT U86 ( .A1(n115), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n65) );
  AOI22D1BWP30P140LVT U87 ( .A1(n180), .A2(i_data_bus[233]), .B1(n116), .B2(
        i_data_bus[73]), .ZN(n64) );
  ND4D1BWP30P140LVT U88 ( .A1(n67), .A2(n66), .A3(n65), .A4(n64), .ZN(N378) );
  AOI22D1BWP30P140LVT U89 ( .A1(n114), .A2(i_data_bus[136]), .B1(n174), .B2(
        i_data_bus[8]), .ZN(n71) );
  AOI22D1BWP30P140LVT U90 ( .A1(n145), .A2(i_data_bus[40]), .B1(n176), .B2(
        i_data_bus[104]), .ZN(n70) );
  AOI22D1BWP30P140LVT U91 ( .A1(n115), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n69) );
  AOI22D1BWP30P140LVT U92 ( .A1(n180), .A2(i_data_bus[232]), .B1(n116), .B2(
        i_data_bus[72]), .ZN(n68) );
  ND4D1BWP30P140LVT U93 ( .A1(n71), .A2(n70), .A3(n69), .A4(n68), .ZN(N377) );
  AOI22D1BWP30P140LVT U94 ( .A1(n114), .A2(i_data_bus[135]), .B1(n174), .B2(
        i_data_bus[7]), .ZN(n75) );
  AOI22D1BWP30P140LVT U95 ( .A1(n145), .A2(i_data_bus[39]), .B1(n176), .B2(
        i_data_bus[103]), .ZN(n74) );
  AOI22D1BWP30P140LVT U96 ( .A1(n115), .A2(i_data_bus[199]), .B1(n1), .B2(
        i_data_bus[167]), .ZN(n73) );
  AOI22D1BWP30P140LVT U97 ( .A1(n180), .A2(i_data_bus[231]), .B1(n116), .B2(
        i_data_bus[71]), .ZN(n72) );
  ND4D1BWP30P140LVT U98 ( .A1(n75), .A2(n74), .A3(n73), .A4(n72), .ZN(N376) );
  AOI22D1BWP30P140LVT U99 ( .A1(n114), .A2(i_data_bus[134]), .B1(n174), .B2(
        i_data_bus[6]), .ZN(n79) );
  AOI22D1BWP30P140LVT U100 ( .A1(n145), .A2(i_data_bus[38]), .B1(n176), .B2(
        i_data_bus[102]), .ZN(n78) );
  AOI22D1BWP30P140LVT U101 ( .A1(n115), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n77) );
  AOI22D1BWP30P140LVT U102 ( .A1(n180), .A2(i_data_bus[230]), .B1(n116), .B2(
        i_data_bus[70]), .ZN(n76) );
  ND4D1BWP30P140LVT U103 ( .A1(n79), .A2(n78), .A3(n77), .A4(n76), .ZN(N375)
         );
  AOI22D1BWP30P140LVT U104 ( .A1(n114), .A2(i_data_bus[133]), .B1(n174), .B2(
        i_data_bus[5]), .ZN(n83) );
  AOI22D1BWP30P140LVT U105 ( .A1(n145), .A2(i_data_bus[37]), .B1(n176), .B2(
        i_data_bus[101]), .ZN(n82) );
  AOI22D1BWP30P140LVT U106 ( .A1(n115), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n81) );
  AOI22D1BWP30P140LVT U107 ( .A1(n180), .A2(i_data_bus[229]), .B1(n116), .B2(
        i_data_bus[69]), .ZN(n80) );
  ND4D1BWP30P140LVT U108 ( .A1(n83), .A2(n82), .A3(n81), .A4(n80), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U109 ( .A1(n114), .A2(i_data_bus[132]), .B1(n174), .B2(
        i_data_bus[4]), .ZN(n87) );
  AOI22D1BWP30P140LVT U110 ( .A1(n145), .A2(i_data_bus[36]), .B1(n176), .B2(
        i_data_bus[100]), .ZN(n86) );
  AOI22D1BWP30P140LVT U111 ( .A1(n115), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n85) );
  AOI22D1BWP30P140LVT U112 ( .A1(n180), .A2(i_data_bus[228]), .B1(n116), .B2(
        i_data_bus[68]), .ZN(n84) );
  ND4D1BWP30P140LVT U113 ( .A1(n87), .A2(n86), .A3(n85), .A4(n84), .ZN(N373)
         );
  AOI22D1BWP30P140LVT U114 ( .A1(n114), .A2(i_data_bus[131]), .B1(n174), .B2(
        i_data_bus[3]), .ZN(n91) );
  AOI22D1BWP30P140LVT U115 ( .A1(n145), .A2(i_data_bus[35]), .B1(n176), .B2(
        i_data_bus[99]), .ZN(n90) );
  AOI22D1BWP30P140LVT U116 ( .A1(n115), .A2(i_data_bus[195]), .B1(n1), .B2(
        i_data_bus[163]), .ZN(n89) );
  AOI22D1BWP30P140LVT U117 ( .A1(n180), .A2(i_data_bus[227]), .B1(n116), .B2(
        i_data_bus[67]), .ZN(n88) );
  ND4D1BWP30P140LVT U118 ( .A1(n91), .A2(n90), .A3(n89), .A4(n88), .ZN(N372)
         );
  AOI22D1BWP30P140LVT U119 ( .A1(n114), .A2(i_data_bus[130]), .B1(n174), .B2(
        i_data_bus[2]), .ZN(n95) );
  AOI22D1BWP30P140LVT U120 ( .A1(n145), .A2(i_data_bus[34]), .B1(n176), .B2(
        i_data_bus[98]), .ZN(n94) );
  AOI22D1BWP30P140LVT U121 ( .A1(n115), .A2(i_data_bus[194]), .B1(n1), .B2(
        i_data_bus[162]), .ZN(n93) );
  AOI22D1BWP30P140LVT U122 ( .A1(n180), .A2(i_data_bus[226]), .B1(n116), .B2(
        i_data_bus[66]), .ZN(n92) );
  ND4D1BWP30P140LVT U123 ( .A1(n95), .A2(n94), .A3(n93), .A4(n92), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U124 ( .A1(n114), .A2(i_data_bus[129]), .B1(n174), .B2(
        i_data_bus[1]), .ZN(n99) );
  AOI22D1BWP30P140LVT U125 ( .A1(n145), .A2(i_data_bus[33]), .B1(n176), .B2(
        i_data_bus[97]), .ZN(n98) );
  AOI22D1BWP30P140LVT U126 ( .A1(n115), .A2(i_data_bus[193]), .B1(n1), .B2(
        i_data_bus[161]), .ZN(n97) );
  AOI22D1BWP30P140LVT U127 ( .A1(n180), .A2(i_data_bus[225]), .B1(n116), .B2(
        i_data_bus[65]), .ZN(n96) );
  ND4D1BWP30P140LVT U128 ( .A1(n99), .A2(n98), .A3(n97), .A4(n96), .ZN(N370)
         );
  AOI22D1BWP30P140LVT U129 ( .A1(n114), .A2(i_data_bus[128]), .B1(n174), .B2(
        i_data_bus[0]), .ZN(n105) );
  AOI22D1BWP30P140LVT U130 ( .A1(n145), .A2(i_data_bus[32]), .B1(n176), .B2(
        i_data_bus[96]), .ZN(n104) );
  INVD1BWP30P140LVT U131 ( .I(n100), .ZN(n101) );
  AOI22D1BWP30P140LVT U132 ( .A1(n101), .A2(i_data_bus[192]), .B1(n1), .B2(
        i_data_bus[160]), .ZN(n103) );
  AOI22D1BWP30P140LVT U133 ( .A1(n180), .A2(i_data_bus[224]), .B1(n116), .B2(
        i_data_bus[64]), .ZN(n102) );
  ND4D1BWP30P140LVT U134 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .ZN(
        N369) );
  AOI22D1BWP30P140LVT U135 ( .A1(n114), .A2(i_data_bus[143]), .B1(n174), .B2(
        i_data_bus[15]), .ZN(n109) );
  AOI22D1BWP30P140LVT U136 ( .A1(n145), .A2(i_data_bus[47]), .B1(n176), .B2(
        i_data_bus[111]), .ZN(n108) );
  AOI22D1BWP30P140LVT U137 ( .A1(n115), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n107) );
  AOI22D1BWP30P140LVT U138 ( .A1(n180), .A2(i_data_bus[239]), .B1(n116), .B2(
        i_data_bus[79]), .ZN(n106) );
  ND4D1BWP30P140LVT U139 ( .A1(n109), .A2(n108), .A3(n107), .A4(n106), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U140 ( .A1(n114), .A2(i_data_bus[142]), .B1(n174), .B2(
        i_data_bus[14]), .ZN(n113) );
  AOI22D1BWP30P140LVT U141 ( .A1(n145), .A2(i_data_bus[46]), .B1(n176), .B2(
        i_data_bus[110]), .ZN(n112) );
  AOI22D1BWP30P140LVT U142 ( .A1(n115), .A2(i_data_bus[206]), .B1(n1), .B2(
        i_data_bus[174]), .ZN(n111) );
  AOI22D1BWP30P140LVT U143 ( .A1(n180), .A2(i_data_bus[238]), .B1(n116), .B2(
        i_data_bus[78]), .ZN(n110) );
  ND4D1BWP30P140LVT U144 ( .A1(n113), .A2(n112), .A3(n111), .A4(n110), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U145 ( .A1(n114), .A2(i_data_bus[141]), .B1(n174), .B2(
        i_data_bus[13]), .ZN(n120) );
  AOI22D1BWP30P140LVT U146 ( .A1(n145), .A2(i_data_bus[45]), .B1(n176), .B2(
        i_data_bus[109]), .ZN(n119) );
  AOI22D1BWP30P140LVT U147 ( .A1(n115), .A2(i_data_bus[205]), .B1(n1), .B2(
        i_data_bus[173]), .ZN(n118) );
  AOI22D1BWP30P140LVT U148 ( .A1(n180), .A2(i_data_bus[237]), .B1(n116), .B2(
        i_data_bus[77]), .ZN(n117) );
  ND4D1BWP30P140LVT U149 ( .A1(n120), .A2(n119), .A3(n118), .A4(n117), .ZN(
        N382) );
  AOI22D1BWP30P140LVT U150 ( .A1(n175), .A2(i_data_bus[159]), .B1(n174), .B2(
        i_data_bus[31]), .ZN(n124) );
  AOI22D1BWP30P140LVT U151 ( .A1(n145), .A2(i_data_bus[63]), .B1(n176), .B2(
        i_data_bus[127]), .ZN(n123) );
  AOI22D1BWP30P140LVT U152 ( .A1(n178), .A2(i_data_bus[223]), .B1(n1), .B2(
        i_data_bus[191]), .ZN(n122) );
  AOI22D1BWP30P140LVT U153 ( .A1(n180), .A2(i_data_bus[255]), .B1(n179), .B2(
        i_data_bus[95]), .ZN(n121) );
  ND4D1BWP30P140LVT U154 ( .A1(n124), .A2(n123), .A3(n122), .A4(n121), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U155 ( .A1(n175), .A2(i_data_bus[158]), .B1(n174), .B2(
        i_data_bus[30]), .ZN(n128) );
  AOI22D1BWP30P140LVT U156 ( .A1(n145), .A2(i_data_bus[62]), .B1(n176), .B2(
        i_data_bus[126]), .ZN(n127) );
  AOI22D1BWP30P140LVT U157 ( .A1(n178), .A2(i_data_bus[222]), .B1(n1), .B2(
        i_data_bus[190]), .ZN(n126) );
  AOI22D1BWP30P140LVT U158 ( .A1(n180), .A2(i_data_bus[254]), .B1(n179), .B2(
        i_data_bus[94]), .ZN(n125) );
  ND4D1BWP30P140LVT U159 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U160 ( .A1(n175), .A2(i_data_bus[157]), .B1(n174), .B2(
        i_data_bus[29]), .ZN(n132) );
  AOI22D1BWP30P140LVT U161 ( .A1(n145), .A2(i_data_bus[61]), .B1(n176), .B2(
        i_data_bus[125]), .ZN(n131) );
  AOI22D1BWP30P140LVT U162 ( .A1(n178), .A2(i_data_bus[221]), .B1(n1), .B2(
        i_data_bus[189]), .ZN(n130) );
  AOI22D1BWP30P140LVT U163 ( .A1(n180), .A2(i_data_bus[253]), .B1(n179), .B2(
        i_data_bus[93]), .ZN(n129) );
  ND4D1BWP30P140LVT U164 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U165 ( .A1(n175), .A2(i_data_bus[156]), .B1(n174), .B2(
        i_data_bus[28]), .ZN(n136) );
  AOI22D1BWP30P140LVT U166 ( .A1(n145), .A2(i_data_bus[60]), .B1(n176), .B2(
        i_data_bus[124]), .ZN(n135) );
  AOI22D1BWP30P140LVT U167 ( .A1(n178), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n134) );
  AOI22D1BWP30P140LVT U168 ( .A1(n180), .A2(i_data_bus[252]), .B1(n179), .B2(
        i_data_bus[92]), .ZN(n133) );
  ND4D1BWP30P140LVT U169 ( .A1(n136), .A2(n135), .A3(n134), .A4(n133), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U170 ( .A1(n175), .A2(i_data_bus[155]), .B1(n174), .B2(
        i_data_bus[27]), .ZN(n140) );
  AOI22D1BWP30P140LVT U171 ( .A1(n145), .A2(i_data_bus[59]), .B1(n176), .B2(
        i_data_bus[123]), .ZN(n139) );
  AOI22D1BWP30P140LVT U172 ( .A1(n178), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n138) );
  AOI22D1BWP30P140LVT U173 ( .A1(n180), .A2(i_data_bus[251]), .B1(n179), .B2(
        i_data_bus[91]), .ZN(n137) );
  ND4D1BWP30P140LVT U174 ( .A1(n140), .A2(n139), .A3(n138), .A4(n137), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U175 ( .A1(n175), .A2(i_data_bus[154]), .B1(n174), .B2(
        i_data_bus[26]), .ZN(n144) );
  AOI22D1BWP30P140LVT U176 ( .A1(n145), .A2(i_data_bus[58]), .B1(n176), .B2(
        i_data_bus[122]), .ZN(n143) );
  AOI22D1BWP30P140LVT U177 ( .A1(n178), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n142) );
  AOI22D1BWP30P140LVT U178 ( .A1(n180), .A2(i_data_bus[250]), .B1(n179), .B2(
        i_data_bus[90]), .ZN(n141) );
  ND4D1BWP30P140LVT U179 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U180 ( .A1(n175), .A2(i_data_bus[153]), .B1(n174), .B2(
        i_data_bus[25]), .ZN(n149) );
  AOI22D1BWP30P140LVT U181 ( .A1(n145), .A2(i_data_bus[57]), .B1(n176), .B2(
        i_data_bus[121]), .ZN(n148) );
  AOI22D1BWP30P140LVT U182 ( .A1(n178), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n147) );
  AOI22D1BWP30P140LVT U183 ( .A1(n180), .A2(i_data_bus[249]), .B1(n179), .B2(
        i_data_bus[89]), .ZN(n146) );
  ND4D1BWP30P140LVT U184 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U185 ( .A1(n175), .A2(i_data_bus[152]), .B1(n174), .B2(
        i_data_bus[24]), .ZN(n153) );
  AOI22D1BWP30P140LVT U186 ( .A1(n177), .A2(i_data_bus[56]), .B1(n176), .B2(
        i_data_bus[120]), .ZN(n152) );
  AOI22D1BWP30P140LVT U187 ( .A1(n178), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n151) );
  AOI22D1BWP30P140LVT U188 ( .A1(n180), .A2(i_data_bus[248]), .B1(n179), .B2(
        i_data_bus[88]), .ZN(n150) );
  ND4D1BWP30P140LVT U189 ( .A1(n153), .A2(n152), .A3(n151), .A4(n150), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U190 ( .A1(n175), .A2(i_data_bus[151]), .B1(n174), .B2(
        i_data_bus[23]), .ZN(n157) );
  AOI22D1BWP30P140LVT U191 ( .A1(n177), .A2(i_data_bus[55]), .B1(n176), .B2(
        i_data_bus[119]), .ZN(n156) );
  AOI22D1BWP30P140LVT U192 ( .A1(n178), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n155) );
  AOI22D1BWP30P140LVT U193 ( .A1(n180), .A2(i_data_bus[247]), .B1(n179), .B2(
        i_data_bus[87]), .ZN(n154) );
  ND4D1BWP30P140LVT U194 ( .A1(n157), .A2(n156), .A3(n155), .A4(n154), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U195 ( .A1(n175), .A2(i_data_bus[150]), .B1(n174), .B2(
        i_data_bus[22]), .ZN(n161) );
  AOI22D1BWP30P140LVT U196 ( .A1(n177), .A2(i_data_bus[54]), .B1(n176), .B2(
        i_data_bus[118]), .ZN(n160) );
  AOI22D1BWP30P140LVT U197 ( .A1(n178), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n159) );
  AOI22D1BWP30P140LVT U198 ( .A1(n180), .A2(i_data_bus[246]), .B1(n179), .B2(
        i_data_bus[86]), .ZN(n158) );
  ND4D1BWP30P140LVT U199 ( .A1(n161), .A2(n160), .A3(n159), .A4(n158), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U200 ( .A1(n175), .A2(i_data_bus[149]), .B1(n174), .B2(
        i_data_bus[21]), .ZN(n165) );
  AOI22D1BWP30P140LVT U201 ( .A1(n177), .A2(i_data_bus[53]), .B1(n176), .B2(
        i_data_bus[117]), .ZN(n164) );
  AOI22D1BWP30P140LVT U202 ( .A1(n178), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n163) );
  AOI22D1BWP30P140LVT U203 ( .A1(n180), .A2(i_data_bus[245]), .B1(n179), .B2(
        i_data_bus[85]), .ZN(n162) );
  ND4D1BWP30P140LVT U204 ( .A1(n165), .A2(n164), .A3(n163), .A4(n162), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U205 ( .A1(n175), .A2(i_data_bus[148]), .B1(n174), .B2(
        i_data_bus[20]), .ZN(n169) );
  AOI22D1BWP30P140LVT U206 ( .A1(n177), .A2(i_data_bus[52]), .B1(n176), .B2(
        i_data_bus[116]), .ZN(n168) );
  AOI22D1BWP30P140LVT U207 ( .A1(n178), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n167) );
  AOI22D1BWP30P140LVT U208 ( .A1(n180), .A2(i_data_bus[244]), .B1(n179), .B2(
        i_data_bus[84]), .ZN(n166) );
  ND4D1BWP30P140LVT U209 ( .A1(n169), .A2(n168), .A3(n167), .A4(n166), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U210 ( .A1(n175), .A2(i_data_bus[147]), .B1(n174), .B2(
        i_data_bus[19]), .ZN(n173) );
  AOI22D1BWP30P140LVT U211 ( .A1(n177), .A2(i_data_bus[51]), .B1(n176), .B2(
        i_data_bus[115]), .ZN(n172) );
  AOI22D1BWP30P140LVT U212 ( .A1(n178), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n171) );
  AOI22D1BWP30P140LVT U213 ( .A1(n180), .A2(i_data_bus[243]), .B1(n179), .B2(
        i_data_bus[83]), .ZN(n170) );
  ND4D1BWP30P140LVT U214 ( .A1(n173), .A2(n172), .A3(n171), .A4(n170), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U215 ( .A1(n175), .A2(i_data_bus[146]), .B1(n174), .B2(
        i_data_bus[18]), .ZN(n184) );
  AOI22D1BWP30P140LVT U216 ( .A1(n177), .A2(i_data_bus[50]), .B1(n176), .B2(
        i_data_bus[114]), .ZN(n183) );
  AOI22D1BWP30P140LVT U217 ( .A1(n178), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n182) );
  AOI22D1BWP30P140LVT U218 ( .A1(n180), .A2(i_data_bus[242]), .B1(n179), .B2(
        i_data_bus[82]), .ZN(n181) );
  ND4D1BWP30P140LVT U219 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .ZN(
        N387) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_5 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  BUFFD2BWP30P140LVT U3 ( .I(n130), .Z(n183) );
  BUFFD2BWP30P140LVT U4 ( .I(n130), .Z(n155) );
  INVD1BWP30P140LVT U5 ( .I(n36), .ZN(n101) );
  INVD1BWP30P140LVT U6 ( .I(n31), .ZN(n141) );
  INVD3BWP30P140LVT U7 ( .I(n72), .ZN(n156) );
  INVD2BWP30P140LVT U8 ( .I(n18), .ZN(n47) );
  NR2D1BWP30P140LVT U9 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n34) );
  NR4D1BWP30P140LVT U10 ( .A1(n17), .A2(i_cmd[6]), .A3(n16), .A4(n15), .ZN(n18) );
  CKND2D3BWP30P140LVT U11 ( .A1(n22), .A2(n4), .ZN(n32) );
  INVD1BWP30P140LVT U12 ( .I(i_cmd[3]), .ZN(n7) );
  NR2D2BWP30P140LVT U13 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n9) );
  INVD1BWP30P140LVT U14 ( .I(n14), .ZN(n72) );
  INVD8BWP30P140LVT U15 ( .I(n47), .ZN(n2) );
  INVD2BWP30P140LVT U16 ( .I(n101), .ZN(n154) );
  INVD4BWP30P140LVT U17 ( .I(n141), .ZN(n1) );
  INVD3BWP30P140LVT U18 ( .I(n44), .ZN(n184) );
  AOI22D1BWP30P140LVT U19 ( .A1(n156), .A2(i_data_bus[208]), .B1(n2), .B2(
        i_data_bus[176]), .ZN(n19) );
  INR2D2BWP30P140LVT U20 ( .A1(n11), .B1(n32), .ZN(n27) );
  INR2D2BWP30P140LVT U21 ( .A1(n8), .B1(i_cmd[7]), .ZN(n4) );
  INVD1BWP30P140LVT U22 ( .I(i_cmd[5]), .ZN(n16) );
  NR4D1BWP30P140LVT U23 ( .A1(n17), .A2(i_cmd[5]), .A3(n13), .A4(n12), .ZN(n14) );
  INVD1BWP30P140LVT U24 ( .I(i_cmd[4]), .ZN(n35) );
  NR4D0BWP30P140LVT U25 ( .A1(n30), .A2(i_cmd[1]), .A3(n29), .A4(n28), .ZN(n31) );
  INVD1BWP30P140LVT U26 ( .I(i_cmd[2]), .ZN(n29) );
  INVD1BWP30P140LVT U27 ( .I(n131), .ZN(n44) );
  INVD1BWP30P140LVT U28 ( .I(n26), .ZN(n17) );
  INVD1BWP30P140LVT U29 ( .I(n27), .ZN(n30) );
  ND3D1BWP30P140LVT U30 ( .A1(n34), .A2(i_valid[1]), .A3(i_cmd[1]), .ZN(n6) );
  INVD3BWP30P140LVT U31 ( .I(n40), .ZN(n181) );
  INVD1BWP30P140LVT U32 ( .I(n39), .ZN(n40) );
  INVD1BWP30P140LVT U33 ( .I(i_cmd[0]), .ZN(n38) );
  NR2D1BWP30P140LVT U34 ( .A1(n24), .A2(n23), .ZN(n25) );
  ND2D1BWP30P140LVT U35 ( .A1(i_cmd[7]), .A2(i_valid[7]), .ZN(n23) );
  ND2D1BWP30P140LVT U36 ( .A1(n46), .A2(n45), .ZN(N402) );
  AN2D2BWP30P140LVT U37 ( .A1(n26), .A2(n25), .Z(n3) );
  INR2D2BWP30P140LVT U38 ( .A1(n27), .B1(n5), .ZN(n130) );
  NR2D3BWP30P140LVT U39 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n11) );
  NR2OPTPAD4BWP30P140LVT U40 ( .A1(i_cmd[5]), .A2(i_cmd[6]), .ZN(n22) );
  INR2D1BWP30P140LVT U41 ( .A1(i_en), .B1(rst), .ZN(n8) );
  ND3D1BWP30P140LVT U42 ( .A1(i_cmd[3]), .A2(i_valid[3]), .A3(n9), .ZN(n5) );
  INR2D2BWP30P140LVT U43 ( .A1(n27), .B1(n6), .ZN(n131) );
  AOI22D1BWP30P140LVT U44 ( .A1(i_data_bus[112]), .A2(n130), .B1(n131), .B2(
        i_data_bus[48]), .ZN(n21) );
  ND3OPTPAD2BWP30P140LVT U45 ( .A1(n9), .A2(n8), .A3(n7), .ZN(n10) );
  INR2D2BWP30P140LVT U46 ( .A1(n11), .B1(n10), .ZN(n26) );
  IND2D1BWP30P140LVT U47 ( .A1(i_cmd[7]), .B1(i_valid[6]), .ZN(n13) );
  INVD1BWP30P140LVT U48 ( .I(i_cmd[6]), .ZN(n12) );
  IND2D1BWP30P140LVT U49 ( .A1(i_cmd[7]), .B1(i_valid[5]), .ZN(n15) );
  INVD1BWP30P140LVT U50 ( .I(n19), .ZN(n20) );
  INR2D1BWP30P140LVT U51 ( .A1(n21), .B1(n20), .ZN(n43) );
  INVD1BWP30P140LVT U52 ( .I(n22), .ZN(n24) );
  IND2D1BWP30P140LVT U53 ( .A1(i_cmd[3]), .B1(i_valid[2]), .ZN(n28) );
  AOI22D1BWP30P140LVT U54 ( .A1(n3), .A2(i_data_bus[240]), .B1(n1), .B2(
        i_data_bus[80]), .ZN(n42) );
  INVD2BWP30P140LVT U55 ( .I(n32), .ZN(n33) );
  IND3D4BWP30P140LVT U56 ( .A1(i_cmd[1]), .B1(n34), .B2(n33), .ZN(n37) );
  INR4D1BWP30P140LVT U57 ( .A1(i_valid[4]), .B1(i_cmd[0]), .B2(n35), .B3(n37), 
        .ZN(n36) );
  INVD2BWP30P140LVT U58 ( .I(n101), .ZN(n182) );
  INR4D1BWP30P140LVT U59 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n38), .B3(n37), 
        .ZN(n39) );
  AOI22D1BWP30P140LVT U60 ( .A1(n182), .A2(i_data_bus[144]), .B1(n181), .B2(
        i_data_bus[16]), .ZN(n41) );
  ND3D1BWP30P140LVT U61 ( .A1(n43), .A2(n42), .A3(n41), .ZN(N385) );
  NR4D0BWP30P140LVT U62 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .ZN(n46)
         );
  INVD2BWP30P140LVT U63 ( .I(n72), .ZN(n185) );
  NR4D0BWP30P140LVT U64 ( .A1(n3), .A2(n185), .A3(n1), .A4(n2), .ZN(n45) );
  AOI22D1BWP30P140LVT U65 ( .A1(n154), .A2(i_data_bus[140]), .B1(n181), .B2(
        i_data_bus[12]), .ZN(n51) );
  AOI22D1BWP30P140LVT U66 ( .A1(n184), .A2(i_data_bus[44]), .B1(n155), .B2(
        i_data_bus[108]), .ZN(n50) );
  AOI22D1BWP30P140LVT U67 ( .A1(n156), .A2(i_data_bus[204]), .B1(n2), .B2(
        i_data_bus[172]), .ZN(n49) );
  AOI22D1BWP30P140LVT U68 ( .A1(n3), .A2(i_data_bus[236]), .B1(n1), .B2(
        i_data_bus[76]), .ZN(n48) );
  ND4D1BWP30P140LVT U69 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(N381) );
  AOI22D1BWP30P140LVT U70 ( .A1(n154), .A2(i_data_bus[139]), .B1(n181), .B2(
        i_data_bus[11]), .ZN(n55) );
  AOI22D1BWP30P140LVT U71 ( .A1(n184), .A2(i_data_bus[43]), .B1(n155), .B2(
        i_data_bus[107]), .ZN(n54) );
  AOI22D1BWP30P140LVT U72 ( .A1(n156), .A2(i_data_bus[203]), .B1(n2), .B2(
        i_data_bus[171]), .ZN(n53) );
  AOI22D1BWP30P140LVT U73 ( .A1(n3), .A2(i_data_bus[235]), .B1(n1), .B2(
        i_data_bus[75]), .ZN(n52) );
  ND4D1BWP30P140LVT U74 ( .A1(n55), .A2(n54), .A3(n53), .A4(n52), .ZN(N380) );
  AOI22D1BWP30P140LVT U75 ( .A1(n154), .A2(i_data_bus[136]), .B1(n181), .B2(
        i_data_bus[8]), .ZN(n59) );
  AOI22D1BWP30P140LVT U76 ( .A1(n184), .A2(i_data_bus[40]), .B1(n155), .B2(
        i_data_bus[104]), .ZN(n58) );
  AOI22D1BWP30P140LVT U77 ( .A1(n156), .A2(i_data_bus[200]), .B1(n2), .B2(
        i_data_bus[168]), .ZN(n57) );
  AOI22D1BWP30P140LVT U78 ( .A1(n3), .A2(i_data_bus[232]), .B1(n1), .B2(
        i_data_bus[72]), .ZN(n56) );
  ND4D1BWP30P140LVT U79 ( .A1(n59), .A2(n58), .A3(n57), .A4(n56), .ZN(N377) );
  AOI22D1BWP30P140LVT U80 ( .A1(n154), .A2(i_data_bus[134]), .B1(n181), .B2(
        i_data_bus[6]), .ZN(n63) );
  AOI22D1BWP30P140LVT U81 ( .A1(n184), .A2(i_data_bus[38]), .B1(n155), .B2(
        i_data_bus[102]), .ZN(n62) );
  AOI22D1BWP30P140LVT U82 ( .A1(n156), .A2(i_data_bus[198]), .B1(n2), .B2(
        i_data_bus[166]), .ZN(n61) );
  AOI22D1BWP30P140LVT U83 ( .A1(n3), .A2(i_data_bus[230]), .B1(n1), .B2(
        i_data_bus[70]), .ZN(n60) );
  ND4D1BWP30P140LVT U84 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .ZN(N375) );
  AOI22D1BWP30P140LVT U85 ( .A1(n154), .A2(i_data_bus[133]), .B1(n181), .B2(
        i_data_bus[5]), .ZN(n67) );
  AOI22D1BWP30P140LVT U86 ( .A1(n184), .A2(i_data_bus[37]), .B1(n155), .B2(
        i_data_bus[101]), .ZN(n66) );
  AOI22D1BWP30P140LVT U87 ( .A1(n156), .A2(i_data_bus[197]), .B1(n2), .B2(
        i_data_bus[165]), .ZN(n65) );
  AOI22D1BWP30P140LVT U88 ( .A1(n3), .A2(i_data_bus[229]), .B1(n1), .B2(
        i_data_bus[69]), .ZN(n64) );
  ND4D1BWP30P140LVT U89 ( .A1(n67), .A2(n66), .A3(n65), .A4(n64), .ZN(N374) );
  AOI22D1BWP30P140LVT U90 ( .A1(n154), .A2(i_data_bus[130]), .B1(n181), .B2(
        i_data_bus[2]), .ZN(n71) );
  AOI22D1BWP30P140LVT U91 ( .A1(n184), .A2(i_data_bus[34]), .B1(n155), .B2(
        i_data_bus[98]), .ZN(n70) );
  AOI22D1BWP30P140LVT U92 ( .A1(n156), .A2(i_data_bus[194]), .B1(n2), .B2(
        i_data_bus[162]), .ZN(n69) );
  AOI22D1BWP30P140LVT U93 ( .A1(n3), .A2(i_data_bus[226]), .B1(n1), .B2(
        i_data_bus[66]), .ZN(n68) );
  ND4D1BWP30P140LVT U94 ( .A1(n71), .A2(n70), .A3(n69), .A4(n68), .ZN(N371) );
  AOI22D1BWP30P140LVT U95 ( .A1(n154), .A2(i_data_bus[128]), .B1(n181), .B2(
        i_data_bus[0]), .ZN(n76) );
  AOI22D1BWP30P140LVT U96 ( .A1(n184), .A2(i_data_bus[32]), .B1(n155), .B2(
        i_data_bus[96]), .ZN(n75) );
  AOI22D1BWP30P140LVT U97 ( .A1(n185), .A2(i_data_bus[192]), .B1(n2), .B2(
        i_data_bus[160]), .ZN(n74) );
  AOI22D1BWP30P140LVT U98 ( .A1(n3), .A2(i_data_bus[224]), .B1(n1), .B2(
        i_data_bus[64]), .ZN(n73) );
  ND4D1BWP30P140LVT U99 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(N369) );
  AOI22D1BWP30P140LVT U100 ( .A1(n154), .A2(i_data_bus[138]), .B1(n181), .B2(
        i_data_bus[10]), .ZN(n80) );
  AOI22D1BWP30P140LVT U101 ( .A1(n131), .A2(i_data_bus[42]), .B1(n130), .B2(
        i_data_bus[106]), .ZN(n79) );
  AOI22D1BWP30P140LVT U102 ( .A1(n156), .A2(i_data_bus[202]), .B1(n2), .B2(
        i_data_bus[170]), .ZN(n78) );
  AOI22D1BWP30P140LVT U103 ( .A1(n3), .A2(i_data_bus[234]), .B1(n1), .B2(
        i_data_bus[74]), .ZN(n77) );
  ND4D1BWP30P140LVT U104 ( .A1(n80), .A2(n79), .A3(n78), .A4(n77), .ZN(N379)
         );
  AOI22D1BWP30P140LVT U105 ( .A1(n154), .A2(i_data_bus[137]), .B1(n181), .B2(
        i_data_bus[9]), .ZN(n84) );
  AOI22D1BWP30P140LVT U106 ( .A1(n131), .A2(i_data_bus[41]), .B1(n130), .B2(
        i_data_bus[105]), .ZN(n83) );
  AOI22D1BWP30P140LVT U107 ( .A1(n156), .A2(i_data_bus[201]), .B1(n2), .B2(
        i_data_bus[169]), .ZN(n82) );
  AOI22D1BWP30P140LVT U108 ( .A1(n3), .A2(i_data_bus[233]), .B1(n1), .B2(
        i_data_bus[73]), .ZN(n81) );
  ND4D1BWP30P140LVT U109 ( .A1(n84), .A2(n83), .A3(n82), .A4(n81), .ZN(N378)
         );
  INVD1BWP30P140LVT U110 ( .I(i_data_bus[135]), .ZN(n85) );
  MAOI22D1BWP30P140LVT U111 ( .A1(n181), .A2(i_data_bus[7]), .B1(n101), .B2(
        n85), .ZN(n89) );
  AOI22D1BWP30P140LVT U112 ( .A1(n131), .A2(i_data_bus[39]), .B1(n130), .B2(
        i_data_bus[103]), .ZN(n88) );
  AOI22D1BWP30P140LVT U113 ( .A1(n156), .A2(i_data_bus[199]), .B1(n2), .B2(
        i_data_bus[167]), .ZN(n87) );
  AOI22D1BWP30P140LVT U114 ( .A1(n3), .A2(i_data_bus[231]), .B1(n1), .B2(
        i_data_bus[71]), .ZN(n86) );
  ND4D1BWP30P140LVT U115 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(N376)
         );
  INVD1BWP30P140LVT U116 ( .I(i_data_bus[132]), .ZN(n90) );
  MAOI22D1BWP30P140LVT U117 ( .A1(n181), .A2(i_data_bus[4]), .B1(n101), .B2(
        n90), .ZN(n94) );
  AOI22D1BWP30P140LVT U118 ( .A1(n184), .A2(i_data_bus[36]), .B1(n155), .B2(
        i_data_bus[100]), .ZN(n93) );
  AOI22D1BWP30P140LVT U119 ( .A1(n156), .A2(i_data_bus[196]), .B1(n2), .B2(
        i_data_bus[164]), .ZN(n92) );
  AOI22D1BWP30P140LVT U120 ( .A1(n3), .A2(i_data_bus[228]), .B1(n1), .B2(
        i_data_bus[68]), .ZN(n91) );
  ND4D1BWP30P140LVT U121 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .ZN(N373)
         );
  INVD1BWP30P140LVT U122 ( .I(i_data_bus[131]), .ZN(n95) );
  MAOI22D1BWP30P140LVT U123 ( .A1(n181), .A2(i_data_bus[3]), .B1(n101), .B2(
        n95), .ZN(n99) );
  AOI22D1BWP30P140LVT U124 ( .A1(n131), .A2(i_data_bus[35]), .B1(n130), .B2(
        i_data_bus[99]), .ZN(n98) );
  AOI22D1BWP30P140LVT U125 ( .A1(n156), .A2(i_data_bus[195]), .B1(n2), .B2(
        i_data_bus[163]), .ZN(n97) );
  AOI22D1BWP30P140LVT U126 ( .A1(n3), .A2(i_data_bus[227]), .B1(n1), .B2(
        i_data_bus[67]), .ZN(n96) );
  ND4D1BWP30P140LVT U127 ( .A1(n99), .A2(n98), .A3(n97), .A4(n96), .ZN(N372)
         );
  INVD1BWP30P140LVT U128 ( .I(i_data_bus[129]), .ZN(n100) );
  MAOI22D1BWP30P140LVT U129 ( .A1(n181), .A2(i_data_bus[1]), .B1(n101), .B2(
        n100), .ZN(n105) );
  AOI22D1BWP30P140LVT U130 ( .A1(n184), .A2(i_data_bus[33]), .B1(n155), .B2(
        i_data_bus[97]), .ZN(n104) );
  AOI22D1BWP30P140LVT U131 ( .A1(n156), .A2(i_data_bus[193]), .B1(n2), .B2(
        i_data_bus[161]), .ZN(n103) );
  AOI22D1BWP30P140LVT U132 ( .A1(n3), .A2(i_data_bus[225]), .B1(n1), .B2(
        i_data_bus[65]), .ZN(n102) );
  ND4D1BWP30P140LVT U133 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .ZN(
        N370) );
  AOI22D1BWP30P140LVT U134 ( .A1(n182), .A2(i_data_bus[159]), .B1(n181), .B2(
        i_data_bus[31]), .ZN(n109) );
  AOI22D1BWP30P140LVT U135 ( .A1(n131), .A2(i_data_bus[63]), .B1(n130), .B2(
        i_data_bus[127]), .ZN(n108) );
  AOI22D1BWP30P140LVT U136 ( .A1(n185), .A2(i_data_bus[223]), .B1(n2), .B2(
        i_data_bus[191]), .ZN(n107) );
  AOI22D1BWP30P140LVT U137 ( .A1(n3), .A2(i_data_bus[255]), .B1(n1), .B2(
        i_data_bus[95]), .ZN(n106) );
  ND4D1BWP30P140LVT U138 ( .A1(n109), .A2(n108), .A3(n107), .A4(n106), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U139 ( .A1(n182), .A2(i_data_bus[158]), .B1(n181), .B2(
        i_data_bus[30]), .ZN(n113) );
  AOI22D1BWP30P140LVT U140 ( .A1(n184), .A2(i_data_bus[62]), .B1(n183), .B2(
        i_data_bus[126]), .ZN(n112) );
  AOI22D1BWP30P140LVT U141 ( .A1(n185), .A2(i_data_bus[222]), .B1(n2), .B2(
        i_data_bus[190]), .ZN(n111) );
  AOI22D1BWP30P140LVT U142 ( .A1(n3), .A2(i_data_bus[254]), .B1(n1), .B2(
        i_data_bus[94]), .ZN(n110) );
  ND4D1BWP30P140LVT U143 ( .A1(n113), .A2(n112), .A3(n111), .A4(n110), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U144 ( .A1(n182), .A2(i_data_bus[156]), .B1(n181), .B2(
        i_data_bus[28]), .ZN(n117) );
  AOI22D1BWP30P140LVT U145 ( .A1(n184), .A2(i_data_bus[60]), .B1(n183), .B2(
        i_data_bus[124]), .ZN(n116) );
  AOI22D1BWP30P140LVT U146 ( .A1(n185), .A2(i_data_bus[220]), .B1(n2), .B2(
        i_data_bus[188]), .ZN(n115) );
  AOI22D1BWP30P140LVT U147 ( .A1(n3), .A2(i_data_bus[252]), .B1(n1), .B2(
        i_data_bus[92]), .ZN(n114) );
  ND4D1BWP30P140LVT U148 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U149 ( .A1(n182), .A2(i_data_bus[155]), .B1(n181), .B2(
        i_data_bus[27]), .ZN(n121) );
  AOI22D1BWP30P140LVT U150 ( .A1(n131), .A2(i_data_bus[59]), .B1(n130), .B2(
        i_data_bus[123]), .ZN(n120) );
  AOI22D1BWP30P140LVT U151 ( .A1(n185), .A2(i_data_bus[219]), .B1(n2), .B2(
        i_data_bus[187]), .ZN(n119) );
  AOI22D1BWP30P140LVT U152 ( .A1(n3), .A2(i_data_bus[251]), .B1(n1), .B2(
        i_data_bus[91]), .ZN(n118) );
  ND4D1BWP30P140LVT U153 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U154 ( .A1(n182), .A2(i_data_bus[153]), .B1(n181), .B2(
        i_data_bus[25]), .ZN(n125) );
  AOI22D1BWP30P140LVT U155 ( .A1(n184), .A2(i_data_bus[57]), .B1(n183), .B2(
        i_data_bus[121]), .ZN(n124) );
  AOI22D1BWP30P140LVT U156 ( .A1(n185), .A2(i_data_bus[217]), .B1(n2), .B2(
        i_data_bus[185]), .ZN(n123) );
  AOI22D1BWP30P140LVT U157 ( .A1(n3), .A2(i_data_bus[249]), .B1(n1), .B2(
        i_data_bus[89]), .ZN(n122) );
  ND4D1BWP30P140LVT U158 ( .A1(n125), .A2(n124), .A3(n123), .A4(n122), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U159 ( .A1(n182), .A2(i_data_bus[152]), .B1(n181), .B2(
        i_data_bus[24]), .ZN(n129) );
  AOI22D1BWP30P140LVT U160 ( .A1(n184), .A2(i_data_bus[56]), .B1(n183), .B2(
        i_data_bus[120]), .ZN(n128) );
  AOI22D1BWP30P140LVT U161 ( .A1(n185), .A2(i_data_bus[216]), .B1(n2), .B2(
        i_data_bus[184]), .ZN(n127) );
  AOI22D1BWP30P140LVT U162 ( .A1(n3), .A2(i_data_bus[248]), .B1(n1), .B2(
        i_data_bus[88]), .ZN(n126) );
  ND4D1BWP30P140LVT U163 ( .A1(n129), .A2(n128), .A3(n127), .A4(n126), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U164 ( .A1(n154), .A2(i_data_bus[143]), .B1(n181), .B2(
        i_data_bus[15]), .ZN(n135) );
  AOI22D1BWP30P140LVT U165 ( .A1(n131), .A2(i_data_bus[47]), .B1(n130), .B2(
        i_data_bus[111]), .ZN(n134) );
  AOI22D1BWP30P140LVT U166 ( .A1(n156), .A2(i_data_bus[207]), .B1(n2), .B2(
        i_data_bus[175]), .ZN(n133) );
  AOI22D1BWP30P140LVT U167 ( .A1(n3), .A2(i_data_bus[239]), .B1(n1), .B2(
        i_data_bus[79]), .ZN(n132) );
  ND4D1BWP30P140LVT U168 ( .A1(n135), .A2(n134), .A3(n133), .A4(n132), .ZN(
        N384) );
  AOI22D1BWP30P140LVT U169 ( .A1(n154), .A2(i_data_bus[141]), .B1(n181), .B2(
        i_data_bus[13]), .ZN(n139) );
  AOI22D1BWP30P140LVT U170 ( .A1(n184), .A2(i_data_bus[45]), .B1(n155), .B2(
        i_data_bus[109]), .ZN(n138) );
  AOI22D1BWP30P140LVT U171 ( .A1(n156), .A2(i_data_bus[205]), .B1(n2), .B2(
        i_data_bus[173]), .ZN(n137) );
  AOI22D1BWP30P140LVT U172 ( .A1(n3), .A2(i_data_bus[237]), .B1(n1), .B2(
        i_data_bus[77]), .ZN(n136) );
  ND4D1BWP30P140LVT U173 ( .A1(n139), .A2(n138), .A3(n137), .A4(n136), .ZN(
        N382) );
  AOI22D1BWP30P140LVT U174 ( .A1(n182), .A2(i_data_bus[157]), .B1(n181), .B2(
        i_data_bus[29]), .ZN(n145) );
  AOI22D1BWP30P140LVT U175 ( .A1(n184), .A2(i_data_bus[61]), .B1(n183), .B2(
        i_data_bus[125]), .ZN(n144) );
  AOI22D1BWP30P140LVT U176 ( .A1(n185), .A2(i_data_bus[221]), .B1(n2), .B2(
        i_data_bus[189]), .ZN(n143) );
  INVD1BWP30P140LVT U177 ( .I(i_data_bus[93]), .ZN(n140) );
  MAOI22D1BWP30P140LVT U178 ( .A1(n3), .A2(i_data_bus[253]), .B1(n141), .B2(
        n140), .ZN(n142) );
  ND4D1BWP30P140LVT U179 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U180 ( .A1(n182), .A2(i_data_bus[154]), .B1(n181), .B2(
        i_data_bus[26]), .ZN(n149) );
  AOI22D1BWP30P140LVT U181 ( .A1(n184), .A2(i_data_bus[58]), .B1(n155), .B2(
        i_data_bus[122]), .ZN(n148) );
  AOI22D1BWP30P140LVT U182 ( .A1(n185), .A2(i_data_bus[218]), .B1(n2), .B2(
        i_data_bus[186]), .ZN(n147) );
  AOI22D1BWP30P140LVT U183 ( .A1(n3), .A2(i_data_bus[250]), .B1(n1), .B2(
        i_data_bus[90]), .ZN(n146) );
  ND4D1BWP30P140LVT U184 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U185 ( .A1(n182), .A2(i_data_bus[151]), .B1(n181), .B2(
        i_data_bus[23]), .ZN(n153) );
  AOI22D1BWP30P140LVT U186 ( .A1(n184), .A2(i_data_bus[55]), .B1(n183), .B2(
        i_data_bus[119]), .ZN(n152) );
  AOI22D1BWP30P140LVT U187 ( .A1(n185), .A2(i_data_bus[215]), .B1(n2), .B2(
        i_data_bus[183]), .ZN(n151) );
  AOI22D1BWP30P140LVT U188 ( .A1(n3), .A2(i_data_bus[247]), .B1(n1), .B2(
        i_data_bus[87]), .ZN(n150) );
  ND4D1BWP30P140LVT U189 ( .A1(n153), .A2(n152), .A3(n151), .A4(n150), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U190 ( .A1(n154), .A2(i_data_bus[142]), .B1(n181), .B2(
        i_data_bus[14]), .ZN(n160) );
  AOI22D1BWP30P140LVT U191 ( .A1(n184), .A2(i_data_bus[46]), .B1(n155), .B2(
        i_data_bus[110]), .ZN(n159) );
  AOI22D1BWP30P140LVT U192 ( .A1(n156), .A2(i_data_bus[206]), .B1(n2), .B2(
        i_data_bus[174]), .ZN(n158) );
  AOI22D1BWP30P140LVT U193 ( .A1(n3), .A2(i_data_bus[238]), .B1(n1), .B2(
        i_data_bus[78]), .ZN(n157) );
  ND4D1BWP30P140LVT U194 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(
        N383) );
  AOI22D1BWP30P140LVT U195 ( .A1(n182), .A2(i_data_bus[150]), .B1(n181), .B2(
        i_data_bus[22]), .ZN(n164) );
  AOI22D1BWP30P140LVT U196 ( .A1(n184), .A2(i_data_bus[54]), .B1(n183), .B2(
        i_data_bus[118]), .ZN(n163) );
  AOI22D1BWP30P140LVT U197 ( .A1(n185), .A2(i_data_bus[214]), .B1(n2), .B2(
        i_data_bus[182]), .ZN(n162) );
  AOI22D1BWP30P140LVT U198 ( .A1(n3), .A2(i_data_bus[246]), .B1(n1), .B2(
        i_data_bus[86]), .ZN(n161) );
  ND4D1BWP30P140LVT U199 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U200 ( .A1(n182), .A2(i_data_bus[149]), .B1(n181), .B2(
        i_data_bus[21]), .ZN(n168) );
  AOI22D1BWP30P140LVT U201 ( .A1(n184), .A2(i_data_bus[53]), .B1(n183), .B2(
        i_data_bus[117]), .ZN(n167) );
  AOI22D1BWP30P140LVT U202 ( .A1(n185), .A2(i_data_bus[213]), .B1(n2), .B2(
        i_data_bus[181]), .ZN(n166) );
  AOI22D1BWP30P140LVT U203 ( .A1(n3), .A2(i_data_bus[245]), .B1(n1), .B2(
        i_data_bus[85]), .ZN(n165) );
  ND4D1BWP30P140LVT U204 ( .A1(n168), .A2(n167), .A3(n166), .A4(n165), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U205 ( .A1(n182), .A2(i_data_bus[148]), .B1(n181), .B2(
        i_data_bus[20]), .ZN(n172) );
  AOI22D1BWP30P140LVT U206 ( .A1(n184), .A2(i_data_bus[52]), .B1(n183), .B2(
        i_data_bus[116]), .ZN(n171) );
  AOI22D1BWP30P140LVT U207 ( .A1(n185), .A2(i_data_bus[212]), .B1(n2), .B2(
        i_data_bus[180]), .ZN(n170) );
  AOI22D1BWP30P140LVT U208 ( .A1(n3), .A2(i_data_bus[244]), .B1(n1), .B2(
        i_data_bus[84]), .ZN(n169) );
  ND4D1BWP30P140LVT U209 ( .A1(n172), .A2(n171), .A3(n170), .A4(n169), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U210 ( .A1(n182), .A2(i_data_bus[147]), .B1(n181), .B2(
        i_data_bus[19]), .ZN(n176) );
  AOI22D1BWP30P140LVT U211 ( .A1(n184), .A2(i_data_bus[51]), .B1(n183), .B2(
        i_data_bus[115]), .ZN(n175) );
  AOI22D1BWP30P140LVT U212 ( .A1(n185), .A2(i_data_bus[211]), .B1(n2), .B2(
        i_data_bus[179]), .ZN(n174) );
  AOI22D1BWP30P140LVT U213 ( .A1(n3), .A2(i_data_bus[243]), .B1(n1), .B2(
        i_data_bus[83]), .ZN(n173) );
  ND4D1BWP30P140LVT U214 ( .A1(n176), .A2(n175), .A3(n174), .A4(n173), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U215 ( .A1(n182), .A2(i_data_bus[146]), .B1(n181), .B2(
        i_data_bus[18]), .ZN(n180) );
  AOI22D1BWP30P140LVT U216 ( .A1(n184), .A2(i_data_bus[50]), .B1(n183), .B2(
        i_data_bus[114]), .ZN(n179) );
  AOI22D1BWP30P140LVT U217 ( .A1(n185), .A2(i_data_bus[210]), .B1(n2), .B2(
        i_data_bus[178]), .ZN(n178) );
  AOI22D1BWP30P140LVT U218 ( .A1(n3), .A2(i_data_bus[242]), .B1(n1), .B2(
        i_data_bus[82]), .ZN(n177) );
  ND4D1BWP30P140LVT U219 ( .A1(n180), .A2(n179), .A3(n178), .A4(n177), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U220 ( .A1(n182), .A2(i_data_bus[145]), .B1(n181), .B2(
        i_data_bus[17]), .ZN(n189) );
  AOI22D1BWP30P140LVT U221 ( .A1(n184), .A2(i_data_bus[49]), .B1(n183), .B2(
        i_data_bus[113]), .ZN(n188) );
  AOI22D1BWP30P140LVT U222 ( .A1(n185), .A2(i_data_bus[209]), .B1(n2), .B2(
        i_data_bus[177]), .ZN(n187) );
  AOI22D1BWP30P140LVT U223 ( .A1(n3), .A2(i_data_bus[241]), .B1(n1), .B2(
        i_data_bus[81]), .ZN(n186) );
  ND4D1BWP30P140LVT U224 ( .A1(n189), .A2(n188), .A3(n187), .A4(n186), .ZN(
        N386) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_6 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD1BWP30P140LVT U3 ( .I(n15), .ZN(n16) );
  INVD1BWP30P140LVT U4 ( .I(n37), .ZN(n40) );
  NR4D1BWP30P140LVT U5 ( .A1(n36), .A2(i_cmd[6]), .A3(n35), .A4(n34), .ZN(n37)
         );
  NR2D1BWP30P140LVT U6 ( .A1(i_cmd[7]), .A2(i_cmd[5]), .ZN(n3) );
  INR2D1BWP30P140LVT U7 ( .A1(n18), .B1(i_cmd[6]), .ZN(n2) );
  INVD1BWP30P140LVT U8 ( .I(n28), .ZN(n90) );
  INVD6BWP30P140LVT U9 ( .I(n40), .ZN(n1) );
  INVD6BWP30P140LVT U10 ( .I(n16), .ZN(n177) );
  NR2OPTPAD2BWP30P140LVT U11 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n19) );
  INVD1BWP30P140LVT U12 ( .I(i_cmd[2]), .ZN(n31) );
  INVD1BWP30P140LVT U13 ( .I(i_cmd[6]), .ZN(n26) );
  INVD2BWP30P140LVT U14 ( .I(n29), .ZN(n32) );
  IND3D2BWP30P140LVT U15 ( .A1(i_cmd[1]), .B1(n10), .B2(n9), .ZN(n13) );
  INVD2BWP30P140LVT U16 ( .I(n8), .ZN(n9) );
  INVD1BWP30P140LVT U17 ( .I(i_cmd[5]), .ZN(n35) );
  NR2D2BWP30P140LVT U18 ( .A1(n4), .A2(n8), .ZN(n29) );
  INVD1BWP30P140LVT U19 ( .I(n21), .ZN(n4) );
  INVD2BWP30P140LVT U20 ( .I(n12), .ZN(n176) );
  INVD1BWP30P140LVT U21 ( .I(i_cmd[4]), .ZN(n11) );
  INVD2BWP30P140LVT U22 ( .I(n176), .ZN(n147) );
  INVD2BWP30P140LVT U23 ( .I(n176), .ZN(n157) );
  BUFFD4BWP30P140LVT U24 ( .I(n24), .Z(n181) );
  BUFFD4BWP30P140LVT U25 ( .I(n6), .Z(n178) );
  ND2D1BWP30P140LVT U26 ( .A1(n39), .A2(n38), .ZN(N402) );
  NR4D1BWP30P140LVT U27 ( .A1(n32), .A2(i_cmd[1]), .A3(n31), .A4(n30), .ZN(n33) );
  INVD1BWP30P140LVT U28 ( .I(i_cmd[0]), .ZN(n14) );
  NR2OPTPAD1BWP30P140LVT U29 ( .A1(i_cmd[4]), .A2(i_cmd[0]), .ZN(n21) );
  INR2D1BWP30P140LVT U30 ( .A1(i_en), .B1(rst), .ZN(n18) );
  ND2OPTIBD2BWP30P140LVT U31 ( .A1(n3), .A2(n2), .ZN(n8) );
  NR2OPTPAD1BWP30P140LVT U32 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n10) );
  ND3D1BWP30P140LVT U33 ( .A1(i_cmd[1]), .A2(i_valid[1]), .A3(n10), .ZN(n5) );
  INR2D1BWP30P140LVT U34 ( .A1(n29), .B1(n5), .ZN(n6) );
  ND3D1BWP30P140LVT U35 ( .A1(n19), .A2(i_valid[3]), .A3(i_cmd[3]), .ZN(n7) );
  INR2D4BWP30P140LVT U36 ( .A1(n29), .B1(n7), .ZN(n164) );
  INR4D1BWP30P140LVT U37 ( .A1(i_valid[4]), .B1(i_cmd[0]), .B2(n11), .B3(n13), 
        .ZN(n12) );
  INR4D1BWP30P140LVT U38 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n14), .B3(n13), 
        .ZN(n15) );
  NR4D0BWP30P140LVT U39 ( .A1(n178), .A2(n164), .A3(n147), .A4(n177), .ZN(n39)
         );
  INVD2BWP30P140LVT U40 ( .I(i_cmd[3]), .ZN(n17) );
  ND3OPTPAD2BWP30P140LVT U41 ( .A1(n19), .A2(n18), .A3(n17), .ZN(n20) );
  INR2D2BWP30P140LVT U42 ( .A1(n21), .B1(n20), .ZN(n25) );
  NR2D1BWP30P140LVT U43 ( .A1(i_cmd[6]), .A2(i_cmd[5]), .ZN(n22) );
  ND3D1BWP30P140LVT U44 ( .A1(n22), .A2(i_valid[7]), .A3(i_cmd[7]), .ZN(n23)
         );
  INR2D1BWP30P140LVT U45 ( .A1(n25), .B1(n23), .ZN(n24) );
  INVD2BWP30P140LVT U46 ( .I(n25), .ZN(n36) );
  IND2D1BWP30P140LVT U47 ( .A1(i_cmd[7]), .B1(i_valid[6]), .ZN(n27) );
  NR4D1BWP30P140LVT U48 ( .A1(n36), .A2(i_cmd[5]), .A3(n27), .A4(n26), .ZN(n28) );
  INVD2BWP30P140LVT U49 ( .I(n90), .ZN(n170) );
  IND2D1BWP30P140LVT U50 ( .A1(i_cmd[3]), .B1(i_valid[2]), .ZN(n30) );
  INVD2BWP30P140LVT U51 ( .I(n33), .ZN(n41) );
  INVD2BWP30P140LVT U52 ( .I(n41), .ZN(n180) );
  IND2D1BWP30P140LVT U53 ( .A1(i_cmd[7]), .B1(i_valid[5]), .ZN(n34) );
  NR4D0BWP30P140LVT U54 ( .A1(n181), .A2(n170), .A3(n180), .A4(n1), .ZN(n38)
         );
  AOI22D1BWP30P140LVT U55 ( .A1(n157), .A2(i_data_bus[140]), .B1(n177), .B2(
        i_data_bus[12]), .ZN(n45) );
  AOI22D1BWP30P140LVT U56 ( .A1(n178), .A2(i_data_bus[44]), .B1(n164), .B2(
        i_data_bus[108]), .ZN(n44) );
  INVD2BWP30P140LVT U57 ( .I(n90), .ZN(n179) );
  AOI22D1BWP30P140LVT U58 ( .A1(n179), .A2(i_data_bus[204]), .B1(n1), .B2(
        i_data_bus[172]), .ZN(n43) );
  INVD2BWP30P140LVT U59 ( .I(n41), .ZN(n158) );
  AOI22D1BWP30P140LVT U60 ( .A1(n181), .A2(i_data_bus[236]), .B1(n158), .B2(
        i_data_bus[76]), .ZN(n42) );
  ND4D1BWP30P140LVT U61 ( .A1(n45), .A2(n44), .A3(n43), .A4(n42), .ZN(N381) );
  AOI22D1BWP30P140LVT U62 ( .A1(n157), .A2(i_data_bus[139]), .B1(n177), .B2(
        i_data_bus[11]), .ZN(n49) );
  AOI22D1BWP30P140LVT U63 ( .A1(n178), .A2(i_data_bus[43]), .B1(n164), .B2(
        i_data_bus[107]), .ZN(n48) );
  AOI22D1BWP30P140LVT U64 ( .A1(n179), .A2(i_data_bus[203]), .B1(n1), .B2(
        i_data_bus[171]), .ZN(n47) );
  AOI22D1BWP30P140LVT U65 ( .A1(n181), .A2(i_data_bus[235]), .B1(n158), .B2(
        i_data_bus[75]), .ZN(n46) );
  ND4D1BWP30P140LVT U66 ( .A1(n49), .A2(n48), .A3(n47), .A4(n46), .ZN(N380) );
  AOI22D1BWP30P140LVT U67 ( .A1(n157), .A2(i_data_bus[138]), .B1(n177), .B2(
        i_data_bus[10]), .ZN(n53) );
  AOI22D1BWP30P140LVT U68 ( .A1(n178), .A2(i_data_bus[42]), .B1(n164), .B2(
        i_data_bus[106]), .ZN(n52) );
  AOI22D1BWP30P140LVT U69 ( .A1(n179), .A2(i_data_bus[202]), .B1(n1), .B2(
        i_data_bus[170]), .ZN(n51) );
  AOI22D1BWP30P140LVT U70 ( .A1(n181), .A2(i_data_bus[234]), .B1(n158), .B2(
        i_data_bus[74]), .ZN(n50) );
  ND4D1BWP30P140LVT U71 ( .A1(n53), .A2(n52), .A3(n51), .A4(n50), .ZN(N379) );
  AOI22D1BWP30P140LVT U72 ( .A1(n157), .A2(i_data_bus[137]), .B1(n177), .B2(
        i_data_bus[9]), .ZN(n57) );
  AOI22D1BWP30P140LVT U73 ( .A1(n178), .A2(i_data_bus[41]), .B1(n164), .B2(
        i_data_bus[105]), .ZN(n56) );
  AOI22D1BWP30P140LVT U74 ( .A1(n179), .A2(i_data_bus[201]), .B1(n1), .B2(
        i_data_bus[169]), .ZN(n55) );
  AOI22D1BWP30P140LVT U75 ( .A1(n181), .A2(i_data_bus[233]), .B1(n158), .B2(
        i_data_bus[73]), .ZN(n54) );
  ND4D1BWP30P140LVT U76 ( .A1(n57), .A2(n56), .A3(n55), .A4(n54), .ZN(N378) );
  AOI22D1BWP30P140LVT U77 ( .A1(n157), .A2(i_data_bus[136]), .B1(n177), .B2(
        i_data_bus[8]), .ZN(n61) );
  AOI22D1BWP30P140LVT U78 ( .A1(n178), .A2(i_data_bus[40]), .B1(n164), .B2(
        i_data_bus[104]), .ZN(n60) );
  AOI22D1BWP30P140LVT U79 ( .A1(n179), .A2(i_data_bus[200]), .B1(n1), .B2(
        i_data_bus[168]), .ZN(n59) );
  AOI22D1BWP30P140LVT U80 ( .A1(n181), .A2(i_data_bus[232]), .B1(n158), .B2(
        i_data_bus[72]), .ZN(n58) );
  ND4D1BWP30P140LVT U81 ( .A1(n61), .A2(n60), .A3(n59), .A4(n58), .ZN(N377) );
  AOI22D1BWP30P140LVT U82 ( .A1(n157), .A2(i_data_bus[135]), .B1(n177), .B2(
        i_data_bus[7]), .ZN(n65) );
  AOI22D1BWP30P140LVT U83 ( .A1(n178), .A2(i_data_bus[39]), .B1(n164), .B2(
        i_data_bus[103]), .ZN(n64) );
  AOI22D1BWP30P140LVT U84 ( .A1(n179), .A2(i_data_bus[199]), .B1(n1), .B2(
        i_data_bus[167]), .ZN(n63) );
  AOI22D1BWP30P140LVT U85 ( .A1(n181), .A2(i_data_bus[231]), .B1(n158), .B2(
        i_data_bus[71]), .ZN(n62) );
  ND4D1BWP30P140LVT U86 ( .A1(n65), .A2(n64), .A3(n63), .A4(n62), .ZN(N376) );
  AOI22D1BWP30P140LVT U87 ( .A1(n157), .A2(i_data_bus[134]), .B1(n177), .B2(
        i_data_bus[6]), .ZN(n69) );
  AOI22D1BWP30P140LVT U88 ( .A1(n178), .A2(i_data_bus[38]), .B1(n164), .B2(
        i_data_bus[102]), .ZN(n68) );
  AOI22D1BWP30P140LVT U89 ( .A1(n179), .A2(i_data_bus[198]), .B1(n1), .B2(
        i_data_bus[166]), .ZN(n67) );
  AOI22D1BWP30P140LVT U90 ( .A1(n181), .A2(i_data_bus[230]), .B1(n158), .B2(
        i_data_bus[70]), .ZN(n66) );
  ND4D1BWP30P140LVT U91 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(N375) );
  AOI22D1BWP30P140LVT U92 ( .A1(n157), .A2(i_data_bus[133]), .B1(n177), .B2(
        i_data_bus[5]), .ZN(n73) );
  AOI22D1BWP30P140LVT U93 ( .A1(n178), .A2(i_data_bus[37]), .B1(n164), .B2(
        i_data_bus[101]), .ZN(n72) );
  AOI22D1BWP30P140LVT U94 ( .A1(n179), .A2(i_data_bus[197]), .B1(n1), .B2(
        i_data_bus[165]), .ZN(n71) );
  AOI22D1BWP30P140LVT U95 ( .A1(n181), .A2(i_data_bus[229]), .B1(n158), .B2(
        i_data_bus[69]), .ZN(n70) );
  ND4D1BWP30P140LVT U96 ( .A1(n73), .A2(n72), .A3(n71), .A4(n70), .ZN(N374) );
  AOI22D1BWP30P140LVT U97 ( .A1(n157), .A2(i_data_bus[132]), .B1(n177), .B2(
        i_data_bus[4]), .ZN(n77) );
  AOI22D1BWP30P140LVT U98 ( .A1(n178), .A2(i_data_bus[36]), .B1(n164), .B2(
        i_data_bus[100]), .ZN(n76) );
  AOI22D1BWP30P140LVT U99 ( .A1(n179), .A2(i_data_bus[196]), .B1(n1), .B2(
        i_data_bus[164]), .ZN(n75) );
  AOI22D1BWP30P140LVT U100 ( .A1(n181), .A2(i_data_bus[228]), .B1(n158), .B2(
        i_data_bus[68]), .ZN(n74) );
  ND4D1BWP30P140LVT U101 ( .A1(n77), .A2(n76), .A3(n75), .A4(n74), .ZN(N373)
         );
  AOI22D1BWP30P140LVT U102 ( .A1(n157), .A2(i_data_bus[131]), .B1(n177), .B2(
        i_data_bus[3]), .ZN(n81) );
  AOI22D1BWP30P140LVT U103 ( .A1(n178), .A2(i_data_bus[35]), .B1(n164), .B2(
        i_data_bus[99]), .ZN(n80) );
  AOI22D1BWP30P140LVT U104 ( .A1(n179), .A2(i_data_bus[195]), .B1(n1), .B2(
        i_data_bus[163]), .ZN(n79) );
  AOI22D1BWP30P140LVT U105 ( .A1(n181), .A2(i_data_bus[227]), .B1(n158), .B2(
        i_data_bus[67]), .ZN(n78) );
  ND4D1BWP30P140LVT U106 ( .A1(n81), .A2(n80), .A3(n79), .A4(n78), .ZN(N372)
         );
  AOI22D1BWP30P140LVT U107 ( .A1(n157), .A2(i_data_bus[130]), .B1(n177), .B2(
        i_data_bus[2]), .ZN(n85) );
  AOI22D1BWP30P140LVT U108 ( .A1(n178), .A2(i_data_bus[34]), .B1(n164), .B2(
        i_data_bus[98]), .ZN(n84) );
  AOI22D1BWP30P140LVT U109 ( .A1(n179), .A2(i_data_bus[194]), .B1(n1), .B2(
        i_data_bus[162]), .ZN(n83) );
  AOI22D1BWP30P140LVT U110 ( .A1(n181), .A2(i_data_bus[226]), .B1(n158), .B2(
        i_data_bus[66]), .ZN(n82) );
  ND4D1BWP30P140LVT U111 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U112 ( .A1(n157), .A2(i_data_bus[129]), .B1(n177), .B2(
        i_data_bus[1]), .ZN(n89) );
  AOI22D1BWP30P140LVT U113 ( .A1(n178), .A2(i_data_bus[33]), .B1(n164), .B2(
        i_data_bus[97]), .ZN(n88) );
  AOI22D1BWP30P140LVT U114 ( .A1(n179), .A2(i_data_bus[193]), .B1(n1), .B2(
        i_data_bus[161]), .ZN(n87) );
  AOI22D1BWP30P140LVT U115 ( .A1(n181), .A2(i_data_bus[225]), .B1(n158), .B2(
        i_data_bus[65]), .ZN(n86) );
  ND4D1BWP30P140LVT U116 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(N370)
         );
  AOI22D1BWP30P140LVT U117 ( .A1(n157), .A2(i_data_bus[128]), .B1(n177), .B2(
        i_data_bus[0]), .ZN(n94) );
  AOI22D1BWP30P140LVT U118 ( .A1(n178), .A2(i_data_bus[32]), .B1(n164), .B2(
        i_data_bus[96]), .ZN(n93) );
  AOI22D1BWP30P140LVT U119 ( .A1(n170), .A2(i_data_bus[192]), .B1(n1), .B2(
        i_data_bus[160]), .ZN(n92) );
  AOI22D1BWP30P140LVT U120 ( .A1(n181), .A2(i_data_bus[224]), .B1(n158), .B2(
        i_data_bus[64]), .ZN(n91) );
  ND4D1BWP30P140LVT U121 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .ZN(N369)
         );
  AOI22D1BWP30P140LVT U122 ( .A1(n157), .A2(i_data_bus[143]), .B1(n177), .B2(
        i_data_bus[15]), .ZN(n98) );
  AOI22D1BWP30P140LVT U123 ( .A1(n178), .A2(i_data_bus[47]), .B1(n164), .B2(
        i_data_bus[111]), .ZN(n97) );
  AOI22D1BWP30P140LVT U124 ( .A1(n179), .A2(i_data_bus[207]), .B1(n1), .B2(
        i_data_bus[175]), .ZN(n96) );
  AOI22D1BWP30P140LVT U125 ( .A1(n181), .A2(i_data_bus[239]), .B1(n158), .B2(
        i_data_bus[79]), .ZN(n95) );
  ND4D1BWP30P140LVT U126 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .ZN(N384)
         );
  AOI22D1BWP30P140LVT U127 ( .A1(n157), .A2(i_data_bus[142]), .B1(n177), .B2(
        i_data_bus[14]), .ZN(n102) );
  AOI22D1BWP30P140LVT U128 ( .A1(n178), .A2(i_data_bus[46]), .B1(n164), .B2(
        i_data_bus[110]), .ZN(n101) );
  AOI22D1BWP30P140LVT U129 ( .A1(n179), .A2(i_data_bus[206]), .B1(n1), .B2(
        i_data_bus[174]), .ZN(n100) );
  AOI22D1BWP30P140LVT U130 ( .A1(n181), .A2(i_data_bus[238]), .B1(n158), .B2(
        i_data_bus[78]), .ZN(n99) );
  ND4D1BWP30P140LVT U131 ( .A1(n102), .A2(n101), .A3(n100), .A4(n99), .ZN(N383) );
  AOI22D1BWP30P140LVT U132 ( .A1(n147), .A2(i_data_bus[159]), .B1(n177), .B2(
        i_data_bus[31]), .ZN(n106) );
  AOI22D1BWP30P140LVT U133 ( .A1(n178), .A2(i_data_bus[63]), .B1(n164), .B2(
        i_data_bus[127]), .ZN(n105) );
  AOI22D1BWP30P140LVT U134 ( .A1(n170), .A2(i_data_bus[223]), .B1(n1), .B2(
        i_data_bus[191]), .ZN(n104) );
  AOI22D1BWP30P140LVT U135 ( .A1(n181), .A2(i_data_bus[255]), .B1(n180), .B2(
        i_data_bus[95]), .ZN(n103) );
  ND4D1BWP30P140LVT U136 ( .A1(n106), .A2(n105), .A3(n104), .A4(n103), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U137 ( .A1(n147), .A2(i_data_bus[158]), .B1(n177), .B2(
        i_data_bus[30]), .ZN(n110) );
  AOI22D1BWP30P140LVT U138 ( .A1(n178), .A2(i_data_bus[62]), .B1(n164), .B2(
        i_data_bus[126]), .ZN(n109) );
  AOI22D1BWP30P140LVT U139 ( .A1(n170), .A2(i_data_bus[222]), .B1(n1), .B2(
        i_data_bus[190]), .ZN(n108) );
  AOI22D1BWP30P140LVT U140 ( .A1(n181), .A2(i_data_bus[254]), .B1(n180), .B2(
        i_data_bus[94]), .ZN(n107) );
  ND4D1BWP30P140LVT U141 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U142 ( .A1(n147), .A2(i_data_bus[157]), .B1(n177), .B2(
        i_data_bus[29]), .ZN(n114) );
  AOI22D1BWP30P140LVT U143 ( .A1(n178), .A2(i_data_bus[61]), .B1(n164), .B2(
        i_data_bus[125]), .ZN(n113) );
  AOI22D1BWP30P140LVT U144 ( .A1(n170), .A2(i_data_bus[221]), .B1(n1), .B2(
        i_data_bus[189]), .ZN(n112) );
  AOI22D1BWP30P140LVT U145 ( .A1(n181), .A2(i_data_bus[253]), .B1(n180), .B2(
        i_data_bus[93]), .ZN(n111) );
  ND4D1BWP30P140LVT U146 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U147 ( .A1(n147), .A2(i_data_bus[156]), .B1(n177), .B2(
        i_data_bus[28]), .ZN(n118) );
  AOI22D1BWP30P140LVT U148 ( .A1(n178), .A2(i_data_bus[60]), .B1(n164), .B2(
        i_data_bus[124]), .ZN(n117) );
  AOI22D1BWP30P140LVT U149 ( .A1(n170), .A2(i_data_bus[220]), .B1(n1), .B2(
        i_data_bus[188]), .ZN(n116) );
  AOI22D1BWP30P140LVT U150 ( .A1(n181), .A2(i_data_bus[252]), .B1(n180), .B2(
        i_data_bus[92]), .ZN(n115) );
  ND4D1BWP30P140LVT U151 ( .A1(n118), .A2(n117), .A3(n116), .A4(n115), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U152 ( .A1(n147), .A2(i_data_bus[155]), .B1(n177), .B2(
        i_data_bus[27]), .ZN(n122) );
  AOI22D1BWP30P140LVT U153 ( .A1(n178), .A2(i_data_bus[59]), .B1(n164), .B2(
        i_data_bus[123]), .ZN(n121) );
  AOI22D1BWP30P140LVT U154 ( .A1(n170), .A2(i_data_bus[219]), .B1(n1), .B2(
        i_data_bus[187]), .ZN(n120) );
  AOI22D1BWP30P140LVT U155 ( .A1(n181), .A2(i_data_bus[251]), .B1(n180), .B2(
        i_data_bus[91]), .ZN(n119) );
  ND4D1BWP30P140LVT U156 ( .A1(n122), .A2(n121), .A3(n120), .A4(n119), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U157 ( .A1(n147), .A2(i_data_bus[154]), .B1(n177), .B2(
        i_data_bus[26]), .ZN(n126) );
  AOI22D1BWP30P140LVT U158 ( .A1(n178), .A2(i_data_bus[58]), .B1(n164), .B2(
        i_data_bus[122]), .ZN(n125) );
  AOI22D1BWP30P140LVT U159 ( .A1(n170), .A2(i_data_bus[218]), .B1(n1), .B2(
        i_data_bus[186]), .ZN(n124) );
  AOI22D1BWP30P140LVT U160 ( .A1(n181), .A2(i_data_bus[250]), .B1(n180), .B2(
        i_data_bus[90]), .ZN(n123) );
  ND4D1BWP30P140LVT U161 ( .A1(n126), .A2(n125), .A3(n124), .A4(n123), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U162 ( .A1(n147), .A2(i_data_bus[153]), .B1(n177), .B2(
        i_data_bus[25]), .ZN(n130) );
  AOI22D1BWP30P140LVT U163 ( .A1(n178), .A2(i_data_bus[57]), .B1(n164), .B2(
        i_data_bus[121]), .ZN(n129) );
  AOI22D1BWP30P140LVT U164 ( .A1(n170), .A2(i_data_bus[217]), .B1(n1), .B2(
        i_data_bus[185]), .ZN(n128) );
  AOI22D1BWP30P140LVT U165 ( .A1(n181), .A2(i_data_bus[249]), .B1(n180), .B2(
        i_data_bus[89]), .ZN(n127) );
  ND4D1BWP30P140LVT U166 ( .A1(n130), .A2(n129), .A3(n128), .A4(n127), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U167 ( .A1(n147), .A2(i_data_bus[152]), .B1(n177), .B2(
        i_data_bus[24]), .ZN(n134) );
  AOI22D1BWP30P140LVT U168 ( .A1(n178), .A2(i_data_bus[56]), .B1(n164), .B2(
        i_data_bus[120]), .ZN(n133) );
  AOI22D1BWP30P140LVT U169 ( .A1(n170), .A2(i_data_bus[216]), .B1(n1), .B2(
        i_data_bus[184]), .ZN(n132) );
  AOI22D1BWP30P140LVT U170 ( .A1(n181), .A2(i_data_bus[248]), .B1(n180), .B2(
        i_data_bus[88]), .ZN(n131) );
  ND4D1BWP30P140LVT U171 ( .A1(n134), .A2(n133), .A3(n132), .A4(n131), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U172 ( .A1(n147), .A2(i_data_bus[151]), .B1(n177), .B2(
        i_data_bus[23]), .ZN(n138) );
  AOI22D1BWP30P140LVT U173 ( .A1(n178), .A2(i_data_bus[55]), .B1(n164), .B2(
        i_data_bus[119]), .ZN(n137) );
  AOI22D1BWP30P140LVT U174 ( .A1(n170), .A2(i_data_bus[215]), .B1(n1), .B2(
        i_data_bus[183]), .ZN(n136) );
  AOI22D1BWP30P140LVT U175 ( .A1(n181), .A2(i_data_bus[247]), .B1(n180), .B2(
        i_data_bus[87]), .ZN(n135) );
  ND4D1BWP30P140LVT U176 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U177 ( .A1(n147), .A2(i_data_bus[150]), .B1(n177), .B2(
        i_data_bus[22]), .ZN(n142) );
  AOI22D1BWP30P140LVT U178 ( .A1(n178), .A2(i_data_bus[54]), .B1(n164), .B2(
        i_data_bus[118]), .ZN(n141) );
  AOI22D1BWP30P140LVT U179 ( .A1(n170), .A2(i_data_bus[214]), .B1(n1), .B2(
        i_data_bus[182]), .ZN(n140) );
  AOI22D1BWP30P140LVT U180 ( .A1(n181), .A2(i_data_bus[246]), .B1(n180), .B2(
        i_data_bus[86]), .ZN(n139) );
  ND4D1BWP30P140LVT U181 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U182 ( .A1(n147), .A2(i_data_bus[149]), .B1(n177), .B2(
        i_data_bus[21]), .ZN(n146) );
  AOI22D1BWP30P140LVT U183 ( .A1(n178), .A2(i_data_bus[53]), .B1(n164), .B2(
        i_data_bus[117]), .ZN(n145) );
  AOI22D1BWP30P140LVT U184 ( .A1(n170), .A2(i_data_bus[213]), .B1(n1), .B2(
        i_data_bus[181]), .ZN(n144) );
  AOI22D1BWP30P140LVT U185 ( .A1(n181), .A2(i_data_bus[245]), .B1(n180), .B2(
        i_data_bus[85]), .ZN(n143) );
  ND4D1BWP30P140LVT U186 ( .A1(n146), .A2(n145), .A3(n144), .A4(n143), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U187 ( .A1(n147), .A2(i_data_bus[148]), .B1(n177), .B2(
        i_data_bus[20]), .ZN(n151) );
  AOI22D1BWP30P140LVT U188 ( .A1(n178), .A2(i_data_bus[52]), .B1(n164), .B2(
        i_data_bus[116]), .ZN(n150) );
  AOI22D1BWP30P140LVT U189 ( .A1(n170), .A2(i_data_bus[212]), .B1(n1), .B2(
        i_data_bus[180]), .ZN(n149) );
  AOI22D1BWP30P140LVT U190 ( .A1(n181), .A2(i_data_bus[244]), .B1(n180), .B2(
        i_data_bus[84]), .ZN(n148) );
  ND4D1BWP30P140LVT U191 ( .A1(n151), .A2(n150), .A3(n149), .A4(n148), .ZN(
        N389) );
  INVD1BWP30P140LVT U192 ( .I(i_data_bus[147]), .ZN(n152) );
  MAOI22D1BWP30P140LVT U193 ( .A1(n177), .A2(i_data_bus[19]), .B1(n176), .B2(
        n152), .ZN(n156) );
  AOI22D1BWP30P140LVT U194 ( .A1(n178), .A2(i_data_bus[51]), .B1(n164), .B2(
        i_data_bus[115]), .ZN(n155) );
  AOI22D1BWP30P140LVT U195 ( .A1(n170), .A2(i_data_bus[211]), .B1(n1), .B2(
        i_data_bus[179]), .ZN(n154) );
  AOI22D1BWP30P140LVT U196 ( .A1(n181), .A2(i_data_bus[243]), .B1(n180), .B2(
        i_data_bus[83]), .ZN(n153) );
  ND4D1BWP30P140LVT U197 ( .A1(n156), .A2(n155), .A3(n154), .A4(n153), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U198 ( .A1(n157), .A2(i_data_bus[141]), .B1(n177), .B2(
        i_data_bus[13]), .ZN(n162) );
  AOI22D1BWP30P140LVT U199 ( .A1(n178), .A2(i_data_bus[45]), .B1(n164), .B2(
        i_data_bus[109]), .ZN(n161) );
  AOI22D1BWP30P140LVT U200 ( .A1(n179), .A2(i_data_bus[205]), .B1(n1), .B2(
        i_data_bus[173]), .ZN(n160) );
  AOI22D1BWP30P140LVT U201 ( .A1(n181), .A2(i_data_bus[237]), .B1(n158), .B2(
        i_data_bus[77]), .ZN(n159) );
  ND4D1BWP30P140LVT U202 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .ZN(
        N382) );
  INVD1BWP30P140LVT U203 ( .I(i_data_bus[146]), .ZN(n163) );
  MAOI22D1BWP30P140LVT U204 ( .A1(n177), .A2(i_data_bus[18]), .B1(n176), .B2(
        n163), .ZN(n168) );
  AOI22D1BWP30P140LVT U205 ( .A1(n178), .A2(i_data_bus[50]), .B1(n164), .B2(
        i_data_bus[114]), .ZN(n167) );
  AOI22D1BWP30P140LVT U206 ( .A1(n170), .A2(i_data_bus[210]), .B1(n1), .B2(
        i_data_bus[178]), .ZN(n166) );
  AOI22D1BWP30P140LVT U207 ( .A1(n181), .A2(i_data_bus[242]), .B1(n180), .B2(
        i_data_bus[82]), .ZN(n165) );
  ND4D1BWP30P140LVT U208 ( .A1(n168), .A2(n167), .A3(n166), .A4(n165), .ZN(
        N387) );
  INVD1BWP30P140LVT U209 ( .I(i_data_bus[145]), .ZN(n169) );
  MAOI22D1BWP30P140LVT U210 ( .A1(n177), .A2(i_data_bus[17]), .B1(n176), .B2(
        n169), .ZN(n174) );
  AOI22D1BWP30P140LVT U211 ( .A1(n178), .A2(i_data_bus[49]), .B1(n164), .B2(
        i_data_bus[113]), .ZN(n173) );
  AOI22D1BWP30P140LVT U212 ( .A1(n170), .A2(i_data_bus[209]), .B1(n1), .B2(
        i_data_bus[177]), .ZN(n172) );
  AOI22D1BWP30P140LVT U213 ( .A1(n181), .A2(i_data_bus[241]), .B1(n180), .B2(
        i_data_bus[81]), .ZN(n171) );
  ND4D1BWP30P140LVT U214 ( .A1(n174), .A2(n173), .A3(n172), .A4(n171), .ZN(
        N386) );
  INVD1BWP30P140LVT U215 ( .I(i_data_bus[144]), .ZN(n175) );
  MAOI22D1BWP30P140LVT U216 ( .A1(n177), .A2(i_data_bus[16]), .B1(n176), .B2(
        n175), .ZN(n185) );
  AOI22D1BWP30P140LVT U217 ( .A1(i_data_bus[112]), .A2(n164), .B1(n178), .B2(
        i_data_bus[48]), .ZN(n184) );
  AOI22D1BWP30P140LVT U218 ( .A1(n179), .A2(i_data_bus[208]), .B1(n1), .B2(
        i_data_bus[176]), .ZN(n183) );
  AOI22D1BWP30P140LVT U219 ( .A1(n181), .A2(i_data_bus[240]), .B1(n180), .B2(
        i_data_bus[80]), .ZN(n182) );
  ND4D1BWP30P140LVT U220 ( .A1(n185), .A2(n184), .A3(n183), .A4(n182), .ZN(
        N385) );
endmodule


module mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_7 ( CLK, 
        rst, i_valid, i_data_bus, o_valid, o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [0:0] o_valid;
  output [31:0] o_data_bus;
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  wire   N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N402, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;

  DFQD1BWP30P140LVT o_valid_reg_reg_0_ ( .D(N402), .CP(CLK), .Q(o_valid[0]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N400), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N399), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N398), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N397), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N396), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N395), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N394), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(N393), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(N392), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(N391), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(N390), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(N389), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(N388), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(N387), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(N386), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(N385), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(N384), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(N383), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(N382), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(N381), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(N380), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(N379), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(N378), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(N377), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(N376), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(N375), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(N374), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(N373), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(N372), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(N371), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(N370), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD1BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(N369), .CP(CLK), .Q(
        o_data_bus[0]) );
  INVD4BWP30P140LVT U3 ( .I(n54), .ZN(n184) );
  INVD3BWP30P140LVT U4 ( .I(n15), .ZN(n186) );
  INVD4BWP30P140LVT U5 ( .I(n54), .ZN(n104) );
  INVD1BWP30P140LVT U6 ( .I(n23), .ZN(n43) );
  BUFFD4BWP30P140LVT U7 ( .I(n33), .Z(n183) );
  INR2D1BWP30P140LVT U8 ( .A1(n13), .B1(n12), .ZN(n14) );
  INR2D1BWP30P140LVT U9 ( .A1(n36), .B1(n32), .ZN(n33) );
  INVD0P7BWP30P140LVT U10 ( .I(i_cmd[4]), .ZN(n26) );
  NR2D2BWP30P140LVT U11 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n31) );
  CKND2D3BWP30P140LVT U12 ( .A1(n18), .A2(n17), .ZN(n24) );
  NR2OPTPAD2BWP30P140LVT U13 ( .A1(i_cmd[5]), .A2(i_cmd[6]), .ZN(n18) );
  INR2D2BWP30P140LVT U14 ( .A1(n16), .B1(i_cmd[7]), .ZN(n17) );
  INVD1BWP30P140LVT U15 ( .I(n13), .ZN(n8) );
  INVD1BWP30P140LVT U16 ( .I(n14), .ZN(n15) );
  ND2D1BWP30P140LVT U17 ( .A1(n47), .A2(n46), .ZN(n48) );
  INR2D2BWP30P140LVT U18 ( .A1(n19), .B1(n24), .ZN(n36) );
  NR2D3BWP30P140LVT U19 ( .A1(i_cmd[0]), .A2(i_cmd[4]), .ZN(n19) );
  NR4D1BWP30P140LVT U20 ( .A1(n8), .A2(i_cmd[5]), .A3(n4), .A4(n3), .ZN(n5) );
  INVD1BWP30P140LVT U21 ( .I(i_cmd[6]), .ZN(n3) );
  NR4D1BWP30P140LVT U22 ( .A1(n8), .A2(i_cmd[6]), .A3(n7), .A4(n6), .ZN(n9) );
  INVD1BWP30P140LVT U23 ( .I(i_cmd[5]), .ZN(n7) );
  INVD1BWP30P140LVT U24 ( .I(n36), .ZN(n22) );
  INVD1BWP30P140LVT U25 ( .I(i_cmd[0]), .ZN(n29) );
  INR2D4BWP30P140LVT U26 ( .A1(n36), .B1(n35), .ZN(n182) );
  ND2D1BWP30P140LVT U27 ( .A1(n53), .A2(n52), .ZN(N402) );
  INVD1BWP30P140LVT U28 ( .I(n5), .ZN(n103) );
  NR2D3BWP30P140LVT U29 ( .A1(i_cmd[1]), .A2(i_cmd[2]), .ZN(n34) );
  INR2D1BWP30P140LVT U30 ( .A1(i_en), .B1(rst), .ZN(n16) );
  INR2D1BWP30P140LVT U31 ( .A1(n16), .B1(i_cmd[3]), .ZN(n1) );
  ND2OPTIBD1BWP30P140LVT U32 ( .A1(n34), .A2(n1), .ZN(n2) );
  INR2D2BWP30P140LVT U33 ( .A1(n19), .B1(n2), .ZN(n13) );
  IND2D1BWP30P140LVT U34 ( .A1(i_cmd[7]), .B1(i_valid[6]), .ZN(n4) );
  INVD2BWP30P140LVT U35 ( .I(n103), .ZN(n122) );
  IND2D1BWP30P140LVT U36 ( .A1(i_cmd[7]), .B1(i_valid[5]), .ZN(n6) );
  INVD2BWP30P140LVT U37 ( .I(n9), .ZN(n54) );
  AOI22D1BWP30P140LVT U38 ( .A1(n122), .A2(i_data_bus[206]), .B1(n184), .B2(
        i_data_bus[174]), .ZN(n42) );
  INVD1BWP30P140LVT U39 ( .I(i_cmd[7]), .ZN(n10) );
  INR2D1BWP30P140LVT U40 ( .A1(i_valid[7]), .B1(n10), .ZN(n11) );
  ND2OPTIBD1BWP30P140LVT U41 ( .A1(n18), .A2(n11), .ZN(n12) );
  INVD1BWP30P140LVT U42 ( .I(i_cmd[2]), .ZN(n21) );
  IND2D1BWP30P140LVT U43 ( .A1(i_cmd[3]), .B1(i_valid[2]), .ZN(n20) );
  NR4D0BWP30P140LVT U44 ( .A1(n22), .A2(i_cmd[1]), .A3(n21), .A4(n20), .ZN(n23) );
  INVD2BWP30P140LVT U45 ( .I(n43), .ZN(n123) );
  AOI22D1BWP30P140LVT U46 ( .A1(n186), .A2(i_data_bus[238]), .B1(n123), .B2(
        i_data_bus[78]), .ZN(n41) );
  INVD2BWP30P140LVT U47 ( .I(n24), .ZN(n25) );
  IND3D4BWP30P140LVT U48 ( .A1(i_cmd[1]), .B1(n31), .B2(n25), .ZN(n28) );
  INR4D1BWP30P140LVT U49 ( .A1(i_valid[4]), .B1(i_cmd[0]), .B2(n26), .B3(n28), 
        .ZN(n27) );
  INVD2BWP30P140LVT U50 ( .I(n27), .ZN(n116) );
  INVD2BWP30P140LVT U51 ( .I(n116), .ZN(n121) );
  INR4D1BWP30P140LVT U52 ( .A1(i_valid[0]), .B1(i_cmd[4]), .B2(n29), .B3(n28), 
        .ZN(n30) );
  INVD2BWP30P140LVT U53 ( .I(n30), .ZN(n110) );
  INVD8BWP30P140LVT U54 ( .I(n110), .ZN(n180) );
  AOI22D4BWP30P140LVT U55 ( .A1(n121), .A2(i_data_bus[142]), .B1(n180), .B2(
        i_data_bus[14]), .ZN(n38) );
  ND3D1BWP30P140LVT U56 ( .A1(n31), .A2(i_valid[1]), .A3(i_cmd[1]), .ZN(n32)
         );
  ND3D2BWP30P140LVT U57 ( .A1(n34), .A2(i_valid[3]), .A3(i_cmd[3]), .ZN(n35)
         );
  AOI22D1BWP30P140LVT U58 ( .A1(n183), .A2(i_data_bus[46]), .B1(n182), .B2(
        i_data_bus[110]), .ZN(n37) );
  ND2D2BWP30P140LVT U59 ( .A1(n38), .A2(n37), .ZN(n39) );
  INVD1BWP30P140LVT U60 ( .I(n39), .ZN(n40) );
  ND3D1BWP30P140LVT U61 ( .A1(n42), .A2(n41), .A3(n40), .ZN(N383) );
  INVD2BWP30P140LVT U62 ( .I(n43), .ZN(n44) );
  AOI22D1BWP30P140LVT U63 ( .A1(n186), .A2(i_data_bus[240]), .B1(n44), .B2(
        i_data_bus[80]), .ZN(n51) );
  AOI22D1BWP30P140LVT U64 ( .A1(n122), .A2(i_data_bus[208]), .B1(n184), .B2(
        i_data_bus[176]), .ZN(n50) );
  INVD2BWP30P140LVT U65 ( .I(n116), .ZN(n181) );
  INVD1BWP30P140LVT U66 ( .I(i_data_bus[16]), .ZN(n45) );
  MAOI22D1BWP30P140LVT U67 ( .A1(n181), .A2(i_data_bus[144]), .B1(n110), .B2(
        n45), .ZN(n47) );
  AOI22D1BWP30P140LVT U68 ( .A1(n183), .A2(i_data_bus[48]), .B1(n182), .B2(
        i_data_bus[112]), .ZN(n46) );
  INVD1BWP30P140LVT U69 ( .I(n48), .ZN(n49) );
  ND3D1BWP30P140LVT U70 ( .A1(n51), .A2(n50), .A3(n49), .ZN(N385) );
  NR4D0BWP30P140LVT U71 ( .A1(n183), .A2(n182), .A3(n181), .A4(n180), .ZN(n53)
         );
  INVD2BWP30P140LVT U72 ( .I(n103), .ZN(n185) );
  NR4D0BWP30P140LVT U73 ( .A1(n186), .A2(n185), .A3(n44), .A4(n184), .ZN(n52)
         );
  AOI22D1BWP30P140LVT U74 ( .A1(n121), .A2(i_data_bus[140]), .B1(n180), .B2(
        i_data_bus[12]), .ZN(n58) );
  AOI22D1BWP30P140LVT U75 ( .A1(n183), .A2(i_data_bus[44]), .B1(n182), .B2(
        i_data_bus[108]), .ZN(n57) );
  AOI22D1BWP30P140LVT U76 ( .A1(n122), .A2(i_data_bus[204]), .B1(n104), .B2(
        i_data_bus[172]), .ZN(n56) );
  AOI22D1BWP30P140LVT U77 ( .A1(n186), .A2(i_data_bus[236]), .B1(n123), .B2(
        i_data_bus[76]), .ZN(n55) );
  ND4D1BWP30P140LVT U78 ( .A1(n58), .A2(n57), .A3(n56), .A4(n55), .ZN(N381) );
  AOI22D1BWP30P140LVT U79 ( .A1(n121), .A2(i_data_bus[139]), .B1(n180), .B2(
        i_data_bus[11]), .ZN(n62) );
  AOI22D1BWP30P140LVT U80 ( .A1(n183), .A2(i_data_bus[43]), .B1(n182), .B2(
        i_data_bus[107]), .ZN(n61) );
  AOI22D1BWP30P140LVT U81 ( .A1(n122), .A2(i_data_bus[203]), .B1(n104), .B2(
        i_data_bus[171]), .ZN(n60) );
  AOI22D1BWP30P140LVT U82 ( .A1(n186), .A2(i_data_bus[235]), .B1(n123), .B2(
        i_data_bus[75]), .ZN(n59) );
  ND4D1BWP30P140LVT U83 ( .A1(n62), .A2(n61), .A3(n60), .A4(n59), .ZN(N380) );
  AOI22D1BWP30P140LVT U84 ( .A1(n121), .A2(i_data_bus[138]), .B1(n180), .B2(
        i_data_bus[10]), .ZN(n66) );
  AOI22D1BWP30P140LVT U85 ( .A1(n183), .A2(i_data_bus[42]), .B1(n182), .B2(
        i_data_bus[106]), .ZN(n65) );
  AOI22D1BWP30P140LVT U86 ( .A1(n122), .A2(i_data_bus[202]), .B1(n104), .B2(
        i_data_bus[170]), .ZN(n64) );
  AOI22D1BWP30P140LVT U87 ( .A1(n186), .A2(i_data_bus[234]), .B1(n123), .B2(
        i_data_bus[74]), .ZN(n63) );
  ND4D1BWP30P140LVT U88 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(N379) );
  AOI22D1BWP30P140LVT U89 ( .A1(n121), .A2(i_data_bus[137]), .B1(n180), .B2(
        i_data_bus[9]), .ZN(n70) );
  AOI22D1BWP30P140LVT U90 ( .A1(n183), .A2(i_data_bus[41]), .B1(n182), .B2(
        i_data_bus[105]), .ZN(n69) );
  AOI22D1BWP30P140LVT U91 ( .A1(n122), .A2(i_data_bus[201]), .B1(n104), .B2(
        i_data_bus[169]), .ZN(n68) );
  AOI22D1BWP30P140LVT U92 ( .A1(n186), .A2(i_data_bus[233]), .B1(n123), .B2(
        i_data_bus[73]), .ZN(n67) );
  ND4D1BWP30P140LVT U93 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(N378) );
  AOI22D1BWP30P140LVT U94 ( .A1(n121), .A2(i_data_bus[136]), .B1(n180), .B2(
        i_data_bus[8]), .ZN(n74) );
  AOI22D1BWP30P140LVT U95 ( .A1(n183), .A2(i_data_bus[40]), .B1(n182), .B2(
        i_data_bus[104]), .ZN(n73) );
  AOI22D1BWP30P140LVT U96 ( .A1(n122), .A2(i_data_bus[200]), .B1(n104), .B2(
        i_data_bus[168]), .ZN(n72) );
  AOI22D1BWP30P140LVT U97 ( .A1(n186), .A2(i_data_bus[232]), .B1(n123), .B2(
        i_data_bus[72]), .ZN(n71) );
  ND4D1BWP30P140LVT U98 ( .A1(n74), .A2(n73), .A3(n72), .A4(n71), .ZN(N377) );
  AOI22D1BWP30P140LVT U99 ( .A1(n121), .A2(i_data_bus[135]), .B1(n180), .B2(
        i_data_bus[7]), .ZN(n78) );
  AOI22D1BWP30P140LVT U100 ( .A1(n183), .A2(i_data_bus[39]), .B1(n182), .B2(
        i_data_bus[103]), .ZN(n77) );
  AOI22D1BWP30P140LVT U101 ( .A1(n122), .A2(i_data_bus[199]), .B1(n104), .B2(
        i_data_bus[167]), .ZN(n76) );
  AOI22D1BWP30P140LVT U102 ( .A1(n186), .A2(i_data_bus[231]), .B1(n123), .B2(
        i_data_bus[71]), .ZN(n75) );
  ND4D1BWP30P140LVT U103 ( .A1(n78), .A2(n77), .A3(n76), .A4(n75), .ZN(N376)
         );
  AOI22D1BWP30P140LVT U104 ( .A1(n121), .A2(i_data_bus[134]), .B1(n180), .B2(
        i_data_bus[6]), .ZN(n82) );
  AOI22D1BWP30P140LVT U105 ( .A1(n183), .A2(i_data_bus[38]), .B1(n182), .B2(
        i_data_bus[102]), .ZN(n81) );
  AOI22D1BWP30P140LVT U106 ( .A1(n122), .A2(i_data_bus[198]), .B1(n104), .B2(
        i_data_bus[166]), .ZN(n80) );
  AOI22D1BWP30P140LVT U107 ( .A1(n186), .A2(i_data_bus[230]), .B1(n123), .B2(
        i_data_bus[70]), .ZN(n79) );
  ND4D1BWP30P140LVT U108 ( .A1(n82), .A2(n81), .A3(n80), .A4(n79), .ZN(N375)
         );
  AOI22D1BWP30P140LVT U109 ( .A1(n121), .A2(i_data_bus[133]), .B1(n180), .B2(
        i_data_bus[5]), .ZN(n86) );
  AOI22D1BWP30P140LVT U110 ( .A1(n183), .A2(i_data_bus[37]), .B1(n182), .B2(
        i_data_bus[101]), .ZN(n85) );
  AOI22D1BWP30P140LVT U111 ( .A1(n122), .A2(i_data_bus[197]), .B1(n104), .B2(
        i_data_bus[165]), .ZN(n84) );
  AOI22D1BWP30P140LVT U112 ( .A1(n186), .A2(i_data_bus[229]), .B1(n123), .B2(
        i_data_bus[69]), .ZN(n83) );
  ND4D1BWP30P140LVT U113 ( .A1(n86), .A2(n85), .A3(n84), .A4(n83), .ZN(N374)
         );
  AOI22D1BWP30P140LVT U114 ( .A1(n121), .A2(i_data_bus[132]), .B1(n180), .B2(
        i_data_bus[4]), .ZN(n90) );
  AOI22D1BWP30P140LVT U115 ( .A1(n183), .A2(i_data_bus[36]), .B1(n182), .B2(
        i_data_bus[100]), .ZN(n89) );
  AOI22D1BWP30P140LVT U116 ( .A1(n122), .A2(i_data_bus[196]), .B1(n104), .B2(
        i_data_bus[164]), .ZN(n88) );
  AOI22D1BWP30P140LVT U117 ( .A1(n186), .A2(i_data_bus[228]), .B1(n123), .B2(
        i_data_bus[68]), .ZN(n87) );
  ND4D1BWP30P140LVT U118 ( .A1(n90), .A2(n89), .A3(n88), .A4(n87), .ZN(N373)
         );
  AOI22D1BWP30P140LVT U119 ( .A1(n121), .A2(i_data_bus[131]), .B1(n180), .B2(
        i_data_bus[3]), .ZN(n94) );
  AOI22D1BWP30P140LVT U120 ( .A1(n183), .A2(i_data_bus[35]), .B1(n182), .B2(
        i_data_bus[99]), .ZN(n93) );
  AOI22D1BWP30P140LVT U121 ( .A1(n122), .A2(i_data_bus[195]), .B1(n104), .B2(
        i_data_bus[163]), .ZN(n92) );
  AOI22D1BWP30P140LVT U122 ( .A1(n186), .A2(i_data_bus[227]), .B1(n123), .B2(
        i_data_bus[67]), .ZN(n91) );
  ND4D1BWP30P140LVT U123 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .ZN(N372)
         );
  AOI22D1BWP30P140LVT U124 ( .A1(n121), .A2(i_data_bus[130]), .B1(n180), .B2(
        i_data_bus[2]), .ZN(n98) );
  AOI22D1BWP30P140LVT U125 ( .A1(n183), .A2(i_data_bus[34]), .B1(n182), .B2(
        i_data_bus[98]), .ZN(n97) );
  AOI22D1BWP30P140LVT U126 ( .A1(n122), .A2(i_data_bus[194]), .B1(n104), .B2(
        i_data_bus[162]), .ZN(n96) );
  AOI22D1BWP30P140LVT U127 ( .A1(n186), .A2(i_data_bus[226]), .B1(n123), .B2(
        i_data_bus[66]), .ZN(n95) );
  ND4D1BWP30P140LVT U128 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .ZN(N371)
         );
  AOI22D1BWP30P140LVT U129 ( .A1(n121), .A2(i_data_bus[129]), .B1(n180), .B2(
        i_data_bus[1]), .ZN(n102) );
  AOI22D1BWP30P140LVT U130 ( .A1(n183), .A2(i_data_bus[33]), .B1(n182), .B2(
        i_data_bus[97]), .ZN(n101) );
  AOI22D1BWP30P140LVT U131 ( .A1(n122), .A2(i_data_bus[193]), .B1(n104), .B2(
        i_data_bus[161]), .ZN(n100) );
  AOI22D1BWP30P140LVT U132 ( .A1(n186), .A2(i_data_bus[225]), .B1(n123), .B2(
        i_data_bus[65]), .ZN(n99) );
  ND4D1BWP30P140LVT U133 ( .A1(n102), .A2(n101), .A3(n100), .A4(n99), .ZN(N370) );
  AOI22D1BWP30P140LVT U134 ( .A1(n121), .A2(i_data_bus[128]), .B1(n180), .B2(
        i_data_bus[0]), .ZN(n108) );
  AOI22D1BWP30P140LVT U135 ( .A1(n183), .A2(i_data_bus[32]), .B1(n182), .B2(
        i_data_bus[96]), .ZN(n107) );
  AOI22D1BWP30P140LVT U136 ( .A1(n185), .A2(i_data_bus[192]), .B1(n104), .B2(
        i_data_bus[160]), .ZN(n106) );
  AOI22D1BWP30P140LVT U137 ( .A1(n186), .A2(i_data_bus[224]), .B1(n123), .B2(
        i_data_bus[64]), .ZN(n105) );
  ND4D1BWP30P140LVT U138 ( .A1(n108), .A2(n107), .A3(n106), .A4(n105), .ZN(
        N369) );
  INVD1BWP30P140LVT U139 ( .I(i_data_bus[15]), .ZN(n109) );
  MAOI22D1BWP30P140LVT U140 ( .A1(n121), .A2(i_data_bus[143]), .B1(n110), .B2(
        n109), .ZN(n114) );
  AOI22D1BWP30P140LVT U141 ( .A1(n183), .A2(i_data_bus[47]), .B1(n182), .B2(
        i_data_bus[111]), .ZN(n113) );
  AOI22D1BWP30P140LVT U142 ( .A1(n122), .A2(i_data_bus[207]), .B1(n184), .B2(
        i_data_bus[175]), .ZN(n112) );
  AOI22D1BWP30P140LVT U143 ( .A1(n186), .A2(i_data_bus[239]), .B1(n123), .B2(
        i_data_bus[79]), .ZN(n111) );
  ND4D1BWP30P140LVT U144 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(
        N384) );
  INVD1BWP30P140LVT U145 ( .I(i_data_bus[152]), .ZN(n115) );
  MAOI22D1BWP30P140LVT U146 ( .A1(n180), .A2(i_data_bus[24]), .B1(n116), .B2(
        n115), .ZN(n120) );
  AOI22D1BWP30P140LVT U147 ( .A1(n183), .A2(i_data_bus[56]), .B1(n182), .B2(
        i_data_bus[120]), .ZN(n119) );
  AOI22D1BWP30P140LVT U148 ( .A1(n185), .A2(i_data_bus[216]), .B1(n184), .B2(
        i_data_bus[184]), .ZN(n118) );
  AOI22D1BWP30P140LVT U149 ( .A1(n186), .A2(i_data_bus[248]), .B1(n44), .B2(
        i_data_bus[88]), .ZN(n117) );
  ND4D1BWP30P140LVT U150 ( .A1(n120), .A2(n119), .A3(n118), .A4(n117), .ZN(
        N393) );
  AOI22D1BWP30P140LVT U151 ( .A1(n121), .A2(i_data_bus[141]), .B1(n180), .B2(
        i_data_bus[13]), .ZN(n127) );
  AOI22D1BWP30P140LVT U152 ( .A1(n183), .A2(i_data_bus[45]), .B1(n182), .B2(
        i_data_bus[109]), .ZN(n126) );
  AOI22D1BWP30P140LVT U153 ( .A1(n122), .A2(i_data_bus[205]), .B1(n184), .B2(
        i_data_bus[173]), .ZN(n125) );
  AOI22D1BWP30P140LVT U154 ( .A1(n186), .A2(i_data_bus[237]), .B1(n123), .B2(
        i_data_bus[77]), .ZN(n124) );
  ND4D1BWP30P140LVT U155 ( .A1(n127), .A2(n126), .A3(n125), .A4(n124), .ZN(
        N382) );
  AOI22D1BWP30P140LVT U156 ( .A1(n181), .A2(i_data_bus[159]), .B1(n180), .B2(
        i_data_bus[31]), .ZN(n131) );
  AOI22D1BWP30P140LVT U157 ( .A1(n183), .A2(i_data_bus[63]), .B1(n182), .B2(
        i_data_bus[127]), .ZN(n130) );
  AOI22D1BWP30P140LVT U158 ( .A1(n185), .A2(i_data_bus[223]), .B1(n184), .B2(
        i_data_bus[191]), .ZN(n129) );
  AOI22D1BWP30P140LVT U159 ( .A1(n186), .A2(i_data_bus[255]), .B1(n44), .B2(
        i_data_bus[95]), .ZN(n128) );
  ND4D1BWP30P140LVT U160 ( .A1(n131), .A2(n130), .A3(n129), .A4(n128), .ZN(
        N400) );
  AOI22D1BWP30P140LVT U161 ( .A1(n181), .A2(i_data_bus[158]), .B1(n180), .B2(
        i_data_bus[30]), .ZN(n135) );
  AOI22D1BWP30P140LVT U162 ( .A1(n183), .A2(i_data_bus[62]), .B1(n182), .B2(
        i_data_bus[126]), .ZN(n134) );
  AOI22D1BWP30P140LVT U163 ( .A1(n185), .A2(i_data_bus[222]), .B1(n184), .B2(
        i_data_bus[190]), .ZN(n133) );
  AOI22D1BWP30P140LVT U164 ( .A1(n186), .A2(i_data_bus[254]), .B1(n44), .B2(
        i_data_bus[94]), .ZN(n132) );
  ND4D1BWP30P140LVT U165 ( .A1(n135), .A2(n134), .A3(n133), .A4(n132), .ZN(
        N399) );
  AOI22D1BWP30P140LVT U166 ( .A1(n181), .A2(i_data_bus[157]), .B1(n180), .B2(
        i_data_bus[29]), .ZN(n139) );
  AOI22D1BWP30P140LVT U167 ( .A1(n183), .A2(i_data_bus[61]), .B1(n182), .B2(
        i_data_bus[125]), .ZN(n138) );
  AOI22D1BWP30P140LVT U168 ( .A1(n185), .A2(i_data_bus[221]), .B1(n184), .B2(
        i_data_bus[189]), .ZN(n137) );
  AOI22D1BWP30P140LVT U169 ( .A1(n186), .A2(i_data_bus[253]), .B1(n44), .B2(
        i_data_bus[93]), .ZN(n136) );
  ND4D1BWP30P140LVT U170 ( .A1(n139), .A2(n138), .A3(n137), .A4(n136), .ZN(
        N398) );
  AOI22D1BWP30P140LVT U171 ( .A1(n181), .A2(i_data_bus[156]), .B1(n180), .B2(
        i_data_bus[28]), .ZN(n143) );
  AOI22D1BWP30P140LVT U172 ( .A1(n183), .A2(i_data_bus[60]), .B1(n182), .B2(
        i_data_bus[124]), .ZN(n142) );
  AOI22D1BWP30P140LVT U173 ( .A1(n185), .A2(i_data_bus[220]), .B1(n184), .B2(
        i_data_bus[188]), .ZN(n141) );
  AOI22D1BWP30P140LVT U174 ( .A1(n186), .A2(i_data_bus[252]), .B1(n44), .B2(
        i_data_bus[92]), .ZN(n140) );
  ND4D1BWP30P140LVT U175 ( .A1(n143), .A2(n142), .A3(n141), .A4(n140), .ZN(
        N397) );
  AOI22D1BWP30P140LVT U176 ( .A1(n181), .A2(i_data_bus[155]), .B1(n180), .B2(
        i_data_bus[27]), .ZN(n147) );
  AOI22D1BWP30P140LVT U177 ( .A1(n183), .A2(i_data_bus[59]), .B1(n182), .B2(
        i_data_bus[123]), .ZN(n146) );
  AOI22D1BWP30P140LVT U178 ( .A1(n185), .A2(i_data_bus[219]), .B1(n184), .B2(
        i_data_bus[187]), .ZN(n145) );
  AOI22D1BWP30P140LVT U179 ( .A1(n186), .A2(i_data_bus[251]), .B1(n44), .B2(
        i_data_bus[91]), .ZN(n144) );
  ND4D1BWP30P140LVT U180 ( .A1(n147), .A2(n146), .A3(n145), .A4(n144), .ZN(
        N396) );
  AOI22D1BWP30P140LVT U181 ( .A1(n181), .A2(i_data_bus[154]), .B1(n180), .B2(
        i_data_bus[26]), .ZN(n151) );
  AOI22D1BWP30P140LVT U182 ( .A1(n183), .A2(i_data_bus[58]), .B1(n182), .B2(
        i_data_bus[122]), .ZN(n150) );
  AOI22D1BWP30P140LVT U183 ( .A1(n185), .A2(i_data_bus[218]), .B1(n184), .B2(
        i_data_bus[186]), .ZN(n149) );
  AOI22D1BWP30P140LVT U184 ( .A1(n186), .A2(i_data_bus[250]), .B1(n44), .B2(
        i_data_bus[90]), .ZN(n148) );
  ND4D1BWP30P140LVT U185 ( .A1(n151), .A2(n150), .A3(n149), .A4(n148), .ZN(
        N395) );
  AOI22D1BWP30P140LVT U186 ( .A1(n181), .A2(i_data_bus[153]), .B1(n180), .B2(
        i_data_bus[25]), .ZN(n155) );
  AOI22D1BWP30P140LVT U187 ( .A1(n183), .A2(i_data_bus[57]), .B1(n182), .B2(
        i_data_bus[121]), .ZN(n154) );
  AOI22D1BWP30P140LVT U188 ( .A1(n185), .A2(i_data_bus[217]), .B1(n184), .B2(
        i_data_bus[185]), .ZN(n153) );
  AOI22D1BWP30P140LVT U189 ( .A1(n186), .A2(i_data_bus[249]), .B1(n44), .B2(
        i_data_bus[89]), .ZN(n152) );
  ND4D1BWP30P140LVT U190 ( .A1(n155), .A2(n154), .A3(n153), .A4(n152), .ZN(
        N394) );
  AOI22D1BWP30P140LVT U191 ( .A1(n181), .A2(i_data_bus[151]), .B1(n180), .B2(
        i_data_bus[23]), .ZN(n159) );
  AOI22D1BWP30P140LVT U192 ( .A1(n183), .A2(i_data_bus[55]), .B1(n182), .B2(
        i_data_bus[119]), .ZN(n158) );
  AOI22D1BWP30P140LVT U193 ( .A1(n185), .A2(i_data_bus[215]), .B1(n184), .B2(
        i_data_bus[183]), .ZN(n157) );
  AOI22D1BWP30P140LVT U194 ( .A1(n186), .A2(i_data_bus[247]), .B1(n44), .B2(
        i_data_bus[87]), .ZN(n156) );
  ND4D1BWP30P140LVT U195 ( .A1(n159), .A2(n158), .A3(n157), .A4(n156), .ZN(
        N392) );
  AOI22D1BWP30P140LVT U196 ( .A1(n181), .A2(i_data_bus[150]), .B1(n180), .B2(
        i_data_bus[22]), .ZN(n163) );
  AOI22D1BWP30P140LVT U197 ( .A1(n183), .A2(i_data_bus[54]), .B1(n182), .B2(
        i_data_bus[118]), .ZN(n162) );
  AOI22D1BWP30P140LVT U198 ( .A1(n185), .A2(i_data_bus[214]), .B1(n184), .B2(
        i_data_bus[182]), .ZN(n161) );
  AOI22D1BWP30P140LVT U199 ( .A1(n186), .A2(i_data_bus[246]), .B1(n44), .B2(
        i_data_bus[86]), .ZN(n160) );
  ND4D1BWP30P140LVT U200 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .ZN(
        N391) );
  AOI22D1BWP30P140LVT U201 ( .A1(n181), .A2(i_data_bus[149]), .B1(n180), .B2(
        i_data_bus[21]), .ZN(n167) );
  AOI22D1BWP30P140LVT U202 ( .A1(n183), .A2(i_data_bus[53]), .B1(n182), .B2(
        i_data_bus[117]), .ZN(n166) );
  AOI22D1BWP30P140LVT U203 ( .A1(n185), .A2(i_data_bus[213]), .B1(n184), .B2(
        i_data_bus[181]), .ZN(n165) );
  AOI22D1BWP30P140LVT U204 ( .A1(n186), .A2(i_data_bus[245]), .B1(n44), .B2(
        i_data_bus[85]), .ZN(n164) );
  ND4D1BWP30P140LVT U205 ( .A1(n167), .A2(n166), .A3(n165), .A4(n164), .ZN(
        N390) );
  AOI22D1BWP30P140LVT U206 ( .A1(n181), .A2(i_data_bus[148]), .B1(n180), .B2(
        i_data_bus[20]), .ZN(n171) );
  AOI22D1BWP30P140LVT U207 ( .A1(n183), .A2(i_data_bus[52]), .B1(n182), .B2(
        i_data_bus[116]), .ZN(n170) );
  AOI22D1BWP30P140LVT U208 ( .A1(n185), .A2(i_data_bus[212]), .B1(n184), .B2(
        i_data_bus[180]), .ZN(n169) );
  AOI22D1BWP30P140LVT U209 ( .A1(n186), .A2(i_data_bus[244]), .B1(n44), .B2(
        i_data_bus[84]), .ZN(n168) );
  ND4D1BWP30P140LVT U210 ( .A1(n171), .A2(n170), .A3(n169), .A4(n168), .ZN(
        N389) );
  AOI22D1BWP30P140LVT U211 ( .A1(n181), .A2(i_data_bus[147]), .B1(n180), .B2(
        i_data_bus[19]), .ZN(n175) );
  AOI22D1BWP30P140LVT U212 ( .A1(n183), .A2(i_data_bus[51]), .B1(n182), .B2(
        i_data_bus[115]), .ZN(n174) );
  AOI22D1BWP30P140LVT U213 ( .A1(n185), .A2(i_data_bus[211]), .B1(n184), .B2(
        i_data_bus[179]), .ZN(n173) );
  AOI22D1BWP30P140LVT U214 ( .A1(n186), .A2(i_data_bus[243]), .B1(n44), .B2(
        i_data_bus[83]), .ZN(n172) );
  ND4D1BWP30P140LVT U215 ( .A1(n175), .A2(n174), .A3(n173), .A4(n172), .ZN(
        N388) );
  AOI22D1BWP30P140LVT U216 ( .A1(n181), .A2(i_data_bus[146]), .B1(n180), .B2(
        i_data_bus[18]), .ZN(n179) );
  AOI22D1BWP30P140LVT U217 ( .A1(n183), .A2(i_data_bus[50]), .B1(n182), .B2(
        i_data_bus[114]), .ZN(n178) );
  AOI22D1BWP30P140LVT U218 ( .A1(n185), .A2(i_data_bus[210]), .B1(n184), .B2(
        i_data_bus[178]), .ZN(n177) );
  AOI22D1BWP30P140LVT U219 ( .A1(n186), .A2(i_data_bus[242]), .B1(n44), .B2(
        i_data_bus[82]), .ZN(n176) );
  ND4D1BWP30P140LVT U220 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(
        N387) );
  AOI22D1BWP30P140LVT U221 ( .A1(n181), .A2(i_data_bus[145]), .B1(n180), .B2(
        i_data_bus[17]), .ZN(n190) );
  AOI22D1BWP30P140LVT U222 ( .A1(n183), .A2(i_data_bus[49]), .B1(n182), .B2(
        i_data_bus[113]), .ZN(n189) );
  AOI22D1BWP30P140LVT U223 ( .A1(n185), .A2(i_data_bus[209]), .B1(n184), .B2(
        i_data_bus[177]), .ZN(n188) );
  AOI22D1BWP30P140LVT U224 ( .A1(n186), .A2(i_data_bus[241]), .B1(n44), .B2(
        i_data_bus[81]), .ZN(n187) );
  ND4D1BWP30P140LVT U225 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(
        N386) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;
  tri   CLK;
  tri   rst;
  tri   i_en;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;
  tri   CLK;
  tri   rst;
  tri   i_en;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;
  tri   CLK;
  tri   rst;
  tri   i_en;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;
  tri   CLK;
  tri   rst;
  tri   i_en;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;
  tri   CLK;
  tri   rst;
  tri   i_en;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;
  tri   CLK;
  tri   rst;
  tri   i_en;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule



    module cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 ( 
        CLK, rst, o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, 
        o_cmd_6, o_cmd_7, i_en, i_cmd );
  input [7:0] i_cmd;
  input CLK, rst, i_en;
  output o_cmd_0, o_cmd_1, o_cmd_2, o_cmd_3, o_cmd_4, o_cmd_5, o_cmd_6,
         o_cmd_7;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;
  wire   [7:0] cmd_wire_0__inner_cmd_reg;
  wire   [7:0] cmd_wire_1__inner_cmd_reg;
  wire   [7:0] cmd_wire_2__inner_cmd_reg;
  tri   CLK;
  tri   rst;
  tri   i_en;

  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__7_ ( .D(N10), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__6_ ( .D(N9), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__5_ ( .D(N8), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__4_ ( .D(N7), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__3_ ( .D(N6), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__2_ ( .D(N5), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__1_ ( .D(N4), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_0__inner_cmd_reg_reg_0__0_ ( .D(N3), .CP(CLK), 
        .Q(cmd_wire_0__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__3_ ( .D(
        cmd_wire_0__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__2_ ( .D(
        cmd_wire_0__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_0__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_1__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_0__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_1__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[5]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[7]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_0__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[4]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[6]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[7]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[5]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_1__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[6]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[4]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[1]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[3]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_2__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[0]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[2]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__1_ ( .D(
        cmd_wire_1__inner_cmd_reg[3]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[1]) );
  DFQD1BWP30P140LVT cmd_wire_2__inner_cmd_reg_reg_3__0_ ( .D(
        cmd_wire_1__inner_cmd_reg[2]), .CP(CLK), .Q(
        cmd_wire_2__inner_cmd_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_2_ ( .D(cmd_wire_2__inner_cmd_reg[4]), .CP(
        CLK), .Q(o_cmd_2) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_7_ ( .D(cmd_wire_2__inner_cmd_reg[1]), .CP(
        CLK), .Q(o_cmd_7) );
  DFQD4BWP30P140LVT o_cmd_reg_reg_3_ ( .D(cmd_wire_2__inner_cmd_reg[5]), .CP(
        CLK), .Q(o_cmd_3) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_0_ ( .D(cmd_wire_2__inner_cmd_reg[6]), .CP(
        CLK), .Q(o_cmd_0) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_1_ ( .D(cmd_wire_2__inner_cmd_reg[7]), .CP(
        CLK), .Q(o_cmd_1) );
  DFQD1BWP30P140LVT o_cmd_reg_reg_4_ ( .D(cmd_wire_2__inner_cmd_reg[2]), .CP(
        CLK), .Q(o_cmd_4) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_5_ ( .D(cmd_wire_2__inner_cmd_reg[3]), .CP(
        CLK), .Q(o_cmd_5) );
  DFQD2BWP30P140LVT o_cmd_reg_reg_6_ ( .D(cmd_wire_2__inner_cmd_reg[0]), .CP(
        CLK), .Q(o_cmd_6) );
  INR2D1BWP30P140LVT U3 ( .A1(i_en), .B1(rst), .ZN(n1) );
  CKAN2D1BWP30P140LVT U4 ( .A1(n1), .A2(i_cmd[0]), .Z(N3) );
  CKAN2D1BWP30P140LVT U5 ( .A1(n1), .A2(i_cmd[1]), .Z(N4) );
  CKAN2D1BWP30P140LVT U6 ( .A1(n1), .A2(i_cmd[2]), .Z(N5) );
  CKAN2D1BWP30P140LVT U7 ( .A1(n1), .A2(i_cmd[3]), .Z(N6) );
  CKAN2D1BWP30P140LVT U8 ( .A1(n1), .A2(i_cmd[4]), .Z(N7) );
  CKAN2D1BWP30P140LVT U9 ( .A1(n1), .A2(i_cmd[5]), .Z(N8) );
  CKAN2D1BWP30P140LVT U10 ( .A1(n1), .A2(i_cmd[6]), .Z(N9) );
  CKAN2D1BWP30P140LVT U11 ( .A1(n1), .A2(i_cmd[7]), .Z(N10) );
endmodule


module crossbar_one_hot_seq ( CLK, rst, i_valid, i_data_bus, o_valid, 
        o_data_bus, i_en, i_cmd );
  input [7:0] i_valid;
  input [255:0] i_data_bus;
  output [7:0] o_valid;
  output [255:0] o_data_bus;
  input [63:0] i_cmd;
  input CLK, rst, i_en;
  wire   n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528;
  wire   [63:0] o_inner_cmd_wire;
  tri   CLK;
  tri   rst;
  tri   [7:0] i_valid;
  tri   [255:0] i_data_bus;
  tri   i_en;
  tri   [255:0] bottom_half_0__inner_data_i_mux_tree_wire;
  tri   [7:0] bottom_half_0__inner_valid_i_mux_tree_wire;
  tri   [255:0] bottom_half_1__inner_data_i_mux_tree_wire;
  tri   [7:0] bottom_half_1__inner_valid_i_mux_tree_wire;
  tri   [255:0] bottom_half_2__inner_data_i_mux_tree_wire;
  tri   [7:0] bottom_half_2__inner_valid_i_mux_tree_wire;
  tri   [255:0] bottom_half_3__inner_data_i_mux_tree_wire;
  tri   [7:0] bottom_half_3__inner_valid_i_mux_tree_wire;
  tri   [255:0] bottom_half_4__inner_data_i_mux_tree_wire;
  tri   [7:0] bottom_half_4__inner_valid_i_mux_tree_wire;
  tri   [255:0] bottom_half_5__inner_data_i_mux_tree_wire;
  tri   [7:0] bottom_half_5__inner_valid_i_mux_tree_wire;
  tri   [255:0] bottom_half_6__inner_data_i_mux_tree_wire;
  tri   [7:0] bottom_half_6__inner_valid_i_mux_tree_wire;
  tri   [255:0] bottom_half_7__inner_data_i_mux_tree_wire;
  tri   [7:0] bottom_half_7__inner_valid_i_mux_tree_wire;

  wire_binary_tree_1_8_seq top_half_0__wire_pipeline ( .CLK(CLK), .rst(rst), 
        .i_valid(i_valid[0]), .i_data_bus(i_data_bus[31:0]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[0], 
        bottom_half_6__inner_valid_i_mux_tree_wire[0], 
        bottom_half_5__inner_valid_i_mux_tree_wire[0], 
        bottom_half_4__inner_valid_i_mux_tree_wire[0], 
        bottom_half_3__inner_valid_i_mux_tree_wire[0], 
        bottom_half_2__inner_valid_i_mux_tree_wire[0], 
        bottom_half_1__inner_valid_i_mux_tree_wire[0], 
        bottom_half_0__inner_valid_i_mux_tree_wire[0]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_6__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_5__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_4__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_3__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_2__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_1__inner_data_i_mux_tree_wire[31:0], 
        bottom_half_0__inner_data_i_mux_tree_wire[31:0]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq top_half_1__wire_pipeline ( .CLK(CLK), .rst(rst), 
        .i_valid(i_valid[1]), .i_data_bus(i_data_bus[63:32]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[1], 
        bottom_half_6__inner_valid_i_mux_tree_wire[1], 
        bottom_half_5__inner_valid_i_mux_tree_wire[1], 
        bottom_half_4__inner_valid_i_mux_tree_wire[1], 
        bottom_half_3__inner_valid_i_mux_tree_wire[1], 
        bottom_half_2__inner_valid_i_mux_tree_wire[1], 
        bottom_half_1__inner_valid_i_mux_tree_wire[1], 
        bottom_half_0__inner_valid_i_mux_tree_wire[1]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_6__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_5__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_4__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_3__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_2__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_1__inner_data_i_mux_tree_wire[63:32], 
        bottom_half_0__inner_data_i_mux_tree_wire[63:32]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq top_half_2__wire_pipeline ( .CLK(CLK), .rst(rst), 
        .i_valid(i_valid[2]), .i_data_bus(i_data_bus[95:64]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[2], 
        bottom_half_6__inner_valid_i_mux_tree_wire[2], 
        bottom_half_5__inner_valid_i_mux_tree_wire[2], 
        bottom_half_4__inner_valid_i_mux_tree_wire[2], 
        bottom_half_3__inner_valid_i_mux_tree_wire[2], 
        bottom_half_2__inner_valid_i_mux_tree_wire[2], 
        bottom_half_1__inner_valid_i_mux_tree_wire[2], 
        bottom_half_0__inner_valid_i_mux_tree_wire[2]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_6__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_5__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_4__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_3__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_2__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_1__inner_data_i_mux_tree_wire[95:64], 
        bottom_half_0__inner_data_i_mux_tree_wire[95:64]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq top_half_3__wire_pipeline ( .CLK(CLK), .rst(rst), 
        .i_valid(i_valid[3]), .i_data_bus(i_data_bus[127:96]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[3], 
        bottom_half_6__inner_valid_i_mux_tree_wire[3], 
        bottom_half_5__inner_valid_i_mux_tree_wire[3], 
        bottom_half_4__inner_valid_i_mux_tree_wire[3], 
        bottom_half_3__inner_valid_i_mux_tree_wire[3], 
        bottom_half_2__inner_valid_i_mux_tree_wire[3], 
        bottom_half_1__inner_valid_i_mux_tree_wire[3], 
        bottom_half_0__inner_valid_i_mux_tree_wire[3]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_6__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_5__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_4__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_3__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_2__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_1__inner_data_i_mux_tree_wire[127:96], 
        bottom_half_0__inner_data_i_mux_tree_wire[127:96]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq top_half_4__wire_pipeline ( .CLK(CLK), .rst(rst), 
        .i_valid(i_valid[4]), .i_data_bus(i_data_bus[159:128]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[4], 
        bottom_half_6__inner_valid_i_mux_tree_wire[4], 
        bottom_half_5__inner_valid_i_mux_tree_wire[4], 
        bottom_half_4__inner_valid_i_mux_tree_wire[4], 
        bottom_half_3__inner_valid_i_mux_tree_wire[4], 
        bottom_half_2__inner_valid_i_mux_tree_wire[4], 
        bottom_half_1__inner_valid_i_mux_tree_wire[4], 
        bottom_half_0__inner_valid_i_mux_tree_wire[4]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_6__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_5__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_4__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_3__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_2__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_1__inner_data_i_mux_tree_wire[159:128], 
        bottom_half_0__inner_data_i_mux_tree_wire[159:128]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq top_half_5__wire_pipeline ( .CLK(CLK), .rst(rst), 
        .i_valid(i_valid[5]), .i_data_bus(i_data_bus[191:160]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[5], 
        bottom_half_6__inner_valid_i_mux_tree_wire[5], 
        bottom_half_5__inner_valid_i_mux_tree_wire[5], 
        bottom_half_4__inner_valid_i_mux_tree_wire[5], 
        bottom_half_3__inner_valid_i_mux_tree_wire[5], 
        bottom_half_2__inner_valid_i_mux_tree_wire[5], 
        bottom_half_1__inner_valid_i_mux_tree_wire[5], 
        bottom_half_0__inner_valid_i_mux_tree_wire[5]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_6__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_5__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_4__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_3__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_2__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_1__inner_data_i_mux_tree_wire[191:160], 
        bottom_half_0__inner_data_i_mux_tree_wire[191:160]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq top_half_6__wire_pipeline ( .CLK(CLK), .rst(rst), 
        .i_valid(i_valid[6]), .i_data_bus(i_data_bus[223:192]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[6], 
        bottom_half_6__inner_valid_i_mux_tree_wire[6], 
        bottom_half_5__inner_valid_i_mux_tree_wire[6], 
        bottom_half_4__inner_valid_i_mux_tree_wire[6], 
        bottom_half_3__inner_valid_i_mux_tree_wire[6], 
        bottom_half_2__inner_valid_i_mux_tree_wire[6], 
        bottom_half_1__inner_valid_i_mux_tree_wire[6], 
        bottom_half_0__inner_valid_i_mux_tree_wire[6]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_6__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_5__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_4__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_3__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_2__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_1__inner_data_i_mux_tree_wire[223:192], 
        bottom_half_0__inner_data_i_mux_tree_wire[223:192]}), .i_en(i_en) );
  wire_binary_tree_1_8_seq top_half_7__wire_pipeline ( .CLK(CLK), .rst(rst), 
        .i_valid(i_valid[7]), .i_data_bus(i_data_bus[255:224]), .o_valid({
        bottom_half_7__inner_valid_i_mux_tree_wire[7], 
        bottom_half_6__inner_valid_i_mux_tree_wire[7], 
        bottom_half_5__inner_valid_i_mux_tree_wire[7], 
        bottom_half_4__inner_valid_i_mux_tree_wire[7], 
        bottom_half_3__inner_valid_i_mux_tree_wire[7], 
        bottom_half_2__inner_valid_i_mux_tree_wire[7], 
        bottom_half_1__inner_valid_i_mux_tree_wire[7], 
        bottom_half_0__inner_valid_i_mux_tree_wire[7]}), .o_data_bus({
        bottom_half_7__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_6__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_5__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_4__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_3__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_2__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_1__inner_data_i_mux_tree_wire[255:224], 
        bottom_half_0__inner_data_i_mux_tree_wire[255:224]}), .i_en(i_en) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_0 i_cmd_id_0__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[0]), .o_cmd_1(
        o_inner_cmd_wire[8]), .o_cmd_2(o_inner_cmd_wire[16]), .o_cmd_3(
        o_inner_cmd_wire[24]), .o_cmd_4(o_inner_cmd_wire[32]), .o_cmd_5(
        o_inner_cmd_wire[40]), .o_cmd_6(o_inner_cmd_wire[48]), .o_cmd_7(
        o_inner_cmd_wire[56]), .i_en(i_en), .i_cmd(i_cmd[7:0]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_7 i_cmd_id_1__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[1]), .o_cmd_1(
        o_inner_cmd_wire[9]), .o_cmd_2(o_inner_cmd_wire[17]), .o_cmd_3(
        o_inner_cmd_wire[25]), .o_cmd_4(o_inner_cmd_wire[33]), .o_cmd_5(
        o_inner_cmd_wire[41]), .o_cmd_6(o_inner_cmd_wire[49]), .o_cmd_7(
        o_inner_cmd_wire[57]), .i_en(i_en), .i_cmd(i_cmd[15:8]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_6 i_cmd_id_2__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[2]), .o_cmd_1(
        o_inner_cmd_wire[10]), .o_cmd_2(o_inner_cmd_wire[18]), .o_cmd_3(
        o_inner_cmd_wire[26]), .o_cmd_4(o_inner_cmd_wire[34]), .o_cmd_5(
        o_inner_cmd_wire[42]), .o_cmd_6(o_inner_cmd_wire[50]), .o_cmd_7(
        o_inner_cmd_wire[58]), .i_en(i_en), .i_cmd(i_cmd[23:16]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_5 i_cmd_id_3__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[3]), .o_cmd_1(
        o_inner_cmd_wire[11]), .o_cmd_2(o_inner_cmd_wire[19]), .o_cmd_3(
        o_inner_cmd_wire[27]), .o_cmd_4(o_inner_cmd_wire[35]), .o_cmd_5(
        o_inner_cmd_wire[43]), .o_cmd_6(o_inner_cmd_wire[51]), .o_cmd_7(
        o_inner_cmd_wire[59]), .i_en(i_en), .i_cmd(i_cmd[31:24]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_4 i_cmd_id_4__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[4]), .o_cmd_1(
        o_inner_cmd_wire[12]), .o_cmd_2(o_inner_cmd_wire[20]), .o_cmd_3(
        o_inner_cmd_wire[28]), .o_cmd_4(o_inner_cmd_wire[36]), .o_cmd_5(
        o_inner_cmd_wire[44]), .o_cmd_6(o_inner_cmd_wire[52]), .o_cmd_7(
        o_inner_cmd_wire[60]), .i_en(i_en), .i_cmd(i_cmd[39:32]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_3 i_cmd_id_5__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[5]), .o_cmd_1(
        o_inner_cmd_wire[13]), .o_cmd_2(o_inner_cmd_wire[21]), .o_cmd_3(
        o_inner_cmd_wire[29]), .o_cmd_4(o_inner_cmd_wire[37]), .o_cmd_5(
        o_inner_cmd_wire[45]), .o_cmd_6(o_inner_cmd_wire[53]), .o_cmd_7(
        o_inner_cmd_wire[61]), .i_en(i_en), .i_cmd(i_cmd[47:40]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_2 i_cmd_id_6__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[6]), .o_cmd_1(
        o_inner_cmd_wire[14]), .o_cmd_2(o_inner_cmd_wire[22]), .o_cmd_3(
        o_inner_cmd_wire[30]), .o_cmd_4(o_inner_cmd_wire[38]), .o_cmd_5(
        o_inner_cmd_wire[46]), .o_cmd_6(o_inner_cmd_wire[54]), .o_cmd_7(
        o_inner_cmd_wire[62]), .i_en(i_en), .i_cmd(i_cmd[55:48]) );
  cmd_wire_binary_tree_1_8_seq_DATA_WIDTH32_NUM_OUTPUT_DATA8_NUM_INPUT_DATA1_1 i_cmd_id_7__cmd_pipeline ( 
        .CLK(CLK), .rst(rst), .o_cmd_0(o_inner_cmd_wire[7]), .o_cmd_1(
        o_inner_cmd_wire[15]), .o_cmd_2(o_inner_cmd_wire[23]), .o_cmd_3(
        o_inner_cmd_wire[31]), .o_cmd_4(o_inner_cmd_wire[39]), .o_cmd_5(
        o_inner_cmd_wire[47]), .o_cmd_6(o_inner_cmd_wire[55]), .o_cmd_7(
        o_inner_cmd_wire[63]), .i_en(i_en), .i_cmd(i_cmd[63:56]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_0 bottom_half_0__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_0__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_0__inner_data_i_mux_tree_wire), .o_valid(n272), 
        .o_data_bus({n497, n498, n499, n500, n501, n502, n503, n504, n505, 
        n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
        n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[7:0]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_7 bottom_half_1__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_1__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_1__inner_data_i_mux_tree_wire), .o_valid(n271), 
        .o_data_bus({n465, n466, n467, n468, n469, n470, n471, n472, n473, 
        n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, 
        n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[15:8]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_6 bottom_half_2__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_2__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_2__inner_data_i_mux_tree_wire), .o_valid(n270), 
        .o_data_bus({n433, n434, n435, n436, n437, n438, n439, n440, n441, 
        n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
        n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[23:16]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_5 bottom_half_3__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_3__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_3__inner_data_i_mux_tree_wire), .o_valid(n269), 
        .o_data_bus({n401, n402, n403, n404, n405, n406, n407, n408, n409, 
        n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
        n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[31:24]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_4 bottom_half_4__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_4__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_4__inner_data_i_mux_tree_wire), .o_valid(n268), 
        .o_data_bus({n369, n370, n371, n372, n373, n374, n375, n376, n377, 
        n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
        n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[39:32]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_3 bottom_half_5__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_5__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_5__inner_data_i_mux_tree_wire), .o_valid(n267), 
        .o_data_bus({n337, n338, n339, n340, n341, n342, n343, n344, n345, 
        n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
        n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[47:40]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_2 bottom_half_6__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_6__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_6__inner_data_i_mux_tree_wire), .o_valid(n266), 
        .o_data_bus({n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[55:48]) );
  mux_tree_8_1_seq_DATA_WIDTH32_NUM_OUTPUT_DATA1_NUM_INPUT_DATA8_1 bottom_half_7__mux_tree ( 
        .CLK(CLK), .rst(rst), .i_valid(
        bottom_half_7__inner_valid_i_mux_tree_wire), .i_data_bus(
        bottom_half_7__inner_data_i_mux_tree_wire), .o_valid(n265), 
        .o_data_bus({n273, n274, n275, n276, n277, n278, n279, n280, n281, 
        n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
        n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304}), 
        .i_en(i_en), .i_cmd(o_inner_cmd_wire[63:56]) );
  BUFFD6BWP30P140LVT U1 ( .I(n528), .Z(o_data_bus[0]) );
  BUFFD6BWP30P140LVT U2 ( .I(n527), .Z(o_data_bus[1]) );
  BUFFD6BWP30P140LVT U3 ( .I(n526), .Z(o_data_bus[2]) );
  BUFFD6BWP30P140LVT U4 ( .I(n525), .Z(o_data_bus[3]) );
  BUFFD6BWP30P140LVT U5 ( .I(n524), .Z(o_data_bus[4]) );
  BUFFD6BWP30P140LVT U6 ( .I(n523), .Z(o_data_bus[5]) );
  BUFFD6BWP30P140LVT U7 ( .I(n522), .Z(o_data_bus[6]) );
  BUFFD6BWP30P140LVT U8 ( .I(n521), .Z(o_data_bus[7]) );
  BUFFD6BWP30P140LVT U9 ( .I(n520), .Z(o_data_bus[8]) );
  BUFFD6BWP30P140LVT U10 ( .I(n519), .Z(o_data_bus[9]) );
  BUFFD6BWP30P140LVT U11 ( .I(n518), .Z(o_data_bus[10]) );
  BUFFD6BWP30P140LVT U12 ( .I(n517), .Z(o_data_bus[11]) );
  BUFFD6BWP30P140LVT U13 ( .I(n516), .Z(o_data_bus[12]) );
  BUFFD6BWP30P140LVT U14 ( .I(n515), .Z(o_data_bus[13]) );
  BUFFD6BWP30P140LVT U15 ( .I(n514), .Z(o_data_bus[14]) );
  BUFFD6BWP30P140LVT U16 ( .I(n513), .Z(o_data_bus[15]) );
  BUFFD6BWP30P140LVT U17 ( .I(n512), .Z(o_data_bus[16]) );
  BUFFD6BWP30P140LVT U18 ( .I(n511), .Z(o_data_bus[17]) );
  BUFFD6BWP30P140LVT U19 ( .I(n510), .Z(o_data_bus[18]) );
  BUFFD6BWP30P140LVT U20 ( .I(n509), .Z(o_data_bus[19]) );
  BUFFD6BWP30P140LVT U21 ( .I(n508), .Z(o_data_bus[20]) );
  BUFFD6BWP30P140LVT U22 ( .I(n507), .Z(o_data_bus[21]) );
  BUFFD6BWP30P140LVT U23 ( .I(n506), .Z(o_data_bus[22]) );
  BUFFD6BWP30P140LVT U24 ( .I(n505), .Z(o_data_bus[23]) );
  BUFFD6BWP30P140LVT U25 ( .I(n504), .Z(o_data_bus[24]) );
  BUFFD6BWP30P140LVT U26 ( .I(n503), .Z(o_data_bus[25]) );
  BUFFD6BWP30P140LVT U27 ( .I(n502), .Z(o_data_bus[26]) );
  BUFFD6BWP30P140LVT U28 ( .I(n501), .Z(o_data_bus[27]) );
  BUFFD6BWP30P140LVT U29 ( .I(n500), .Z(o_data_bus[28]) );
  BUFFD6BWP30P140LVT U30 ( .I(n499), .Z(o_data_bus[29]) );
  BUFFD6BWP30P140LVT U31 ( .I(n498), .Z(o_data_bus[30]) );
  BUFFD6BWP30P140LVT U32 ( .I(n497), .Z(o_data_bus[31]) );
  BUFFD6BWP30P140LVT U33 ( .I(n496), .Z(o_data_bus[32]) );
  BUFFD6BWP30P140LVT U34 ( .I(n495), .Z(o_data_bus[33]) );
  BUFFD6BWP30P140LVT U35 ( .I(n494), .Z(o_data_bus[34]) );
  BUFFD6BWP30P140LVT U36 ( .I(n493), .Z(o_data_bus[35]) );
  BUFFD6BWP30P140LVT U37 ( .I(n492), .Z(o_data_bus[36]) );
  BUFFD6BWP30P140LVT U38 ( .I(n491), .Z(o_data_bus[37]) );
  BUFFD6BWP30P140LVT U39 ( .I(n490), .Z(o_data_bus[38]) );
  BUFFD6BWP30P140LVT U40 ( .I(n489), .Z(o_data_bus[39]) );
  BUFFD6BWP30P140LVT U41 ( .I(n488), .Z(o_data_bus[40]) );
  BUFFD6BWP30P140LVT U42 ( .I(n487), .Z(o_data_bus[41]) );
  BUFFD6BWP30P140LVT U43 ( .I(n486), .Z(o_data_bus[42]) );
  BUFFD6BWP30P140LVT U44 ( .I(n485), .Z(o_data_bus[43]) );
  BUFFD6BWP30P140LVT U45 ( .I(n484), .Z(o_data_bus[44]) );
  BUFFD6BWP30P140LVT U46 ( .I(n483), .Z(o_data_bus[45]) );
  BUFFD6BWP30P140LVT U47 ( .I(n482), .Z(o_data_bus[46]) );
  BUFFD6BWP30P140LVT U48 ( .I(n481), .Z(o_data_bus[47]) );
  BUFFD6BWP30P140LVT U49 ( .I(n480), .Z(o_data_bus[48]) );
  BUFFD6BWP30P140LVT U50 ( .I(n479), .Z(o_data_bus[49]) );
  BUFFD6BWP30P140LVT U51 ( .I(n478), .Z(o_data_bus[50]) );
  BUFFD6BWP30P140LVT U52 ( .I(n477), .Z(o_data_bus[51]) );
  BUFFD6BWP30P140LVT U53 ( .I(n476), .Z(o_data_bus[52]) );
  BUFFD6BWP30P140LVT U54 ( .I(n475), .Z(o_data_bus[53]) );
  BUFFD6BWP30P140LVT U55 ( .I(n474), .Z(o_data_bus[54]) );
  BUFFD6BWP30P140LVT U56 ( .I(n473), .Z(o_data_bus[55]) );
  BUFFD6BWP30P140LVT U57 ( .I(n472), .Z(o_data_bus[56]) );
  BUFFD6BWP30P140LVT U58 ( .I(n471), .Z(o_data_bus[57]) );
  BUFFD6BWP30P140LVT U59 ( .I(n470), .Z(o_data_bus[58]) );
  BUFFD6BWP30P140LVT U60 ( .I(n469), .Z(o_data_bus[59]) );
  BUFFD6BWP30P140LVT U61 ( .I(n468), .Z(o_data_bus[60]) );
  BUFFD6BWP30P140LVT U62 ( .I(n467), .Z(o_data_bus[61]) );
  BUFFD6BWP30P140LVT U63 ( .I(n466), .Z(o_data_bus[62]) );
  BUFFD6BWP30P140LVT U64 ( .I(n465), .Z(o_data_bus[63]) );
  BUFFD6BWP30P140LVT U65 ( .I(n464), .Z(o_data_bus[64]) );
  BUFFD6BWP30P140LVT U66 ( .I(n463), .Z(o_data_bus[65]) );
  BUFFD6BWP30P140LVT U67 ( .I(n462), .Z(o_data_bus[66]) );
  BUFFD6BWP30P140LVT U68 ( .I(n461), .Z(o_data_bus[67]) );
  BUFFD6BWP30P140LVT U69 ( .I(n460), .Z(o_data_bus[68]) );
  BUFFD6BWP30P140LVT U70 ( .I(n459), .Z(o_data_bus[69]) );
  BUFFD6BWP30P140LVT U71 ( .I(n458), .Z(o_data_bus[70]) );
  BUFFD6BWP30P140LVT U72 ( .I(n457), .Z(o_data_bus[71]) );
  BUFFD6BWP30P140LVT U73 ( .I(n456), .Z(o_data_bus[72]) );
  BUFFD6BWP30P140LVT U74 ( .I(n455), .Z(o_data_bus[73]) );
  BUFFD6BWP30P140LVT U75 ( .I(n454), .Z(o_data_bus[74]) );
  BUFFD6BWP30P140LVT U76 ( .I(n453), .Z(o_data_bus[75]) );
  BUFFD6BWP30P140LVT U77 ( .I(n452), .Z(o_data_bus[76]) );
  BUFFD6BWP30P140LVT U78 ( .I(n451), .Z(o_data_bus[77]) );
  BUFFD6BWP30P140LVT U79 ( .I(n450), .Z(o_data_bus[78]) );
  BUFFD6BWP30P140LVT U80 ( .I(n449), .Z(o_data_bus[79]) );
  BUFFD6BWP30P140LVT U81 ( .I(n448), .Z(o_data_bus[80]) );
  BUFFD6BWP30P140LVT U82 ( .I(n447), .Z(o_data_bus[81]) );
  BUFFD6BWP30P140LVT U83 ( .I(n446), .Z(o_data_bus[82]) );
  BUFFD6BWP30P140LVT U84 ( .I(n445), .Z(o_data_bus[83]) );
  BUFFD6BWP30P140LVT U85 ( .I(n444), .Z(o_data_bus[84]) );
  BUFFD6BWP30P140LVT U86 ( .I(n443), .Z(o_data_bus[85]) );
  BUFFD6BWP30P140LVT U87 ( .I(n442), .Z(o_data_bus[86]) );
  BUFFD6BWP30P140LVT U88 ( .I(n441), .Z(o_data_bus[87]) );
  BUFFD6BWP30P140LVT U89 ( .I(n440), .Z(o_data_bus[88]) );
  BUFFD6BWP30P140LVT U90 ( .I(n439), .Z(o_data_bus[89]) );
  BUFFD6BWP30P140LVT U91 ( .I(n438), .Z(o_data_bus[90]) );
  BUFFD6BWP30P140LVT U92 ( .I(n437), .Z(o_data_bus[91]) );
  BUFFD6BWP30P140LVT U93 ( .I(n436), .Z(o_data_bus[92]) );
  BUFFD6BWP30P140LVT U94 ( .I(n435), .Z(o_data_bus[93]) );
  BUFFD6BWP30P140LVT U95 ( .I(n434), .Z(o_data_bus[94]) );
  BUFFD6BWP30P140LVT U96 ( .I(n433), .Z(o_data_bus[95]) );
  BUFFD6BWP30P140LVT U97 ( .I(n432), .Z(o_data_bus[96]) );
  BUFFD6BWP30P140LVT U98 ( .I(n431), .Z(o_data_bus[97]) );
  BUFFD6BWP30P140LVT U99 ( .I(n430), .Z(o_data_bus[98]) );
  BUFFD6BWP30P140LVT U100 ( .I(n429), .Z(o_data_bus[99]) );
  BUFFD6BWP30P140LVT U101 ( .I(n428), .Z(o_data_bus[100]) );
  BUFFD6BWP30P140LVT U102 ( .I(n427), .Z(o_data_bus[101]) );
  BUFFD6BWP30P140LVT U103 ( .I(n426), .Z(o_data_bus[102]) );
  BUFFD6BWP30P140LVT U104 ( .I(n425), .Z(o_data_bus[103]) );
  BUFFD6BWP30P140LVT U105 ( .I(n424), .Z(o_data_bus[104]) );
  BUFFD6BWP30P140LVT U106 ( .I(n423), .Z(o_data_bus[105]) );
  BUFFD6BWP30P140LVT U107 ( .I(n422), .Z(o_data_bus[106]) );
  BUFFD6BWP30P140LVT U108 ( .I(n421), .Z(o_data_bus[107]) );
  BUFFD6BWP30P140LVT U109 ( .I(n420), .Z(o_data_bus[108]) );
  BUFFD6BWP30P140LVT U110 ( .I(n419), .Z(o_data_bus[109]) );
  BUFFD6BWP30P140LVT U111 ( .I(n418), .Z(o_data_bus[110]) );
  BUFFD6BWP30P140LVT U112 ( .I(n417), .Z(o_data_bus[111]) );
  BUFFD6BWP30P140LVT U113 ( .I(n416), .Z(o_data_bus[112]) );
  BUFFD6BWP30P140LVT U114 ( .I(n415), .Z(o_data_bus[113]) );
  BUFFD6BWP30P140LVT U115 ( .I(n414), .Z(o_data_bus[114]) );
  BUFFD6BWP30P140LVT U116 ( .I(n413), .Z(o_data_bus[115]) );
  BUFFD6BWP30P140LVT U117 ( .I(n412), .Z(o_data_bus[116]) );
  BUFFD6BWP30P140LVT U118 ( .I(n411), .Z(o_data_bus[117]) );
  BUFFD6BWP30P140LVT U119 ( .I(n410), .Z(o_data_bus[118]) );
  BUFFD6BWP30P140LVT U120 ( .I(n409), .Z(o_data_bus[119]) );
  BUFFD6BWP30P140LVT U121 ( .I(n408), .Z(o_data_bus[120]) );
  BUFFD6BWP30P140LVT U122 ( .I(n407), .Z(o_data_bus[121]) );
  BUFFD6BWP30P140LVT U123 ( .I(n406), .Z(o_data_bus[122]) );
  BUFFD6BWP30P140LVT U124 ( .I(n405), .Z(o_data_bus[123]) );
  BUFFD6BWP30P140LVT U125 ( .I(n404), .Z(o_data_bus[124]) );
  BUFFD6BWP30P140LVT U126 ( .I(n403), .Z(o_data_bus[125]) );
  BUFFD6BWP30P140LVT U127 ( .I(n402), .Z(o_data_bus[126]) );
  BUFFD6BWP30P140LVT U128 ( .I(n401), .Z(o_data_bus[127]) );
  BUFFD6BWP30P140LVT U129 ( .I(n400), .Z(o_data_bus[128]) );
  BUFFD6BWP30P140LVT U130 ( .I(n399), .Z(o_data_bus[129]) );
  BUFFD6BWP30P140LVT U131 ( .I(n398), .Z(o_data_bus[130]) );
  BUFFD6BWP30P140LVT U132 ( .I(n397), .Z(o_data_bus[131]) );
  BUFFD6BWP30P140LVT U133 ( .I(n396), .Z(o_data_bus[132]) );
  BUFFD6BWP30P140LVT U134 ( .I(n395), .Z(o_data_bus[133]) );
  BUFFD6BWP30P140LVT U135 ( .I(n394), .Z(o_data_bus[134]) );
  BUFFD6BWP30P140LVT U136 ( .I(n393), .Z(o_data_bus[135]) );
  BUFFD6BWP30P140LVT U137 ( .I(n392), .Z(o_data_bus[136]) );
  BUFFD6BWP30P140LVT U138 ( .I(n391), .Z(o_data_bus[137]) );
  BUFFD6BWP30P140LVT U139 ( .I(n390), .Z(o_data_bus[138]) );
  BUFFD6BWP30P140LVT U140 ( .I(n389), .Z(o_data_bus[139]) );
  BUFFD6BWP30P140LVT U141 ( .I(n388), .Z(o_data_bus[140]) );
  BUFFD6BWP30P140LVT U142 ( .I(n387), .Z(o_data_bus[141]) );
  BUFFD6BWP30P140LVT U143 ( .I(n386), .Z(o_data_bus[142]) );
  BUFFD6BWP30P140LVT U144 ( .I(n385), .Z(o_data_bus[143]) );
  BUFFD6BWP30P140LVT U145 ( .I(n384), .Z(o_data_bus[144]) );
  BUFFD6BWP30P140LVT U146 ( .I(n383), .Z(o_data_bus[145]) );
  BUFFD6BWP30P140LVT U147 ( .I(n382), .Z(o_data_bus[146]) );
  BUFFD6BWP30P140LVT U148 ( .I(n381), .Z(o_data_bus[147]) );
  BUFFD6BWP30P140LVT U149 ( .I(n380), .Z(o_data_bus[148]) );
  BUFFD6BWP30P140LVT U150 ( .I(n379), .Z(o_data_bus[149]) );
  BUFFD6BWP30P140LVT U151 ( .I(n378), .Z(o_data_bus[150]) );
  BUFFD6BWP30P140LVT U152 ( .I(n377), .Z(o_data_bus[151]) );
  BUFFD6BWP30P140LVT U153 ( .I(n376), .Z(o_data_bus[152]) );
  BUFFD6BWP30P140LVT U154 ( .I(n375), .Z(o_data_bus[153]) );
  BUFFD6BWP30P140LVT U155 ( .I(n374), .Z(o_data_bus[154]) );
  BUFFD6BWP30P140LVT U156 ( .I(n373), .Z(o_data_bus[155]) );
  BUFFD6BWP30P140LVT U157 ( .I(n372), .Z(o_data_bus[156]) );
  BUFFD6BWP30P140LVT U158 ( .I(n371), .Z(o_data_bus[157]) );
  BUFFD6BWP30P140LVT U159 ( .I(n370), .Z(o_data_bus[158]) );
  BUFFD6BWP30P140LVT U160 ( .I(n369), .Z(o_data_bus[159]) );
  BUFFD6BWP30P140LVT U161 ( .I(n368), .Z(o_data_bus[160]) );
  BUFFD6BWP30P140LVT U162 ( .I(n367), .Z(o_data_bus[161]) );
  BUFFD6BWP30P140LVT U163 ( .I(n366), .Z(o_data_bus[162]) );
  BUFFD6BWP30P140LVT U164 ( .I(n365), .Z(o_data_bus[163]) );
  BUFFD6BWP30P140LVT U165 ( .I(n364), .Z(o_data_bus[164]) );
  BUFFD6BWP30P140LVT U166 ( .I(n363), .Z(o_data_bus[165]) );
  BUFFD6BWP30P140LVT U167 ( .I(n362), .Z(o_data_bus[166]) );
  BUFFD6BWP30P140LVT U168 ( .I(n361), .Z(o_data_bus[167]) );
  BUFFD6BWP30P140LVT U169 ( .I(n360), .Z(o_data_bus[168]) );
  BUFFD6BWP30P140LVT U170 ( .I(n359), .Z(o_data_bus[169]) );
  BUFFD6BWP30P140LVT U171 ( .I(n358), .Z(o_data_bus[170]) );
  BUFFD6BWP30P140LVT U172 ( .I(n357), .Z(o_data_bus[171]) );
  BUFFD6BWP30P140LVT U173 ( .I(n356), .Z(o_data_bus[172]) );
  BUFFD6BWP30P140LVT U174 ( .I(n355), .Z(o_data_bus[173]) );
  BUFFD6BWP30P140LVT U175 ( .I(n354), .Z(o_data_bus[174]) );
  BUFFD6BWP30P140LVT U176 ( .I(n353), .Z(o_data_bus[175]) );
  BUFFD6BWP30P140LVT U177 ( .I(n352), .Z(o_data_bus[176]) );
  BUFFD6BWP30P140LVT U178 ( .I(n351), .Z(o_data_bus[177]) );
  BUFFD6BWP30P140LVT U179 ( .I(n350), .Z(o_data_bus[178]) );
  BUFFD6BWP30P140LVT U180 ( .I(n349), .Z(o_data_bus[179]) );
  BUFFD6BWP30P140LVT U181 ( .I(n348), .Z(o_data_bus[180]) );
  BUFFD6BWP30P140LVT U182 ( .I(n347), .Z(o_data_bus[181]) );
  BUFFD6BWP30P140LVT U183 ( .I(n346), .Z(o_data_bus[182]) );
  BUFFD6BWP30P140LVT U184 ( .I(n345), .Z(o_data_bus[183]) );
  BUFFD6BWP30P140LVT U185 ( .I(n344), .Z(o_data_bus[184]) );
  BUFFD6BWP30P140LVT U186 ( .I(n343), .Z(o_data_bus[185]) );
  BUFFD6BWP30P140LVT U187 ( .I(n342), .Z(o_data_bus[186]) );
  BUFFD6BWP30P140LVT U188 ( .I(n341), .Z(o_data_bus[187]) );
  BUFFD6BWP30P140LVT U189 ( .I(n340), .Z(o_data_bus[188]) );
  BUFFD6BWP30P140LVT U190 ( .I(n339), .Z(o_data_bus[189]) );
  BUFFD6BWP30P140LVT U191 ( .I(n338), .Z(o_data_bus[190]) );
  BUFFD6BWP30P140LVT U192 ( .I(n337), .Z(o_data_bus[191]) );
  BUFFD6BWP30P140LVT U193 ( .I(n336), .Z(o_data_bus[192]) );
  BUFFD6BWP30P140LVT U194 ( .I(n335), .Z(o_data_bus[193]) );
  BUFFD6BWP30P140LVT U195 ( .I(n334), .Z(o_data_bus[194]) );
  BUFFD6BWP30P140LVT U196 ( .I(n333), .Z(o_data_bus[195]) );
  BUFFD6BWP30P140LVT U197 ( .I(n332), .Z(o_data_bus[196]) );
  BUFFD6BWP30P140LVT U198 ( .I(n331), .Z(o_data_bus[197]) );
  BUFFD6BWP30P140LVT U199 ( .I(n330), .Z(o_data_bus[198]) );
  BUFFD6BWP30P140LVT U200 ( .I(n329), .Z(o_data_bus[199]) );
  BUFFD6BWP30P140LVT U201 ( .I(n328), .Z(o_data_bus[200]) );
  BUFFD6BWP30P140LVT U202 ( .I(n327), .Z(o_data_bus[201]) );
  BUFFD6BWP30P140LVT U203 ( .I(n326), .Z(o_data_bus[202]) );
  BUFFD6BWP30P140LVT U204 ( .I(n325), .Z(o_data_bus[203]) );
  BUFFD6BWP30P140LVT U205 ( .I(n324), .Z(o_data_bus[204]) );
  BUFFD6BWP30P140LVT U206 ( .I(n323), .Z(o_data_bus[205]) );
  BUFFD6BWP30P140LVT U207 ( .I(n322), .Z(o_data_bus[206]) );
  BUFFD6BWP30P140LVT U208 ( .I(n321), .Z(o_data_bus[207]) );
  BUFFD6BWP30P140LVT U209 ( .I(n320), .Z(o_data_bus[208]) );
  BUFFD6BWP30P140LVT U210 ( .I(n319), .Z(o_data_bus[209]) );
  BUFFD6BWP30P140LVT U211 ( .I(n318), .Z(o_data_bus[210]) );
  BUFFD6BWP30P140LVT U212 ( .I(n317), .Z(o_data_bus[211]) );
  BUFFD6BWP30P140LVT U213 ( .I(n316), .Z(o_data_bus[212]) );
  BUFFD6BWP30P140LVT U214 ( .I(n315), .Z(o_data_bus[213]) );
  BUFFD6BWP30P140LVT U215 ( .I(n314), .Z(o_data_bus[214]) );
  BUFFD6BWP30P140LVT U216 ( .I(n313), .Z(o_data_bus[215]) );
  BUFFD6BWP30P140LVT U217 ( .I(n312), .Z(o_data_bus[216]) );
  BUFFD6BWP30P140LVT U218 ( .I(n311), .Z(o_data_bus[217]) );
  BUFFD6BWP30P140LVT U219 ( .I(n310), .Z(o_data_bus[218]) );
  BUFFD6BWP30P140LVT U220 ( .I(n309), .Z(o_data_bus[219]) );
  BUFFD6BWP30P140LVT U221 ( .I(n308), .Z(o_data_bus[220]) );
  BUFFD6BWP30P140LVT U222 ( .I(n307), .Z(o_data_bus[221]) );
  BUFFD6BWP30P140LVT U223 ( .I(n306), .Z(o_data_bus[222]) );
  BUFFD6BWP30P140LVT U224 ( .I(n305), .Z(o_data_bus[223]) );
  BUFFD6BWP30P140LVT U225 ( .I(n304), .Z(o_data_bus[224]) );
  BUFFD6BWP30P140LVT U226 ( .I(n303), .Z(o_data_bus[225]) );
  BUFFD6BWP30P140LVT U227 ( .I(n302), .Z(o_data_bus[226]) );
  BUFFD6BWP30P140LVT U228 ( .I(n301), .Z(o_data_bus[227]) );
  BUFFD6BWP30P140LVT U229 ( .I(n300), .Z(o_data_bus[228]) );
  BUFFD6BWP30P140LVT U230 ( .I(n299), .Z(o_data_bus[229]) );
  BUFFD6BWP30P140LVT U231 ( .I(n298), .Z(o_data_bus[230]) );
  BUFFD6BWP30P140LVT U232 ( .I(n297), .Z(o_data_bus[231]) );
  BUFFD6BWP30P140LVT U233 ( .I(n296), .Z(o_data_bus[232]) );
  BUFFD6BWP30P140LVT U234 ( .I(n295), .Z(o_data_bus[233]) );
  BUFFD6BWP30P140LVT U235 ( .I(n294), .Z(o_data_bus[234]) );
  BUFFD6BWP30P140LVT U236 ( .I(n293), .Z(o_data_bus[235]) );
  BUFFD6BWP30P140LVT U237 ( .I(n292), .Z(o_data_bus[236]) );
  BUFFD6BWP30P140LVT U238 ( .I(n291), .Z(o_data_bus[237]) );
  BUFFD6BWP30P140LVT U239 ( .I(n290), .Z(o_data_bus[238]) );
  BUFFD6BWP30P140LVT U240 ( .I(n289), .Z(o_data_bus[239]) );
  BUFFD6BWP30P140LVT U241 ( .I(n288), .Z(o_data_bus[240]) );
  BUFFD6BWP30P140LVT U242 ( .I(n287), .Z(o_data_bus[241]) );
  BUFFD6BWP30P140LVT U243 ( .I(n286), .Z(o_data_bus[242]) );
  BUFFD6BWP30P140LVT U244 ( .I(n285), .Z(o_data_bus[243]) );
  BUFFD6BWP30P140LVT U245 ( .I(n284), .Z(o_data_bus[244]) );
  BUFFD6BWP30P140LVT U246 ( .I(n283), .Z(o_data_bus[245]) );
  BUFFD6BWP30P140LVT U247 ( .I(n282), .Z(o_data_bus[246]) );
  BUFFD6BWP30P140LVT U248 ( .I(n281), .Z(o_data_bus[247]) );
  BUFFD6BWP30P140LVT U249 ( .I(n280), .Z(o_data_bus[248]) );
  BUFFD6BWP30P140LVT U250 ( .I(n279), .Z(o_data_bus[249]) );
  BUFFD6BWP30P140LVT U251 ( .I(n278), .Z(o_data_bus[250]) );
  BUFFD6BWP30P140LVT U252 ( .I(n277), .Z(o_data_bus[251]) );
  BUFFD6BWP30P140LVT U253 ( .I(n276), .Z(o_data_bus[252]) );
  BUFFD6BWP30P140LVT U254 ( .I(n275), .Z(o_data_bus[253]) );
  BUFFD6BWP30P140LVT U255 ( .I(n274), .Z(o_data_bus[254]) );
  BUFFD6BWP30P140LVT U256 ( .I(n273), .Z(o_data_bus[255]) );
  BUFFD6BWP30P140LVT U257 ( .I(n272), .Z(o_valid[0]) );
  BUFFD6BWP30P140LVT U258 ( .I(n271), .Z(o_valid[1]) );
  BUFFD6BWP30P140LVT U259 ( .I(n270), .Z(o_valid[2]) );
  BUFFD6BWP30P140LVT U260 ( .I(n269), .Z(o_valid[3]) );
  BUFFD6BWP30P140LVT U261 ( .I(n268), .Z(o_valid[4]) );
  BUFFD6BWP30P140LVT U262 ( .I(n267), .Z(o_valid[5]) );
  BUFFD6BWP30P140LVT U263 ( .I(n266), .Z(o_valid[6]) );
  BUFFD6BWP30P140LVT U264 ( .I(n265), .Z(o_valid[7]) );
endmodule

