`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module controller_integrated(CLK, reset, boot_up, start, table_parse, input_valid, glob_scen_noc_input_valid, delay_matrix_element, obj_id_element,from_glob_prefetch_start,  from_glob_prefetch_dest,  scenario_update, local_controller_id, tapping_loc_packet, from_glob_prefetch_stop, hardware_latency1, hardware_latency2, scenario_len, prefetch_bypass_dest_addr_int, prefetch_bypass_cycles, prefetch_bypass_start_addr, addr, data_in, prefetch_bypass_path_input_data,prefetch_bypass_path_input_addr, prefetch_bypass_valid, packet_out_0, packet_out_1, packet_out_2, packet_out_3, from_glob_prefetch_valid, from_glob_prefetch_start_0, from_glob_prefetch_start_1, from_glob_prefetch_start_2, from_glob_prefetch_start_3, from_glob_prefetch_stop_0, from_glob_prefetch_stop_1, from_glob_prefetch_stop_2, from_glob_prefetch_stop_3, from_glob_prefetch_dest_0, from_glob_prefetch_dest_1, from_glob_prefetch_dest_2, from_glob_prefetch_dest_3, from_glob_prefetch_valid0, from_glob_prefetch_valid1, from_glob_prefetch_valid2, from_glob_prefetch_valid3);

    // parameter
    	parameter N_sample = 256;
	parameter datawidth = 16;
	parameter address_vector_width = 4; //can be 200 or 8: 8 for small tapeout
	parameter N_obj = 4; //can be 200 or 8: 8 for small tapeout
	parameter id_width = 6; // 16 local controllers in subscaled system
	parameter sample_address_width = 8; /// assuming 256 words: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	parameter delay_length = 14; // log(id_width*N_sample)
	parameter obj_id_width = 2; // log(N_obj)
	parameter tapping_loc_packet_width = sample_address_width + obj_id_width; // log(N_obj)
	parameter scen_len_width = 11;   //needs to be revised
	

//=== IO Ports ===//

     // Normal Mode Input
    	input CLK; // system clock, generated by VCO
	input reset;
	input start;
	input boot_up;
	input table_parse;
	input input_valid;
	input glob_scen_noc_input_valid;
	input [delay_length - 1:0] delay_matrix_element;
	input [obj_id_width - 1:0] obj_id_element;
	input scenario_update;
	input [delay_length - 1:0] hardware_latency1;   ///keep as config to be input through spi?
	input [delay_length - 1:0] hardware_latency2;   /// keep as config to be input through spi?
	input [scen_len_width - 1:0] scenario_len;   /// keep as config to be input through spi?
	input [2*datawidth - 1:0] data_in;   /// keep as config to be input through spi?

/////// to be removed finally /////////////////////////////////////
	input [sample_address_width - 1:0] from_glob_prefetch_start_0;
	input [sample_address_width - 1:0] from_glob_prefetch_start_1;
	input [sample_address_width - 1:0] from_glob_prefetch_start_2;
	input [sample_address_width - 1:0] from_glob_prefetch_start_3;
	input [sample_address_width - 1:0] from_glob_prefetch_stop_0;
	input [sample_address_width - 1:0] from_glob_prefetch_stop_1;
	input [sample_address_width - 1:0] from_glob_prefetch_stop_2;
	input [sample_address_width - 1:0] from_glob_prefetch_stop_3;
	input [address_vector_width - 1:0] from_glob_prefetch_dest_0;
	input [address_vector_width - 1:0] from_glob_prefetch_dest_1;
	input [address_vector_width - 1:0] from_glob_prefetch_dest_2;
	input [address_vector_width - 1:0] from_glob_prefetch_dest_3;

	input from_glob_prefetch_valid0;
	input from_glob_prefetch_valid1;
	input from_glob_prefetch_valid2;
	input from_glob_prefetch_valid3;

    // output
	output [address_vector_width - 1:0] from_glob_prefetch_dest;
	output [sample_address_width - 1:0] from_glob_prefetch_start;
	output [sample_address_width - 1:0] from_glob_prefetch_stop;
	output [id_width - 1:0] local_controller_id;
	output [tapping_loc_packet_width - 1:0] tapping_loc_packet;
	output [address_vector_width - 1:0] prefetch_bypass_dest_addr_int;
	output [sample_address_width - 1:0] prefetch_bypass_cycles;
	output [delay_length - 1:0] prefetch_bypass_start_addr;

	output [id_width - 1:0] addr;
	output [2*datawidth - 1:0] prefetch_bypass_path_input_data;
	output [address_vector_width - 1:0] prefetch_bypass_path_input_addr;
	output prefetch_bypass_valid;

        output [packet_width-1:0] packet_out_0;   
        output [packet_width-1:0] packet_out_1;   
        output [packet_width-1:0] packet_out_2;   
        output [packet_width-1:0] packet_out_3;   




//////////// internal status regs/signals //////////////////////////////////
	wire [2*datawidth - 1:0] h_tree_input_data;
	wire [id_width - 1:0] h_tree_input_addr;

	wire write_flag_0;
	wire write_flag_1;
	wire write_flag_2;
	wire write_flag_3;

	wire boundary_next_0;
	wire boundary_next_1;
	wire boundary_next_2;
	wire boundary_next_3;
	wire [address_vector_width - 1:0] dest_address_0;
	wire [address_vector_width - 1:0] dest_address_1;
	wire [address_vector_width - 1:0] dest_address_2;
	wire [address_vector_width - 1:0] dest_address_3;


	wire [sample_address_width - 1:0] prefetch_stop_address_0;
	wire [sample_address_width - 1:0] prefetch_stop_address_1;
	wire [sample_address_width - 1:0] prefetch_stop_address_2;
	wire [sample_address_width - 1:0] prefetch_stop_address_3;
	wire [address_vector_width - 1:0] prefetch_dest_addr_0;
	wire [address_vector_width - 1:0] prefetch_dest_addr_1;
	wire [address_vector_width - 1:0] prefetch_dest_addr_2;
	wire [address_vector_width - 1:0] prefetch_dest_addr_3;
	wire prefetch_boundary_prev_0;
	wire prefetch_boundary_prev_1;
	wire prefetch_boundary_prev_2;
	wire prefetch_boundary_prev_3;

	wire [2*datawidth - 1:0] D_0;
	wire [2*datawidth - 1:0] D_1;
	wire [2*datawidth - 1:0] D_2;
	wire [2*datawidth - 1:0] D_3;

////////// to be removed ///////////////////////

	wire write_boundary_next_0;
	wire write_boundary_next_1;
	wire write_boundary_next_2;
	wire write_boundary_next_3;


////////// logic part /////////////////////////////////////////////////////// 
 
////////////sequential logic

    global_controller DUT_global_controller(.CLK(CLK), .reset(reset), .start(start), .boot_up(boot_up),  .table_parse(table_parse), .input_valid(input_valid), .glob_scen_noc_input_valid(glob_scen_noc_input_valid), .delay_matrix_element(delay_matrix_element), .obj_id_element(obj_id_element),.from_glob_prefetch_start(from_glob_prefetch_start),.from_glob_prefetch_dest(from_glob_prefetch_dest),  .scenario_update(scenario_update), .local_controller_id(local_controller_id), .tapping_loc_packet(tapping_loc_packet), .from_glob_prefetch_stop(from_glob_prefetch_stop), .hardware_latency1(hardware_latency1), .hardware_latency2(hardware_latency2), .scenario_len(scenario_len), .prefetch_bypass_dest_addr_int(prefetch_bypass_dest_addr_int), .prefetch_bypass_cycles(prefetch_bypass_cycles), .prefetch_bypass_start_addr(prefetch_bypass_start_addr), .addr(addr), .data_in(data_in), .h_tree_input_data(h_tree_input_data), .h_tree_input_addr(h_tree_input_addr), .prefetch_bypass_path_input_data(prefetch_bypass_path_input_data), .prefetch_bypass_path_input_addr(prefetch_bypass_path_input_addr), .prefetch_bypass_valid(prefetch_bypass_valid));

    Htree_Flat DUT_htree( .CLK(CLK), .addr(h_tree_input_addr), .en(start), .data_in(h_tree_input_data),  .en_sub_0(write_flag_0), .en_sub_1(write_flag_1), .en_sub_2(write_flag_2), .en_sub_3(write_flag_3), .data_in_sub_0(D_0), .data_in_sub_1(D_1), .data_in_sub_2(D_2), .data_in_sub_3(D_3));

 
    local_controller_prefetch_full DUT_local_controller_0(.CLK(CLK), .reset(reset), .boot_up(boot_up), .start(start),     .input_boundary_flag(boundary_next_3), .prev_dest_address(dest_address_3),.packet_out(packet_out_0), .boundary_next(boundary_next_0), .dest_address(dest_address_0), .D(D_0),.write_flag(write_flag_0), .from_glob_prefetch_valid(from_glob_prefetch_valid0), .from_glob_prefetch_start(from_glob_prefetch_start_0), .from_glob_prefetch_stop(from_glob_prefetch_stop_0), .from_glob_prefetch_dest(from_glob_prefetch_dest_0),  .write_boundary_next(write_boundary_next_0), .input_write_boundary(write_boundary_next_3), .prefetch_next_dest_addr(prefetch_dest_addr_1), .prefetch_next_stop_address(prefetch_stop_address_1), .prefetch_boundary_prev(prefetch_boundary_prev_0), .input_prefetch_boundary_flag(prefetch_boundary_prev_1), .prefetch_stop_address(prefetch_stop_address_0), .prefetch_dest_addr(prefetch_dest_addr_0),.scenario_update(scenario_update));

    local_controller_prefetch_full DUT_local_controller_1(.CLK(CLK), .reset(reset),   .boot_up(boot_up), .start(start),     .input_boundary_flag(boundary_next_0), .prev_dest_address(dest_address_0), .packet_out(packet_out_1), .boundary_next(boundary_next_1), .dest_address(dest_address_1), .D(D_1),  .write_flag(write_flag_1), .from_glob_prefetch_valid(from_glob_prefetch_valid1), .from_glob_prefetch_start(from_glob_prefetch_start_1), .from_glob_prefetch_stop(from_glob_prefetch_stop_1), .from_glob_prefetch_dest(from_glob_prefetch_dest_1),   .write_boundary_next(write_boundary_next_1), .input_write_boundary(write_boundary_next_0), .prefetch_next_dest_addr(prefetch_dest_addr_2), .prefetch_next_stop_address(prefetch_stop_address_2), .prefetch_boundary_prev(prefetch_boundary_prev_1), .input_prefetch_boundary_flag(prefetch_boundary_prev_2), .prefetch_stop_address(prefetch_stop_address_1), .prefetch_dest_addr(prefetch_dest_addr_1), .scenario_update(scenario_update));

    local_controller_prefetch_full DUT_local_controller_2(.CLK(CLK), .reset(reset),   .boot_up(boot_up), .start(start),    .input_boundary_flag(boundary_next_1), .prev_dest_address(dest_address_1), .packet_out(packet_out_2), .boundary_next(boundary_next_2), .dest_address(dest_address_2), .D(D_2), .write_flag(write_flag_2), .from_glob_prefetch_valid(from_glob_prefetch_valid2), .from_glob_prefetch_start(from_glob_prefetch_start_2), .from_glob_prefetch_stop(from_glob_prefetch_stop_2), .from_glob_prefetch_dest(from_glob_prefetch_dest_2),  .write_boundary_next(write_boundary_next_2), .input_write_boundary(write_boundary_next_1), .prefetch_next_dest_addr(prefetch_dest_addr_3), .prefetch_next_stop_address(prefetch_stop_address_3), .prefetch_boundary_prev(prefetch_boundary_prev_2), .input_prefetch_boundary_flag(prefetch_boundary_prev_3), .prefetch_stop_address(prefetch_stop_address_2), .prefetch_dest_addr(prefetch_dest_addr_2),  .scenario_update(scenario_update));

    local_controller_prefetch_full DUT_local_controller_3(.CLK(CLK), .reset(reset),   .boot_up(boot_up), .start(start),   .input_boundary_flag(boundary_next_2), .prev_dest_address(dest_address_2),  .packet_out(packet_out_3), .boundary_next(boundary_next_3), .dest_address(dest_address_3), .D(D_3),  .write_flag(write_flag_3), .from_glob_prefetch_valid(from_glob_prefetch_valid3), .from_glob_prefetch_start(from_glob_prefetch_start_3), .from_glob_prefetch_stop(from_glob_prefetch_stop_3), .from_glob_prefetch_dest(from_glob_prefetch_dest_3),  .write_boundary_next(write_boundary_next_3), .input_write_boundary(write_boundary_next_2), .prefetch_next_dest_addr(prefetch_dest_addr_0), .prefetch_next_stop_address(prefetch_stop_address_0), .prefetch_boundary_prev(prefetch_boundary_prev_3), .input_prefetch_boundary_flag(prefetch_boundary_prev_0), .prefetch_stop_address(prefetch_stop_address_3), .prefetch_dest_addr(prefetch_dest_addr_3),  .scenario_update(scenario_update));



	 
	 


   
endmodule
    

