`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Gatech	
// Engineer: Mandovi Mukherjee
// 
// Create Date: 01/08/2021 
// System Name: accelerator
// Module Name: local controller
// Project Name: ARION DRBE
// Description: fetch and push data out to network; assuming the output from
// global controller comes in the form of a packet
// Dependencies:
// Additional Comments: 
/////////////////////////////////////////////////////////////////////////////////////////////////////

module local_controller_simple_negedge(clk, reset, init,  boundary_next );
    // parameter
    parameter N_row = 1024;
	parameter datawidth = 32;
	parameter address_vector_width = 8; //can be 200 or 8: 8 for subscaled system
	parameter id_width = 11; // 1221 local controllers in subscaled system
	parameter row_address_width = 10; /// assuming 1024 rows and 64 columns: needs to change if arrangement is different
	parameter packet_width = 2*datawidth + address_vector_width;
	
	
	
        
    // input
    input clk; // system clock, generated by VCO
	input reset;
	input init;
	input glob_controller_sending; //not used
	input [2*datawidth - 1:0] data_from_sram;
	input [id_width - 1:0] controller_id;
	input input_boundary_flag;
	input write_flag;
	input [address_vector_width - 1:0] prev_dest_address;
	input [address_vector_width - 1:0] from_glob_dest_addr;
	input [row_address_width - 1:0] from_glob_controller_delay;
	input scenario_end_flag;

    // output
    output [packet_width-1:0] packet_out;  
    output reg boundary_next;
    output reg [address_vector_width - 1:0] dest_address;
	
	

    // internal status regs/signals
    reg [row_address_width-1:0] row_address;
	reg [id_width - 1:0] id; 
	reg [packet_width-1:0] packet_out_internal;
	reg coeff_num;
	reg [row_address_width - 1:0] delay;
    

    // logic part  
    assign packet_out = packet_out_internal;


	//sequential logic
	 
	 
	 always @ (posedge clk) begin
		boundary_next <= 0;
		if (reset) begin
			coeff_num <= coeff_num;
			row_address <= row_address;
			dest_address <= dest_address;
		end
		else if (input_boundary_flag == 1) begin
			coeff_num <= 1;
			row_address <= 0;
			dest_address <= prev_dest_address;
		end
		else if (input_boundary_flag == 0) begin
			if (boundary_next == 1) begin
				coeff_num <= 0;
			end
			else begin
				coeff_num <= coeff_num;
			end
			row_address <= row_address;
			dest_address <= dest_address;
			
		end
	 end
	 
	 


   
endmodule
    
