
module linear_network_unicast_seq_1_16 ( CLK, rst, i_valid, i_data_bus, 
        o_valid, o_data_bus, i_en, i_cmd );
  input [24:0] i_data_bus;
  output [15:0] o_valid;
  output [399:0] o_data_bus;
  input [3:0] i_cmd;
  input CLK, rst, i_valid, i_en;
  wire   N155, N156, N157, N158, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N264, N265, N266, N320, N321, N322, N323, N324, N325, N326, N327,
         N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338,
         N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349,
         N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360,
         N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371,
         N373, N374, N453, N454, N455, N456, N457, N458, N459, N460, N461,
         N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, N481, N482, N536, N537,
         N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548,
         N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559,
         N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570,
         N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581,
         N582, N583, N584, N585, N586, N587, N588, N590, N644, N645, N646,
         N647, N648, N649, N650, N651, N652, N653, N654, N655, N656, N657,
         N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668,
         N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679,
         N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690,
         N691, N692, N693, N694, N696, N697, N698, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N805, N806, N860, N861, N862, N863, N864, N865, N866, N867,
         N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878,
         N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889,
         N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900,
         N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911,
         N912, N914, N968, N969, N970, N971, N972, N973, N974, N975, N976,
         N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987,
         N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998,
         N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008,
         N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018,
         N1019, N1020, N1021, N1076, N1077, N1078, N1079, N1080, N1081, N1082,
         N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092,
         N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102,
         N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112,
         N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122,
         N1123, N1124, N1125, N1126, N1128, N1129, N1130, N1209, N1210, N1211,
         N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221,
         N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231,
         N1232, N1233, N1234, N1235, N1236, N1237, N1292, N1293, N1294, N1295,
         N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304, N1305,
         N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315,
         N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325,
         N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335,
         N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1345, N1346,
         N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434,
         N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444,
         N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1508,
         N1509, N1510, N1511, N1512, N1513, N1514, N1515, N1516, N1517, N1518,
         N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528,
         N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538,
         N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548,
         N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558,
         N1559, N1560, N1561, N1616, N1617, N1618, N1619, N1620, N1621, N1622,
         N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632,
         N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642,
         N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652,
         N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662,
         N1663, N1664, N1665, N1666, N1667, N1668, N1670, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259;
  wire   [374:0] o_data_forward_reg;
  wire   [0:14] o_valid_forward_reg;
  wire   [59:0] o_cmd_forward_reg;

  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__3_ ( .D(N158), .CP(CLK), .Q(
        o_cmd_forward_reg[59]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__2_ ( .D(N157), .CP(CLK), .Q(
        o_cmd_forward_reg[58]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__1_ ( .D(N156), .CP(CLK), .Q(
        o_cmd_forward_reg[57]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_0__0_ ( .D(N155), .CP(CLK), .Q(
        o_cmd_forward_reg[56]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__24_ ( .D(n202), .CP(CLK), .Q(
        o_data_forward_reg[374]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__23_ ( .D(n201), .CP(CLK), .Q(
        o_data_forward_reg[373]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__22_ ( .D(n200), .CP(CLK), .Q(
        o_data_forward_reg[372]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__21_ ( .D(n199), .CP(CLK), .Q(
        o_data_forward_reg[371]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__20_ ( .D(n198), .CP(CLK), .Q(
        o_data_forward_reg[370]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__19_ ( .D(n197), .CP(CLK), .Q(
        o_data_forward_reg[369]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__18_ ( .D(n196), .CP(CLK), .Q(
        o_data_forward_reg[368]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__17_ ( .D(n195), .CP(CLK), .Q(
        o_data_forward_reg[367]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__16_ ( .D(n194), .CP(CLK), .Q(
        o_data_forward_reg[366]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__15_ ( .D(n193), .CP(CLK), .Q(
        o_data_forward_reg[365]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__14_ ( .D(n192), .CP(CLK), .Q(
        o_data_forward_reg[364]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__13_ ( .D(n191), .CP(CLK), .Q(
        o_data_forward_reg[363]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__12_ ( .D(n190), .CP(CLK), .Q(
        o_data_forward_reg[362]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__11_ ( .D(n189), .CP(CLK), .Q(
        o_data_forward_reg[361]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__10_ ( .D(n188), .CP(CLK), .Q(
        o_data_forward_reg[360]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__9_ ( .D(n187), .CP(CLK), .Q(
        o_data_forward_reg[359]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__8_ ( .D(n186), .CP(CLK), .Q(
        o_data_forward_reg[358]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__7_ ( .D(n185), .CP(CLK), .Q(
        o_data_forward_reg[357]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__6_ ( .D(n184), .CP(CLK), .Q(
        o_data_forward_reg[356]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__5_ ( .D(n183), .CP(CLK), .Q(
        o_data_forward_reg[355]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__4_ ( .D(n182), .CP(CLK), .Q(
        o_data_forward_reg[354]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__3_ ( .D(n181), .CP(CLK), .Q(
        o_data_forward_reg[353]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__2_ ( .D(n180), .CP(CLK), .Q(
        o_data_forward_reg[352]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__1_ ( .D(n179), .CP(CLK), .Q(
        o_data_forward_reg[351]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_0__0_ ( .D(n178), .CP(CLK), .Q(
        o_data_forward_reg[350]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_0_ ( .D(n250), .CP(CLK), .Q(
        o_valid_forward_reg[0]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__3_ ( .D(N266), .CP(CLK), .Q(
        o_cmd_forward_reg[55]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__2_ ( .D(N265), .CP(CLK), .Q(
        o_cmd_forward_reg[54]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__1_ ( .D(N264), .CP(CLK), .Q(
        o_cmd_forward_reg[53]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_1__0_ ( .D(n251), .CP(CLK), .Q(
        o_cmd_forward_reg[52]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__24_ ( .D(N261), .CP(CLK), .Q(
        o_data_forward_reg[349]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__23_ ( .D(N260), .CP(CLK), .Q(
        o_data_forward_reg[348]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__22_ ( .D(N259), .CP(CLK), .Q(
        o_data_forward_reg[347]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__21_ ( .D(N258), .CP(CLK), .Q(
        o_data_forward_reg[346]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__20_ ( .D(N257), .CP(CLK), .Q(
        o_data_forward_reg[345]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__19_ ( .D(N256), .CP(CLK), .Q(
        o_data_forward_reg[344]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__18_ ( .D(N255), .CP(CLK), .Q(
        o_data_forward_reg[343]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__17_ ( .D(N254), .CP(CLK), .Q(
        o_data_forward_reg[342]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__16_ ( .D(N253), .CP(CLK), .Q(
        o_data_forward_reg[341]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__15_ ( .D(N252), .CP(CLK), .Q(
        o_data_forward_reg[340]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__14_ ( .D(N251), .CP(CLK), .Q(
        o_data_forward_reg[339]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__13_ ( .D(N250), .CP(CLK), .Q(
        o_data_forward_reg[338]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__12_ ( .D(N249), .CP(CLK), .Q(
        o_data_forward_reg[337]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__11_ ( .D(N248), .CP(CLK), .Q(
        o_data_forward_reg[336]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__10_ ( .D(N247), .CP(CLK), .Q(
        o_data_forward_reg[335]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__9_ ( .D(N246), .CP(CLK), .Q(
        o_data_forward_reg[334]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__8_ ( .D(N245), .CP(CLK), .Q(
        o_data_forward_reg[333]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__7_ ( .D(N244), .CP(CLK), .Q(
        o_data_forward_reg[332]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__6_ ( .D(N243), .CP(CLK), .Q(
        o_data_forward_reg[331]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__5_ ( .D(N242), .CP(CLK), .Q(
        o_data_forward_reg[330]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__4_ ( .D(N241), .CP(CLK), .Q(
        o_data_forward_reg[329]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__3_ ( .D(N240), .CP(CLK), .Q(
        o_data_forward_reg[328]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__2_ ( .D(N239), .CP(CLK), .Q(
        o_data_forward_reg[327]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__1_ ( .D(N238), .CP(CLK), .Q(
        o_data_forward_reg[326]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_1__0_ ( .D(N237), .CP(CLK), .Q(
        o_data_forward_reg[325]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_1_ ( .D(N262), .CP(CLK), .Q(
        o_valid_forward_reg[1]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__3_ ( .D(N374), .CP(CLK), .Q(
        o_cmd_forward_reg[51]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__2_ ( .D(N373), .CP(CLK), .Q(
        o_cmd_forward_reg[50]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__1_ ( .D(n249), .CP(CLK), .Q(
        o_cmd_forward_reg[49]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_2__0_ ( .D(N371), .CP(CLK), .Q(
        o_cmd_forward_reg[48]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__24_ ( .D(N369), .CP(CLK), .Q(
        o_data_forward_reg[324]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__23_ ( .D(N368), .CP(CLK), .Q(
        o_data_forward_reg[323]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__22_ ( .D(N367), .CP(CLK), .Q(
        o_data_forward_reg[322]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__21_ ( .D(N366), .CP(CLK), .Q(
        o_data_forward_reg[321]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__20_ ( .D(N365), .CP(CLK), .Q(
        o_data_forward_reg[320]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__19_ ( .D(N364), .CP(CLK), .Q(
        o_data_forward_reg[319]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__18_ ( .D(N363), .CP(CLK), .Q(
        o_data_forward_reg[318]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__17_ ( .D(N362), .CP(CLK), .Q(
        o_data_forward_reg[317]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__16_ ( .D(N361), .CP(CLK), .Q(
        o_data_forward_reg[316]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__15_ ( .D(N360), .CP(CLK), .Q(
        o_data_forward_reg[315]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__14_ ( .D(N359), .CP(CLK), .Q(
        o_data_forward_reg[314]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__13_ ( .D(N358), .CP(CLK), .Q(
        o_data_forward_reg[313]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__12_ ( .D(N357), .CP(CLK), .Q(
        o_data_forward_reg[312]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__11_ ( .D(N356), .CP(CLK), .Q(
        o_data_forward_reg[311]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__10_ ( .D(N355), .CP(CLK), .Q(
        o_data_forward_reg[310]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__9_ ( .D(N354), .CP(CLK), .Q(
        o_data_forward_reg[309]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__8_ ( .D(N353), .CP(CLK), .Q(
        o_data_forward_reg[308]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__7_ ( .D(N352), .CP(CLK), .Q(
        o_data_forward_reg[307]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__6_ ( .D(N351), .CP(CLK), .Q(
        o_data_forward_reg[306]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__5_ ( .D(N350), .CP(CLK), .Q(
        o_data_forward_reg[305]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__4_ ( .D(N349), .CP(CLK), .Q(
        o_data_forward_reg[304]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__3_ ( .D(N348), .CP(CLK), .Q(
        o_data_forward_reg[303]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__2_ ( .D(N347), .CP(CLK), .Q(
        o_data_forward_reg[302]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__1_ ( .D(N346), .CP(CLK), .Q(
        o_data_forward_reg[301]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_2__0_ ( .D(N345), .CP(CLK), .Q(
        o_data_forward_reg[300]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_2_ ( .D(N370), .CP(CLK), .Q(
        o_valid_forward_reg[2]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_3__3_ ( .D(N482), .CP(CLK), .Q(
        o_cmd_forward_reg[47]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_3__2_ ( .D(N481), .CP(CLK), .Q(
        o_cmd_forward_reg[46]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_3__1_ ( .D(n252), .CP(CLK), .Q(
        o_cmd_forward_reg[45]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_3__0_ ( .D(N479), .CP(CLK), .Q(
        o_cmd_forward_reg[44]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__24_ ( .D(N477), .CP(CLK), .Q(
        o_data_forward_reg[299]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__23_ ( .D(N476), .CP(CLK), .Q(
        o_data_forward_reg[298]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__22_ ( .D(N475), .CP(CLK), .Q(
        o_data_forward_reg[297]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__21_ ( .D(N474), .CP(CLK), .Q(
        o_data_forward_reg[296]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__20_ ( .D(N473), .CP(CLK), .Q(
        o_data_forward_reg[295]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__19_ ( .D(N472), .CP(CLK), .Q(
        o_data_forward_reg[294]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__18_ ( .D(N471), .CP(CLK), .Q(
        o_data_forward_reg[293]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__17_ ( .D(N470), .CP(CLK), .Q(
        o_data_forward_reg[292]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__16_ ( .D(N469), .CP(CLK), .Q(
        o_data_forward_reg[291]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__15_ ( .D(N468), .CP(CLK), .Q(
        o_data_forward_reg[290]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__14_ ( .D(N467), .CP(CLK), .Q(
        o_data_forward_reg[289]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__13_ ( .D(N466), .CP(CLK), .Q(
        o_data_forward_reg[288]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__12_ ( .D(N465), .CP(CLK), .Q(
        o_data_forward_reg[287]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__11_ ( .D(N464), .CP(CLK), .Q(
        o_data_forward_reg[286]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__10_ ( .D(N463), .CP(CLK), .Q(
        o_data_forward_reg[285]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__9_ ( .D(N462), .CP(CLK), .Q(
        o_data_forward_reg[284]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__8_ ( .D(N461), .CP(CLK), .Q(
        o_data_forward_reg[283]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__7_ ( .D(N460), .CP(CLK), .Q(
        o_data_forward_reg[282]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__6_ ( .D(N459), .CP(CLK), .Q(
        o_data_forward_reg[281]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__5_ ( .D(N458), .CP(CLK), .Q(
        o_data_forward_reg[280]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__4_ ( .D(N457), .CP(CLK), .Q(
        o_data_forward_reg[279]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__3_ ( .D(N456), .CP(CLK), .Q(
        o_data_forward_reg[278]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__2_ ( .D(N455), .CP(CLK), .Q(
        o_data_forward_reg[277]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__1_ ( .D(N454), .CP(CLK), .Q(
        o_data_forward_reg[276]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_3__0_ ( .D(N453), .CP(CLK), .Q(
        o_data_forward_reg[275]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_3_ ( .D(N478), .CP(CLK), .Q(
        o_valid_forward_reg[3]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_4__3_ ( .D(N590), .CP(CLK), .Q(
        o_cmd_forward_reg[43]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_4__2_ ( .D(n248), .CP(CLK), .Q(
        o_cmd_forward_reg[42]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_4__1_ ( .D(N588), .CP(CLK), .Q(
        o_cmd_forward_reg[41]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_4__0_ ( .D(N587), .CP(CLK), .Q(
        o_cmd_forward_reg[40]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__24_ ( .D(N585), .CP(CLK), .Q(
        o_data_forward_reg[274]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__23_ ( .D(N584), .CP(CLK), .Q(
        o_data_forward_reg[273]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__22_ ( .D(N583), .CP(CLK), .Q(
        o_data_forward_reg[272]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__21_ ( .D(N582), .CP(CLK), .Q(
        o_data_forward_reg[271]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__20_ ( .D(N581), .CP(CLK), .Q(
        o_data_forward_reg[270]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__19_ ( .D(N580), .CP(CLK), .Q(
        o_data_forward_reg[269]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__18_ ( .D(N579), .CP(CLK), .Q(
        o_data_forward_reg[268]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__17_ ( .D(N578), .CP(CLK), .Q(
        o_data_forward_reg[267]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__16_ ( .D(N577), .CP(CLK), .Q(
        o_data_forward_reg[266]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__15_ ( .D(N576), .CP(CLK), .Q(
        o_data_forward_reg[265]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__14_ ( .D(N575), .CP(CLK), .Q(
        o_data_forward_reg[264]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__13_ ( .D(N574), .CP(CLK), .Q(
        o_data_forward_reg[263]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__12_ ( .D(N573), .CP(CLK), .Q(
        o_data_forward_reg[262]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__11_ ( .D(N572), .CP(CLK), .Q(
        o_data_forward_reg[261]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__10_ ( .D(N571), .CP(CLK), .Q(
        o_data_forward_reg[260]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__9_ ( .D(N570), .CP(CLK), .Q(
        o_data_forward_reg[259]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__8_ ( .D(N569), .CP(CLK), .Q(
        o_data_forward_reg[258]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__7_ ( .D(N568), .CP(CLK), .Q(
        o_data_forward_reg[257]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__6_ ( .D(N567), .CP(CLK), .Q(
        o_data_forward_reg[256]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__5_ ( .D(N566), .CP(CLK), .Q(
        o_data_forward_reg[255]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__4_ ( .D(N565), .CP(CLK), .Q(
        o_data_forward_reg[254]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__3_ ( .D(N564), .CP(CLK), .Q(
        o_data_forward_reg[253]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__2_ ( .D(N563), .CP(CLK), .Q(
        o_data_forward_reg[252]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__1_ ( .D(N562), .CP(CLK), .Q(
        o_data_forward_reg[251]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_4__0_ ( .D(N561), .CP(CLK), .Q(
        o_data_forward_reg[250]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_4_ ( .D(N586), .CP(CLK), .Q(
        o_valid_forward_reg[4]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_5__3_ ( .D(N698), .CP(CLK), .Q(
        o_cmd_forward_reg[39]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_5__2_ ( .D(N697), .CP(CLK), .Q(
        o_cmd_forward_reg[38]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_5__1_ ( .D(N696), .CP(CLK), .Q(
        o_cmd_forward_reg[37]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_5__0_ ( .D(n253), .CP(CLK), .Q(
        o_cmd_forward_reg[36]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__24_ ( .D(N693), .CP(CLK), .Q(
        o_data_forward_reg[249]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__23_ ( .D(N692), .CP(CLK), .Q(
        o_data_forward_reg[248]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__22_ ( .D(N691), .CP(CLK), .Q(
        o_data_forward_reg[247]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__21_ ( .D(N690), .CP(CLK), .Q(
        o_data_forward_reg[246]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__20_ ( .D(N689), .CP(CLK), .Q(
        o_data_forward_reg[245]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__19_ ( .D(N688), .CP(CLK), .Q(
        o_data_forward_reg[244]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__18_ ( .D(N687), .CP(CLK), .Q(
        o_data_forward_reg[243]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__17_ ( .D(N686), .CP(CLK), .Q(
        o_data_forward_reg[242]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__16_ ( .D(N685), .CP(CLK), .Q(
        o_data_forward_reg[241]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__15_ ( .D(N684), .CP(CLK), .Q(
        o_data_forward_reg[240]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__14_ ( .D(N683), .CP(CLK), .Q(
        o_data_forward_reg[239]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__13_ ( .D(N682), .CP(CLK), .Q(
        o_data_forward_reg[238]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__12_ ( .D(N681), .CP(CLK), .Q(
        o_data_forward_reg[237]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__11_ ( .D(N680), .CP(CLK), .Q(
        o_data_forward_reg[236]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__10_ ( .D(N679), .CP(CLK), .Q(
        o_data_forward_reg[235]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__9_ ( .D(N678), .CP(CLK), .Q(
        o_data_forward_reg[234]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__8_ ( .D(N677), .CP(CLK), .Q(
        o_data_forward_reg[233]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__7_ ( .D(N676), .CP(CLK), .Q(
        o_data_forward_reg[232]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__6_ ( .D(N675), .CP(CLK), .Q(
        o_data_forward_reg[231]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__5_ ( .D(N674), .CP(CLK), .Q(
        o_data_forward_reg[230]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__4_ ( .D(N673), .CP(CLK), .Q(
        o_data_forward_reg[229]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__3_ ( .D(N672), .CP(CLK), .Q(
        o_data_forward_reg[228]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__2_ ( .D(N671), .CP(CLK), .Q(
        o_data_forward_reg[227]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__1_ ( .D(N670), .CP(CLK), .Q(
        o_data_forward_reg[226]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_5__0_ ( .D(N669), .CP(CLK), .Q(
        o_data_forward_reg[225]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_5_ ( .D(N694), .CP(CLK), .Q(
        o_valid_forward_reg[5]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_6__3_ ( .D(N806), .CP(CLK), .Q(
        o_cmd_forward_reg[35]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_6__2_ ( .D(N805), .CP(CLK), .Q(
        o_cmd_forward_reg[34]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_6__1_ ( .D(n247), .CP(CLK), .Q(
        o_cmd_forward_reg[33]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_6__0_ ( .D(N803), .CP(CLK), .Q(
        o_cmd_forward_reg[32]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__24_ ( .D(N801), .CP(CLK), .Q(
        o_data_forward_reg[224]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__23_ ( .D(N800), .CP(CLK), .Q(
        o_data_forward_reg[223]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__22_ ( .D(N799), .CP(CLK), .Q(
        o_data_forward_reg[222]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__21_ ( .D(N798), .CP(CLK), .Q(
        o_data_forward_reg[221]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__20_ ( .D(N797), .CP(CLK), .Q(
        o_data_forward_reg[220]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__19_ ( .D(N796), .CP(CLK), .Q(
        o_data_forward_reg[219]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__18_ ( .D(N795), .CP(CLK), .Q(
        o_data_forward_reg[218]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__17_ ( .D(N794), .CP(CLK), .Q(
        o_data_forward_reg[217]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__16_ ( .D(N793), .CP(CLK), .Q(
        o_data_forward_reg[216]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__15_ ( .D(N792), .CP(CLK), .Q(
        o_data_forward_reg[215]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__14_ ( .D(N791), .CP(CLK), .Q(
        o_data_forward_reg[214]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__13_ ( .D(N790), .CP(CLK), .Q(
        o_data_forward_reg[213]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__12_ ( .D(N789), .CP(CLK), .Q(
        o_data_forward_reg[212]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__11_ ( .D(N788), .CP(CLK), .Q(
        o_data_forward_reg[211]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__10_ ( .D(N787), .CP(CLK), .Q(
        o_data_forward_reg[210]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__9_ ( .D(N786), .CP(CLK), .Q(
        o_data_forward_reg[209]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__8_ ( .D(N785), .CP(CLK), .Q(
        o_data_forward_reg[208]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__7_ ( .D(N784), .CP(CLK), .Q(
        o_data_forward_reg[207]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__6_ ( .D(N783), .CP(CLK), .Q(
        o_data_forward_reg[206]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__5_ ( .D(N782), .CP(CLK), .Q(
        o_data_forward_reg[205]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__4_ ( .D(N781), .CP(CLK), .Q(
        o_data_forward_reg[204]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__3_ ( .D(N780), .CP(CLK), .Q(
        o_data_forward_reg[203]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__2_ ( .D(N779), .CP(CLK), .Q(
        o_data_forward_reg[202]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__1_ ( .D(N778), .CP(CLK), .Q(
        o_data_forward_reg[201]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_6__0_ ( .D(N777), .CP(CLK), .Q(
        o_data_forward_reg[200]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_6_ ( .D(N802), .CP(CLK), .Q(
        o_valid_forward_reg[6]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_7__3_ ( .D(N914), .CP(CLK), .Q(
        o_cmd_forward_reg[31]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_7__2_ ( .D(n256), .CP(CLK), .Q(
        o_cmd_forward_reg[30]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_7__1_ ( .D(N912), .CP(CLK), .Q(
        o_cmd_forward_reg[29]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_7__0_ ( .D(N911), .CP(CLK), .Q(
        o_cmd_forward_reg[28]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__24_ ( .D(N909), .CP(CLK), .Q(
        o_data_forward_reg[199]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__23_ ( .D(N908), .CP(CLK), .Q(
        o_data_forward_reg[198]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__22_ ( .D(N907), .CP(CLK), .Q(
        o_data_forward_reg[197]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__21_ ( .D(N906), .CP(CLK), .Q(
        o_data_forward_reg[196]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__20_ ( .D(N905), .CP(CLK), .Q(
        o_data_forward_reg[195]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__19_ ( .D(N904), .CP(CLK), .Q(
        o_data_forward_reg[194]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__18_ ( .D(N903), .CP(CLK), .Q(
        o_data_forward_reg[193]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__17_ ( .D(N902), .CP(CLK), .Q(
        o_data_forward_reg[192]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__16_ ( .D(N901), .CP(CLK), .Q(
        o_data_forward_reg[191]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__15_ ( .D(N900), .CP(CLK), .Q(
        o_data_forward_reg[190]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__14_ ( .D(N899), .CP(CLK), .Q(
        o_data_forward_reg[189]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__13_ ( .D(N898), .CP(CLK), .Q(
        o_data_forward_reg[188]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__12_ ( .D(N897), .CP(CLK), .Q(
        o_data_forward_reg[187]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__11_ ( .D(N896), .CP(CLK), .Q(
        o_data_forward_reg[186]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__10_ ( .D(N895), .CP(CLK), .Q(
        o_data_forward_reg[185]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__9_ ( .D(N894), .CP(CLK), .Q(
        o_data_forward_reg[184]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__8_ ( .D(N893), .CP(CLK), .Q(
        o_data_forward_reg[183]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__7_ ( .D(N892), .CP(CLK), .Q(
        o_data_forward_reg[182]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__6_ ( .D(N891), .CP(CLK), .Q(
        o_data_forward_reg[181]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__5_ ( .D(N890), .CP(CLK), .Q(
        o_data_forward_reg[180]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__4_ ( .D(N889), .CP(CLK), .Q(
        o_data_forward_reg[179]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__3_ ( .D(N888), .CP(CLK), .Q(
        o_data_forward_reg[178]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__2_ ( .D(N887), .CP(CLK), .Q(
        o_data_forward_reg[177]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__1_ ( .D(N886), .CP(CLK), .Q(
        o_data_forward_reg[176]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_7__0_ ( .D(N885), .CP(CLK), .Q(
        o_data_forward_reg[175]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_7_ ( .D(N910), .CP(CLK), .Q(
        o_valid_forward_reg[7]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_8__3_ ( .D(n245), .CP(CLK), .Q(
        o_cmd_forward_reg[27]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_8__2_ ( .D(N1021), .CP(CLK), .Q(
        o_cmd_forward_reg[26]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_8__1_ ( .D(N1020), .CP(CLK), .Q(
        o_cmd_forward_reg[25]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_8__0_ ( .D(N1019), .CP(CLK), .Q(
        o_cmd_forward_reg[24]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__24_ ( .D(N1017), .CP(CLK), .Q(
        o_data_forward_reg[174]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__23_ ( .D(N1016), .CP(CLK), .Q(
        o_data_forward_reg[173]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__22_ ( .D(N1015), .CP(CLK), .Q(
        o_data_forward_reg[172]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__21_ ( .D(N1014), .CP(CLK), .Q(
        o_data_forward_reg[171]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__20_ ( .D(N1013), .CP(CLK), .Q(
        o_data_forward_reg[170]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__19_ ( .D(N1012), .CP(CLK), .Q(
        o_data_forward_reg[169]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__18_ ( .D(N1011), .CP(CLK), .Q(
        o_data_forward_reg[168]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__17_ ( .D(N1010), .CP(CLK), .Q(
        o_data_forward_reg[167]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__16_ ( .D(N1009), .CP(CLK), .Q(
        o_data_forward_reg[166]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__15_ ( .D(N1008), .CP(CLK), .Q(
        o_data_forward_reg[165]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__14_ ( .D(N1007), .CP(CLK), .Q(
        o_data_forward_reg[164]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__13_ ( .D(N1006), .CP(CLK), .Q(
        o_data_forward_reg[163]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__12_ ( .D(N1005), .CP(CLK), .Q(
        o_data_forward_reg[162]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__11_ ( .D(N1004), .CP(CLK), .Q(
        o_data_forward_reg[161]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__10_ ( .D(N1003), .CP(CLK), .Q(
        o_data_forward_reg[160]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__9_ ( .D(N1002), .CP(CLK), .Q(
        o_data_forward_reg[159]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__8_ ( .D(N1001), .CP(CLK), .Q(
        o_data_forward_reg[158]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__7_ ( .D(N1000), .CP(CLK), .Q(
        o_data_forward_reg[157]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__6_ ( .D(N999), .CP(CLK), .Q(
        o_data_forward_reg[156]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__5_ ( .D(N998), .CP(CLK), .Q(
        o_data_forward_reg[155]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__4_ ( .D(N997), .CP(CLK), .Q(
        o_data_forward_reg[154]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__3_ ( .D(N996), .CP(CLK), .Q(
        o_data_forward_reg[153]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__2_ ( .D(N995), .CP(CLK), .Q(
        o_data_forward_reg[152]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__1_ ( .D(N994), .CP(CLK), .Q(
        o_data_forward_reg[151]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_8__0_ ( .D(N993), .CP(CLK), .Q(
        o_data_forward_reg[150]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_8_ ( .D(N1018), .CP(CLK), .Q(
        o_valid_forward_reg[8]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_9__3_ ( .D(N1130), .CP(CLK), .Q(
        o_cmd_forward_reg[23]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_9__2_ ( .D(N1129), .CP(CLK), .Q(
        o_cmd_forward_reg[22]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_9__1_ ( .D(N1128), .CP(CLK), .Q(
        o_cmd_forward_reg[21]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_9__0_ ( .D(n254), .CP(CLK), .Q(
        o_cmd_forward_reg[20]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__24_ ( .D(N1125), .CP(CLK), .Q(
        o_data_forward_reg[149]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__23_ ( .D(N1124), .CP(CLK), .Q(
        o_data_forward_reg[148]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__22_ ( .D(N1123), .CP(CLK), .Q(
        o_data_forward_reg[147]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__21_ ( .D(N1122), .CP(CLK), .Q(
        o_data_forward_reg[146]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__20_ ( .D(N1121), .CP(CLK), .Q(
        o_data_forward_reg[145]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__19_ ( .D(N1120), .CP(CLK), .Q(
        o_data_forward_reg[144]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__18_ ( .D(N1119), .CP(CLK), .Q(
        o_data_forward_reg[143]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__17_ ( .D(N1118), .CP(CLK), .Q(
        o_data_forward_reg[142]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__16_ ( .D(N1117), .CP(CLK), .Q(
        o_data_forward_reg[141]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__15_ ( .D(N1116), .CP(CLK), .Q(
        o_data_forward_reg[140]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__14_ ( .D(N1115), .CP(CLK), .Q(
        o_data_forward_reg[139]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__13_ ( .D(N1114), .CP(CLK), .Q(
        o_data_forward_reg[138]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__12_ ( .D(N1113), .CP(CLK), .Q(
        o_data_forward_reg[137]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__11_ ( .D(N1112), .CP(CLK), .Q(
        o_data_forward_reg[136]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__10_ ( .D(N1111), .CP(CLK), .Q(
        o_data_forward_reg[135]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__9_ ( .D(N1110), .CP(CLK), .Q(
        o_data_forward_reg[134]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__8_ ( .D(N1109), .CP(CLK), .Q(
        o_data_forward_reg[133]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__7_ ( .D(N1108), .CP(CLK), .Q(
        o_data_forward_reg[132]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__6_ ( .D(N1107), .CP(CLK), .Q(
        o_data_forward_reg[131]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__5_ ( .D(N1106), .CP(CLK), .Q(
        o_data_forward_reg[130]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__4_ ( .D(N1105), .CP(CLK), .Q(
        o_data_forward_reg[129]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__3_ ( .D(N1104), .CP(CLK), .Q(
        o_data_forward_reg[128]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__2_ ( .D(N1103), .CP(CLK), .Q(
        o_data_forward_reg[127]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__1_ ( .D(N1102), .CP(CLK), .Q(
        o_data_forward_reg[126]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_9__0_ ( .D(N1101), .CP(CLK), .Q(
        o_data_forward_reg[125]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_9_ ( .D(N1126), .CP(CLK), .Q(
        o_valid_forward_reg[9]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_10__3_ ( .D(n255), .CP(CLK), .Q(
        o_cmd_forward_reg[19]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_10__2_ ( .D(N1237), .CP(CLK), .Q(
        o_cmd_forward_reg[18]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_10__1_ ( .D(N1236), .CP(CLK), .Q(
        o_cmd_forward_reg[17]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_10__0_ ( .D(N1235), .CP(CLK), .Q(
        o_cmd_forward_reg[16]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__24_ ( .D(N1233), .CP(CLK), .Q(
        o_data_forward_reg[124]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__23_ ( .D(N1232), .CP(CLK), .Q(
        o_data_forward_reg[123]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__22_ ( .D(N1231), .CP(CLK), .Q(
        o_data_forward_reg[122]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__21_ ( .D(N1230), .CP(CLK), .Q(
        o_data_forward_reg[121]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__20_ ( .D(N1229), .CP(CLK), .Q(
        o_data_forward_reg[120]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__19_ ( .D(N1228), .CP(CLK), .Q(
        o_data_forward_reg[119]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__18_ ( .D(N1227), .CP(CLK), .Q(
        o_data_forward_reg[118]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__17_ ( .D(N1226), .CP(CLK), .Q(
        o_data_forward_reg[117]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__16_ ( .D(N1225), .CP(CLK), .Q(
        o_data_forward_reg[116]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__15_ ( .D(N1224), .CP(CLK), .Q(
        o_data_forward_reg[115]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__14_ ( .D(N1223), .CP(CLK), .Q(
        o_data_forward_reg[114]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__13_ ( .D(N1222), .CP(CLK), .Q(
        o_data_forward_reg[113]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__12_ ( .D(N1221), .CP(CLK), .Q(
        o_data_forward_reg[112]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__11_ ( .D(N1220), .CP(CLK), .Q(
        o_data_forward_reg[111]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__10_ ( .D(N1219), .CP(CLK), .Q(
        o_data_forward_reg[110]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__9_ ( .D(N1218), .CP(CLK), .Q(
        o_data_forward_reg[109]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__8_ ( .D(N1217), .CP(CLK), .Q(
        o_data_forward_reg[108]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__7_ ( .D(N1216), .CP(CLK), .Q(
        o_data_forward_reg[107]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__6_ ( .D(N1215), .CP(CLK), .Q(
        o_data_forward_reg[106]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__5_ ( .D(N1214), .CP(CLK), .Q(
        o_data_forward_reg[105]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__4_ ( .D(N1213), .CP(CLK), .Q(
        o_data_forward_reg[104]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__3_ ( .D(N1212), .CP(CLK), .Q(
        o_data_forward_reg[103]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__2_ ( .D(N1211), .CP(CLK), .Q(
        o_data_forward_reg[102]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__1_ ( .D(N1210), .CP(CLK), .Q(
        o_data_forward_reg[101]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_10__0_ ( .D(N1209), .CP(CLK), .Q(
        o_data_forward_reg[100]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_10_ ( .D(N1234), .CP(CLK), .Q(
        o_valid_forward_reg[10]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_11__3_ ( .D(N1346), .CP(CLK), .Q(
        o_cmd_forward_reg[15]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_11__2_ ( .D(N1345), .CP(CLK), .Q(
        o_cmd_forward_reg[14]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_11__1_ ( .D(n257), .CP(CLK), .Q(
        o_cmd_forward_reg[13]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_11__0_ ( .D(N1343), .CP(CLK), .Q(
        o_cmd_forward_reg[12]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__24_ ( .D(N1341), .CP(CLK), .Q(
        o_data_forward_reg[99]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__23_ ( .D(N1340), .CP(CLK), .Q(
        o_data_forward_reg[98]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__22_ ( .D(N1339), .CP(CLK), .Q(
        o_data_forward_reg[97]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__21_ ( .D(N1338), .CP(CLK), .Q(
        o_data_forward_reg[96]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__20_ ( .D(N1337), .CP(CLK), .Q(
        o_data_forward_reg[95]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__19_ ( .D(N1336), .CP(CLK), .Q(
        o_data_forward_reg[94]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__18_ ( .D(N1335), .CP(CLK), .Q(
        o_data_forward_reg[93]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__17_ ( .D(N1334), .CP(CLK), .Q(
        o_data_forward_reg[92]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__16_ ( .D(N1333), .CP(CLK), .Q(
        o_data_forward_reg[91]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__15_ ( .D(N1332), .CP(CLK), .Q(
        o_data_forward_reg[90]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__14_ ( .D(N1331), .CP(CLK), .Q(
        o_data_forward_reg[89]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__13_ ( .D(N1330), .CP(CLK), .Q(
        o_data_forward_reg[88]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__12_ ( .D(N1329), .CP(CLK), .Q(
        o_data_forward_reg[87]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__11_ ( .D(N1328), .CP(CLK), .Q(
        o_data_forward_reg[86]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__10_ ( .D(N1327), .CP(CLK), .Q(
        o_data_forward_reg[85]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__9_ ( .D(N1326), .CP(CLK), .Q(
        o_data_forward_reg[84]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__8_ ( .D(N1325), .CP(CLK), .Q(
        o_data_forward_reg[83]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__7_ ( .D(N1324), .CP(CLK), .Q(
        o_data_forward_reg[82]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__6_ ( .D(N1323), .CP(CLK), .Q(
        o_data_forward_reg[81]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__5_ ( .D(N1322), .CP(CLK), .Q(
        o_data_forward_reg[80]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__4_ ( .D(N1321), .CP(CLK), .Q(
        o_data_forward_reg[79]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__3_ ( .D(N1320), .CP(CLK), .Q(
        o_data_forward_reg[78]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__2_ ( .D(N1319), .CP(CLK), .Q(
        o_data_forward_reg[77]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__1_ ( .D(N1318), .CP(CLK), .Q(
        o_data_forward_reg[76]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_11__0_ ( .D(N1317), .CP(CLK), .Q(
        o_data_forward_reg[75]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_11_ ( .D(N1342), .CP(CLK), .Q(
        o_valid_forward_reg[11]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_12__3_ ( .D(n259), .CP(CLK), .Q(
        o_cmd_forward_reg[11]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_12__2_ ( .D(N1453), .CP(CLK), .Q(
        o_cmd_forward_reg[10]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_12__1_ ( .D(N1452), .CP(CLK), .Q(
        o_cmd_forward_reg[9]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_12__0_ ( .D(N1451), .CP(CLK), .Q(
        o_cmd_forward_reg[8]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__24_ ( .D(N1449), .CP(CLK), .Q(
        o_data_forward_reg[74]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__23_ ( .D(N1448), .CP(CLK), .Q(
        o_data_forward_reg[73]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__22_ ( .D(N1447), .CP(CLK), .Q(
        o_data_forward_reg[72]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__21_ ( .D(N1446), .CP(CLK), .Q(
        o_data_forward_reg[71]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__20_ ( .D(N1445), .CP(CLK), .Q(
        o_data_forward_reg[70]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__19_ ( .D(N1444), .CP(CLK), .Q(
        o_data_forward_reg[69]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__18_ ( .D(N1443), .CP(CLK), .Q(
        o_data_forward_reg[68]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__17_ ( .D(N1442), .CP(CLK), .Q(
        o_data_forward_reg[67]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__16_ ( .D(N1441), .CP(CLK), .Q(
        o_data_forward_reg[66]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__15_ ( .D(N1440), .CP(CLK), .Q(
        o_data_forward_reg[65]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__14_ ( .D(N1439), .CP(CLK), .Q(
        o_data_forward_reg[64]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__13_ ( .D(N1438), .CP(CLK), .Q(
        o_data_forward_reg[63]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__12_ ( .D(N1437), .CP(CLK), .Q(
        o_data_forward_reg[62]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__11_ ( .D(N1436), .CP(CLK), .Q(
        o_data_forward_reg[61]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__10_ ( .D(N1435), .CP(CLK), .Q(
        o_data_forward_reg[60]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__9_ ( .D(N1434), .CP(CLK), .Q(
        o_data_forward_reg[59]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__8_ ( .D(N1433), .CP(CLK), .Q(
        o_data_forward_reg[58]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__7_ ( .D(N1432), .CP(CLK), .Q(
        o_data_forward_reg[57]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__6_ ( .D(N1431), .CP(CLK), .Q(
        o_data_forward_reg[56]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__5_ ( .D(N1430), .CP(CLK), .Q(
        o_data_forward_reg[55]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__4_ ( .D(N1429), .CP(CLK), .Q(
        o_data_forward_reg[54]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__3_ ( .D(N1428), .CP(CLK), .Q(
        o_data_forward_reg[53]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__2_ ( .D(N1427), .CP(CLK), .Q(
        o_data_forward_reg[52]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__1_ ( .D(N1426), .CP(CLK), .Q(
        o_data_forward_reg[51]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_12__0_ ( .D(N1425), .CP(CLK), .Q(
        o_data_forward_reg[50]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_12_ ( .D(N1450), .CP(CLK), .Q(
        o_valid_forward_reg[12]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_13__3_ ( .D(n258), .CP(CLK), .Q(
        o_cmd_forward_reg[7]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_13__2_ ( .D(N1561), .CP(CLK), .Q(
        o_cmd_forward_reg[6]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_13__1_ ( .D(N1560), .CP(CLK), .Q(
        o_cmd_forward_reg[5]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_13__0_ ( .D(N1559), .CP(CLK), .Q(
        o_cmd_forward_reg[4]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__24_ ( .D(N1557), .CP(CLK), .Q(
        o_data_forward_reg[49]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__23_ ( .D(N1556), .CP(CLK), .Q(
        o_data_forward_reg[48]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__22_ ( .D(N1555), .CP(CLK), .Q(
        o_data_forward_reg[47]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__21_ ( .D(N1554), .CP(CLK), .Q(
        o_data_forward_reg[46]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__20_ ( .D(N1553), .CP(CLK), .Q(
        o_data_forward_reg[45]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__19_ ( .D(N1552), .CP(CLK), .Q(
        o_data_forward_reg[44]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__18_ ( .D(N1551), .CP(CLK), .Q(
        o_data_forward_reg[43]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__17_ ( .D(N1550), .CP(CLK), .Q(
        o_data_forward_reg[42]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__16_ ( .D(N1549), .CP(CLK), .Q(
        o_data_forward_reg[41]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__15_ ( .D(N1548), .CP(CLK), .Q(
        o_data_forward_reg[40]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__14_ ( .D(N1547), .CP(CLK), .Q(
        o_data_forward_reg[39]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__13_ ( .D(N1546), .CP(CLK), .Q(
        o_data_forward_reg[38]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__12_ ( .D(N1545), .CP(CLK), .Q(
        o_data_forward_reg[37]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__11_ ( .D(N1544), .CP(CLK), .Q(
        o_data_forward_reg[36]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__10_ ( .D(N1543), .CP(CLK), .Q(
        o_data_forward_reg[35]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__9_ ( .D(N1542), .CP(CLK), .Q(
        o_data_forward_reg[34]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__8_ ( .D(N1541), .CP(CLK), .Q(
        o_data_forward_reg[33]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__7_ ( .D(N1540), .CP(CLK), .Q(
        o_data_forward_reg[32]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__6_ ( .D(N1539), .CP(CLK), .Q(
        o_data_forward_reg[31]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__5_ ( .D(N1538), .CP(CLK), .Q(
        o_data_forward_reg[30]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__4_ ( .D(N1537), .CP(CLK), .Q(
        o_data_forward_reg[29]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__3_ ( .D(N1536), .CP(CLK), .Q(
        o_data_forward_reg[28]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__2_ ( .D(N1535), .CP(CLK), .Q(
        o_data_forward_reg[27]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__1_ ( .D(N1534), .CP(CLK), .Q(
        o_data_forward_reg[26]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_13__0_ ( .D(N1533), .CP(CLK), .Q(
        o_data_forward_reg[25]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_13_ ( .D(N1558), .CP(CLK), .Q(
        o_valid_forward_reg[13]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_14__3_ ( .D(N1670), .CP(CLK), .Q(
        o_cmd_forward_reg[3]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_14__2_ ( .D(n244), .CP(CLK), .Q(
        o_cmd_forward_reg[2]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_14__1_ ( .D(N1668), .CP(CLK), .Q(
        o_cmd_forward_reg[1]) );
  DFQD1BWP30P140LVT o_cmd_forward_reg_reg_14__0_ ( .D(N1667), .CP(CLK), .Q(
        o_cmd_forward_reg[0]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__24_ ( .D(N1665), .CP(CLK), .Q(
        o_data_forward_reg[24]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__23_ ( .D(N1664), .CP(CLK), .Q(
        o_data_forward_reg[23]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__22_ ( .D(N1663), .CP(CLK), .Q(
        o_data_forward_reg[22]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__21_ ( .D(N1662), .CP(CLK), .Q(
        o_data_forward_reg[21]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__20_ ( .D(N1661), .CP(CLK), .Q(
        o_data_forward_reg[20]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__19_ ( .D(N1660), .CP(CLK), .Q(
        o_data_forward_reg[19]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__18_ ( .D(N1659), .CP(CLK), .Q(
        o_data_forward_reg[18]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__17_ ( .D(N1658), .CP(CLK), .Q(
        o_data_forward_reg[17]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__16_ ( .D(N1657), .CP(CLK), .Q(
        o_data_forward_reg[16]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__15_ ( .D(N1656), .CP(CLK), .Q(
        o_data_forward_reg[15]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__14_ ( .D(N1655), .CP(CLK), .Q(
        o_data_forward_reg[14]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__13_ ( .D(N1654), .CP(CLK), .Q(
        o_data_forward_reg[13]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__12_ ( .D(N1653), .CP(CLK), .Q(
        o_data_forward_reg[12]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__11_ ( .D(N1652), .CP(CLK), .Q(
        o_data_forward_reg[11]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__10_ ( .D(N1651), .CP(CLK), .Q(
        o_data_forward_reg[10]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__9_ ( .D(N1650), .CP(CLK), .Q(
        o_data_forward_reg[9]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__8_ ( .D(N1649), .CP(CLK), .Q(
        o_data_forward_reg[8]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__7_ ( .D(N1648), .CP(CLK), .Q(
        o_data_forward_reg[7]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__6_ ( .D(N1647), .CP(CLK), .Q(
        o_data_forward_reg[6]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__5_ ( .D(N1646), .CP(CLK), .Q(
        o_data_forward_reg[5]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__4_ ( .D(N1645), .CP(CLK), .Q(
        o_data_forward_reg[4]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__3_ ( .D(N1644), .CP(CLK), .Q(
        o_data_forward_reg[3]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__2_ ( .D(N1643), .CP(CLK), .Q(
        o_data_forward_reg[2]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__1_ ( .D(N1642), .CP(CLK), .Q(
        o_data_forward_reg[1]) );
  DFQD1BWP30P140LVT o_data_forward_reg_reg_14__0_ ( .D(N1641), .CP(CLK), .Q(
        o_data_forward_reg[0]) );
  DFQD1BWP30P140LVT o_valid_forward_reg_reg_14_ ( .D(N1666), .CP(CLK), .Q(
        o_valid_forward_reg[14]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_15_ ( .D(n234), .CP(CLK), .Q(o_valid[15])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_14_ ( .D(n243), .CP(CLK), .Q(o_valid[14])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_13_ ( .D(n242), .CP(CLK), .Q(o_valid[13])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_12_ ( .D(n233), .CP(CLK), .Q(o_valid[12])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_11_ ( .D(n241), .CP(CLK), .Q(o_valid[11])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_10_ ( .D(n232), .CP(CLK), .Q(o_valid[10])
         );
  DFQD4BWP30P140LVT o_valid_reg_reg_9_ ( .D(n240), .CP(CLK), .Q(o_valid[9]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_8_ ( .D(n19), .CP(CLK), .Q(o_valid[8]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_7_ ( .D(n246), .CP(CLK), .Q(o_valid[7]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_6_ ( .D(n231), .CP(CLK), .Q(o_valid[6]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_5_ ( .D(n238), .CP(CLK), .Q(o_valid[5]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_4_ ( .D(n21), .CP(CLK), .Q(o_valid[4]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_3_ ( .D(n230), .CP(CLK), .Q(o_valid[3]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_2_ ( .D(n20), .CP(CLK), .Q(o_valid[2]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_1_ ( .D(n22), .CP(CLK), .Q(o_valid[1]) );
  DFQD4BWP30P140LVT o_valid_reg_reg_0_ ( .D(n229), .CP(CLK), .Q(o_valid[0]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_399_ ( .D(n113), .CP(CLK), .Q(
        o_data_bus[399]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_398_ ( .D(n112), .CP(CLK), .Q(
        o_data_bus[398]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_397_ ( .D(n111), .CP(CLK), .Q(
        o_data_bus[397]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_396_ ( .D(n110), .CP(CLK), .Q(
        o_data_bus[396]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_395_ ( .D(n109), .CP(CLK), .Q(
        o_data_bus[395]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_394_ ( .D(n108), .CP(CLK), .Q(
        o_data_bus[394]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_393_ ( .D(n107), .CP(CLK), .Q(
        o_data_bus[393]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_392_ ( .D(n106), .CP(CLK), .Q(
        o_data_bus[392]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_391_ ( .D(n105), .CP(CLK), .Q(
        o_data_bus[391]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_390_ ( .D(n104), .CP(CLK), .Q(
        o_data_bus[390]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_389_ ( .D(n103), .CP(CLK), .Q(
        o_data_bus[389]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_388_ ( .D(n102), .CP(CLK), .Q(
        o_data_bus[388]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_387_ ( .D(n215), .CP(CLK), .Q(
        o_data_bus[387]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_386_ ( .D(n214), .CP(CLK), .Q(
        o_data_bus[386]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_385_ ( .D(n213), .CP(CLK), .Q(
        o_data_bus[385]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_384_ ( .D(n212), .CP(CLK), .Q(
        o_data_bus[384]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_383_ ( .D(n211), .CP(CLK), .Q(
        o_data_bus[383]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_382_ ( .D(n210), .CP(CLK), .Q(
        o_data_bus[382]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_381_ ( .D(n209), .CP(CLK), .Q(
        o_data_bus[381]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_380_ ( .D(n208), .CP(CLK), .Q(
        o_data_bus[380]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_379_ ( .D(n207), .CP(CLK), .Q(
        o_data_bus[379]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_378_ ( .D(n206), .CP(CLK), .Q(
        o_data_bus[378]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_377_ ( .D(n205), .CP(CLK), .Q(
        o_data_bus[377]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_376_ ( .D(n204), .CP(CLK), .Q(
        o_data_bus[376]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_375_ ( .D(n203), .CP(CLK), .Q(
        o_data_bus[375]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_374_ ( .D(N1640), .CP(CLK), .Q(
        o_data_bus[374]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_373_ ( .D(N1639), .CP(CLK), .Q(
        o_data_bus[373]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_372_ ( .D(N1638), .CP(CLK), .Q(
        o_data_bus[372]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_371_ ( .D(N1637), .CP(CLK), .Q(
        o_data_bus[371]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_370_ ( .D(N1636), .CP(CLK), .Q(
        o_data_bus[370]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_369_ ( .D(N1635), .CP(CLK), .Q(
        o_data_bus[369]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_368_ ( .D(N1634), .CP(CLK), .Q(
        o_data_bus[368]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_367_ ( .D(N1633), .CP(CLK), .Q(
        o_data_bus[367]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_366_ ( .D(N1632), .CP(CLK), .Q(
        o_data_bus[366]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_365_ ( .D(N1631), .CP(CLK), .Q(
        o_data_bus[365]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_364_ ( .D(N1630), .CP(CLK), .Q(
        o_data_bus[364]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_363_ ( .D(N1629), .CP(CLK), .Q(
        o_data_bus[363]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_362_ ( .D(N1628), .CP(CLK), .Q(
        o_data_bus[362]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_361_ ( .D(N1627), .CP(CLK), .Q(
        o_data_bus[361]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_360_ ( .D(N1626), .CP(CLK), .Q(
        o_data_bus[360]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_359_ ( .D(N1625), .CP(CLK), .Q(
        o_data_bus[359]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_358_ ( .D(N1624), .CP(CLK), .Q(
        o_data_bus[358]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_357_ ( .D(N1623), .CP(CLK), .Q(
        o_data_bus[357]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_356_ ( .D(N1622), .CP(CLK), .Q(
        o_data_bus[356]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_355_ ( .D(N1621), .CP(CLK), .Q(
        o_data_bus[355]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_354_ ( .D(N1620), .CP(CLK), .Q(
        o_data_bus[354]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_353_ ( .D(N1619), .CP(CLK), .Q(
        o_data_bus[353]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_352_ ( .D(N1618), .CP(CLK), .Q(
        o_data_bus[352]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_351_ ( .D(N1617), .CP(CLK), .Q(
        o_data_bus[351]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_350_ ( .D(N1616), .CP(CLK), .Q(
        o_data_bus[350]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_349_ ( .D(N1532), .CP(CLK), .Q(
        o_data_bus[349]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_348_ ( .D(N1531), .CP(CLK), .Q(
        o_data_bus[348]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_347_ ( .D(N1530), .CP(CLK), .Q(
        o_data_bus[347]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_346_ ( .D(N1529), .CP(CLK), .Q(
        o_data_bus[346]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_345_ ( .D(N1528), .CP(CLK), .Q(
        o_data_bus[345]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_344_ ( .D(N1527), .CP(CLK), .Q(
        o_data_bus[344]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_343_ ( .D(N1526), .CP(CLK), .Q(
        o_data_bus[343]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_342_ ( .D(N1525), .CP(CLK), .Q(
        o_data_bus[342]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_341_ ( .D(N1524), .CP(CLK), .Q(
        o_data_bus[341]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_340_ ( .D(N1523), .CP(CLK), .Q(
        o_data_bus[340]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_339_ ( .D(N1522), .CP(CLK), .Q(
        o_data_bus[339]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_338_ ( .D(N1521), .CP(CLK), .Q(
        o_data_bus[338]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_337_ ( .D(N1520), .CP(CLK), .Q(
        o_data_bus[337]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_336_ ( .D(N1519), .CP(CLK), .Q(
        o_data_bus[336]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_335_ ( .D(N1518), .CP(CLK), .Q(
        o_data_bus[335]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_334_ ( .D(N1517), .CP(CLK), .Q(
        o_data_bus[334]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_333_ ( .D(N1516), .CP(CLK), .Q(
        o_data_bus[333]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_332_ ( .D(N1515), .CP(CLK), .Q(
        o_data_bus[332]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_331_ ( .D(N1514), .CP(CLK), .Q(
        o_data_bus[331]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_330_ ( .D(N1513), .CP(CLK), .Q(
        o_data_bus[330]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_329_ ( .D(N1512), .CP(CLK), .Q(
        o_data_bus[329]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_328_ ( .D(N1511), .CP(CLK), .Q(
        o_data_bus[328]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_327_ ( .D(N1510), .CP(CLK), .Q(
        o_data_bus[327]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_326_ ( .D(N1509), .CP(CLK), .Q(
        o_data_bus[326]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_325_ ( .D(N1508), .CP(CLK), .Q(
        o_data_bus[325]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_324_ ( .D(n101), .CP(CLK), .Q(
        o_data_bus[324]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_323_ ( .D(n100), .CP(CLK), .Q(
        o_data_bus[323]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_322_ ( .D(n99), .CP(CLK), .Q(
        o_data_bus[322]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_321_ ( .D(n98), .CP(CLK), .Q(
        o_data_bus[321]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_320_ ( .D(n97), .CP(CLK), .Q(
        o_data_bus[320]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_319_ ( .D(n96), .CP(CLK), .Q(
        o_data_bus[319]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_318_ ( .D(n95), .CP(CLK), .Q(
        o_data_bus[318]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_317_ ( .D(n94), .CP(CLK), .Q(
        o_data_bus[317]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_316_ ( .D(n93), .CP(CLK), .Q(
        o_data_bus[316]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_315_ ( .D(n92), .CP(CLK), .Q(
        o_data_bus[315]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_314_ ( .D(n91), .CP(CLK), .Q(
        o_data_bus[314]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_313_ ( .D(n90), .CP(CLK), .Q(
        o_data_bus[313]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_312_ ( .D(n165), .CP(CLK), .Q(
        o_data_bus[312]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_311_ ( .D(n164), .CP(CLK), .Q(
        o_data_bus[311]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_310_ ( .D(n163), .CP(CLK), .Q(
        o_data_bus[310]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_309_ ( .D(n162), .CP(CLK), .Q(
        o_data_bus[309]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_308_ ( .D(n161), .CP(CLK), .Q(
        o_data_bus[308]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_307_ ( .D(n160), .CP(CLK), .Q(
        o_data_bus[307]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_306_ ( .D(n159), .CP(CLK), .Q(
        o_data_bus[306]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_305_ ( .D(n158), .CP(CLK), .Q(
        o_data_bus[305]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_304_ ( .D(n157), .CP(CLK), .Q(
        o_data_bus[304]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_303_ ( .D(n156), .CP(CLK), .Q(
        o_data_bus[303]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_302_ ( .D(n155), .CP(CLK), .Q(
        o_data_bus[302]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_301_ ( .D(n154), .CP(CLK), .Q(
        o_data_bus[301]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_300_ ( .D(n153), .CP(CLK), .Q(
        o_data_bus[300]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_299_ ( .D(N1316), .CP(CLK), .Q(
        o_data_bus[299]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_298_ ( .D(N1315), .CP(CLK), .Q(
        o_data_bus[298]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_297_ ( .D(N1314), .CP(CLK), .Q(
        o_data_bus[297]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_296_ ( .D(N1313), .CP(CLK), .Q(
        o_data_bus[296]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_295_ ( .D(N1312), .CP(CLK), .Q(
        o_data_bus[295]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_294_ ( .D(N1311), .CP(CLK), .Q(
        o_data_bus[294]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_293_ ( .D(N1310), .CP(CLK), .Q(
        o_data_bus[293]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_292_ ( .D(N1309), .CP(CLK), .Q(
        o_data_bus[292]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_291_ ( .D(N1308), .CP(CLK), .Q(
        o_data_bus[291]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_290_ ( .D(N1307), .CP(CLK), .Q(
        o_data_bus[290]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_289_ ( .D(N1306), .CP(CLK), .Q(
        o_data_bus[289]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_288_ ( .D(N1305), .CP(CLK), .Q(
        o_data_bus[288]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_287_ ( .D(N1304), .CP(CLK), .Q(
        o_data_bus[287]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_286_ ( .D(N1303), .CP(CLK), .Q(
        o_data_bus[286]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_285_ ( .D(N1302), .CP(CLK), .Q(
        o_data_bus[285]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_284_ ( .D(N1301), .CP(CLK), .Q(
        o_data_bus[284]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_283_ ( .D(N1300), .CP(CLK), .Q(
        o_data_bus[283]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_282_ ( .D(N1299), .CP(CLK), .Q(
        o_data_bus[282]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_281_ ( .D(N1298), .CP(CLK), .Q(
        o_data_bus[281]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_280_ ( .D(N1297), .CP(CLK), .Q(
        o_data_bus[280]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_279_ ( .D(N1296), .CP(CLK), .Q(
        o_data_bus[279]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_278_ ( .D(N1295), .CP(CLK), .Q(
        o_data_bus[278]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_277_ ( .D(N1294), .CP(CLK), .Q(
        o_data_bus[277]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_276_ ( .D(N1293), .CP(CLK), .Q(
        o_data_bus[276]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_275_ ( .D(N1292), .CP(CLK), .Q(
        o_data_bus[275]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_274_ ( .D(n89), .CP(CLK), .Q(
        o_data_bus[274]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_273_ ( .D(n88), .CP(CLK), .Q(
        o_data_bus[273]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_272_ ( .D(n87), .CP(CLK), .Q(
        o_data_bus[272]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_271_ ( .D(n86), .CP(CLK), .Q(
        o_data_bus[271]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_270_ ( .D(n85), .CP(CLK), .Q(
        o_data_bus[270]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_269_ ( .D(n84), .CP(CLK), .Q(
        o_data_bus[269]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_268_ ( .D(n83), .CP(CLK), .Q(
        o_data_bus[268]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_267_ ( .D(n82), .CP(CLK), .Q(
        o_data_bus[267]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_266_ ( .D(n81), .CP(CLK), .Q(
        o_data_bus[266]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_265_ ( .D(n80), .CP(CLK), .Q(
        o_data_bus[265]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_264_ ( .D(n79), .CP(CLK), .Q(
        o_data_bus[264]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_263_ ( .D(n78), .CP(CLK), .Q(
        o_data_bus[263]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_262_ ( .D(n152), .CP(CLK), .Q(
        o_data_bus[262]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_261_ ( .D(n151), .CP(CLK), .Q(
        o_data_bus[261]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_260_ ( .D(n150), .CP(CLK), .Q(
        o_data_bus[260]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_259_ ( .D(n149), .CP(CLK), .Q(
        o_data_bus[259]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_258_ ( .D(n148), .CP(CLK), .Q(
        o_data_bus[258]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_257_ ( .D(n147), .CP(CLK), .Q(
        o_data_bus[257]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_256_ ( .D(n146), .CP(CLK), .Q(
        o_data_bus[256]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_255_ ( .D(n145), .CP(CLK), .Q(
        o_data_bus[255]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_254_ ( .D(n144), .CP(CLK), .Q(
        o_data_bus[254]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_253_ ( .D(n143), .CP(CLK), .Q(
        o_data_bus[253]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_252_ ( .D(n142), .CP(CLK), .Q(
        o_data_bus[252]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_251_ ( .D(n141), .CP(CLK), .Q(
        o_data_bus[251]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_250_ ( .D(n140), .CP(CLK), .Q(
        o_data_bus[250]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_249_ ( .D(N1100), .CP(CLK), .Q(
        o_data_bus[249]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_248_ ( .D(N1099), .CP(CLK), .Q(
        o_data_bus[248]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_247_ ( .D(N1098), .CP(CLK), .Q(
        o_data_bus[247]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_246_ ( .D(N1097), .CP(CLK), .Q(
        o_data_bus[246]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_245_ ( .D(N1096), .CP(CLK), .Q(
        o_data_bus[245]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_244_ ( .D(N1095), .CP(CLK), .Q(
        o_data_bus[244]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_243_ ( .D(N1094), .CP(CLK), .Q(
        o_data_bus[243]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_242_ ( .D(N1093), .CP(CLK), .Q(
        o_data_bus[242]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_241_ ( .D(N1092), .CP(CLK), .Q(
        o_data_bus[241]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_240_ ( .D(N1091), .CP(CLK), .Q(
        o_data_bus[240]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_239_ ( .D(N1090), .CP(CLK), .Q(
        o_data_bus[239]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_238_ ( .D(N1089), .CP(CLK), .Q(
        o_data_bus[238]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_237_ ( .D(N1088), .CP(CLK), .Q(
        o_data_bus[237]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_236_ ( .D(N1087), .CP(CLK), .Q(
        o_data_bus[236]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_235_ ( .D(N1086), .CP(CLK), .Q(
        o_data_bus[235]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_234_ ( .D(N1085), .CP(CLK), .Q(
        o_data_bus[234]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_233_ ( .D(N1084), .CP(CLK), .Q(
        o_data_bus[233]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_232_ ( .D(N1083), .CP(CLK), .Q(
        o_data_bus[232]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_231_ ( .D(N1082), .CP(CLK), .Q(
        o_data_bus[231]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_230_ ( .D(N1081), .CP(CLK), .Q(
        o_data_bus[230]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_229_ ( .D(N1080), .CP(CLK), .Q(
        o_data_bus[229]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_228_ ( .D(N1079), .CP(CLK), .Q(
        o_data_bus[228]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_227_ ( .D(N1078), .CP(CLK), .Q(
        o_data_bus[227]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_226_ ( .D(N1077), .CP(CLK), .Q(
        o_data_bus[226]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_225_ ( .D(N1076), .CP(CLK), .Q(
        o_data_bus[225]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_224_ ( .D(N992), .CP(CLK), .Q(
        o_data_bus[224]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_223_ ( .D(N991), .CP(CLK), .Q(
        o_data_bus[223]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_222_ ( .D(N990), .CP(CLK), .Q(
        o_data_bus[222]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_221_ ( .D(N989), .CP(CLK), .Q(
        o_data_bus[221]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_220_ ( .D(N988), .CP(CLK), .Q(
        o_data_bus[220]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_219_ ( .D(N987), .CP(CLK), .Q(
        o_data_bus[219]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_218_ ( .D(N986), .CP(CLK), .Q(
        o_data_bus[218]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_217_ ( .D(N985), .CP(CLK), .Q(
        o_data_bus[217]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_216_ ( .D(N984), .CP(CLK), .Q(
        o_data_bus[216]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_215_ ( .D(N983), .CP(CLK), .Q(
        o_data_bus[215]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_214_ ( .D(N982), .CP(CLK), .Q(
        o_data_bus[214]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_213_ ( .D(N981), .CP(CLK), .Q(
        o_data_bus[213]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_212_ ( .D(N980), .CP(CLK), .Q(
        o_data_bus[212]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_211_ ( .D(N979), .CP(CLK), .Q(
        o_data_bus[211]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_210_ ( .D(N978), .CP(CLK), .Q(
        o_data_bus[210]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_209_ ( .D(N977), .CP(CLK), .Q(
        o_data_bus[209]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_208_ ( .D(N976), .CP(CLK), .Q(
        o_data_bus[208]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_207_ ( .D(N975), .CP(CLK), .Q(
        o_data_bus[207]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_206_ ( .D(N974), .CP(CLK), .Q(
        o_data_bus[206]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_205_ ( .D(N973), .CP(CLK), .Q(
        o_data_bus[205]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_204_ ( .D(N972), .CP(CLK), .Q(
        o_data_bus[204]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_203_ ( .D(N971), .CP(CLK), .Q(
        o_data_bus[203]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_202_ ( .D(N970), .CP(CLK), .Q(
        o_data_bus[202]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_201_ ( .D(N969), .CP(CLK), .Q(
        o_data_bus[201]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_200_ ( .D(N968), .CP(CLK), .Q(
        o_data_bus[200]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_199_ ( .D(N884), .CP(CLK), .Q(
        o_data_bus[199]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_198_ ( .D(N883), .CP(CLK), .Q(
        o_data_bus[198]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_197_ ( .D(N882), .CP(CLK), .Q(
        o_data_bus[197]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_196_ ( .D(N881), .CP(CLK), .Q(
        o_data_bus[196]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_195_ ( .D(N880), .CP(CLK), .Q(
        o_data_bus[195]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_194_ ( .D(N879), .CP(CLK), .Q(
        o_data_bus[194]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_193_ ( .D(N878), .CP(CLK), .Q(
        o_data_bus[193]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_192_ ( .D(N877), .CP(CLK), .Q(
        o_data_bus[192]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_191_ ( .D(N876), .CP(CLK), .Q(
        o_data_bus[191]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_190_ ( .D(N875), .CP(CLK), .Q(
        o_data_bus[190]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_189_ ( .D(N874), .CP(CLK), .Q(
        o_data_bus[189]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_188_ ( .D(N873), .CP(CLK), .Q(
        o_data_bus[188]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_187_ ( .D(N872), .CP(CLK), .Q(
        o_data_bus[187]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_186_ ( .D(N871), .CP(CLK), .Q(
        o_data_bus[186]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_185_ ( .D(N870), .CP(CLK), .Q(
        o_data_bus[185]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_184_ ( .D(N869), .CP(CLK), .Q(
        o_data_bus[184]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_183_ ( .D(N868), .CP(CLK), .Q(
        o_data_bus[183]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_182_ ( .D(N867), .CP(CLK), .Q(
        o_data_bus[182]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_181_ ( .D(N866), .CP(CLK), .Q(
        o_data_bus[181]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_180_ ( .D(N865), .CP(CLK), .Q(
        o_data_bus[180]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_179_ ( .D(N864), .CP(CLK), .Q(
        o_data_bus[179]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_178_ ( .D(N863), .CP(CLK), .Q(
        o_data_bus[178]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_177_ ( .D(N862), .CP(CLK), .Q(
        o_data_bus[177]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_176_ ( .D(N861), .CP(CLK), .Q(
        o_data_bus[176]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_175_ ( .D(N860), .CP(CLK), .Q(
        o_data_bus[175]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_174_ ( .D(n77), .CP(CLK), .Q(
        o_data_bus[174]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_173_ ( .D(n76), .CP(CLK), .Q(
        o_data_bus[173]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_172_ ( .D(n75), .CP(CLK), .Q(
        o_data_bus[172]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_171_ ( .D(n74), .CP(CLK), .Q(
        o_data_bus[171]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_170_ ( .D(n73), .CP(CLK), .Q(
        o_data_bus[170]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_169_ ( .D(n72), .CP(CLK), .Q(
        o_data_bus[169]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_168_ ( .D(n71), .CP(CLK), .Q(
        o_data_bus[168]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_167_ ( .D(n70), .CP(CLK), .Q(
        o_data_bus[167]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_166_ ( .D(n69), .CP(CLK), .Q(
        o_data_bus[166]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_165_ ( .D(n68), .CP(CLK), .Q(
        o_data_bus[165]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_164_ ( .D(n67), .CP(CLK), .Q(
        o_data_bus[164]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_163_ ( .D(n66), .CP(CLK), .Q(
        o_data_bus[163]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_162_ ( .D(n139), .CP(CLK), .Q(
        o_data_bus[162]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_161_ ( .D(n138), .CP(CLK), .Q(
        o_data_bus[161]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_160_ ( .D(n137), .CP(CLK), .Q(
        o_data_bus[160]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_159_ ( .D(n136), .CP(CLK), .Q(
        o_data_bus[159]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_158_ ( .D(n135), .CP(CLK), .Q(
        o_data_bus[158]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_157_ ( .D(n134), .CP(CLK), .Q(
        o_data_bus[157]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_156_ ( .D(n133), .CP(CLK), .Q(
        o_data_bus[156]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_155_ ( .D(n132), .CP(CLK), .Q(
        o_data_bus[155]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_154_ ( .D(n131), .CP(CLK), .Q(
        o_data_bus[154]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_153_ ( .D(n130), .CP(CLK), .Q(
        o_data_bus[153]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_152_ ( .D(n129), .CP(CLK), .Q(
        o_data_bus[152]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_151_ ( .D(n128), .CP(CLK), .Q(
        o_data_bus[151]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_150_ ( .D(n127), .CP(CLK), .Q(
        o_data_bus[150]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_149_ ( .D(N668), .CP(CLK), .Q(
        o_data_bus[149]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_148_ ( .D(N667), .CP(CLK), .Q(
        o_data_bus[148]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_147_ ( .D(N666), .CP(CLK), .Q(
        o_data_bus[147]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_146_ ( .D(N665), .CP(CLK), .Q(
        o_data_bus[146]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_145_ ( .D(N664), .CP(CLK), .Q(
        o_data_bus[145]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_144_ ( .D(N663), .CP(CLK), .Q(
        o_data_bus[144]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_143_ ( .D(N662), .CP(CLK), .Q(
        o_data_bus[143]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_142_ ( .D(N661), .CP(CLK), .Q(
        o_data_bus[142]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_141_ ( .D(N660), .CP(CLK), .Q(
        o_data_bus[141]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_140_ ( .D(N659), .CP(CLK), .Q(
        o_data_bus[140]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_139_ ( .D(N658), .CP(CLK), .Q(
        o_data_bus[139]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_138_ ( .D(N657), .CP(CLK), .Q(
        o_data_bus[138]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_137_ ( .D(N656), .CP(CLK), .Q(
        o_data_bus[137]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_136_ ( .D(N655), .CP(CLK), .Q(
        o_data_bus[136]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_135_ ( .D(N654), .CP(CLK), .Q(
        o_data_bus[135]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_134_ ( .D(N653), .CP(CLK), .Q(
        o_data_bus[134]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_133_ ( .D(N652), .CP(CLK), .Q(
        o_data_bus[133]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_132_ ( .D(N651), .CP(CLK), .Q(
        o_data_bus[132]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_131_ ( .D(N650), .CP(CLK), .Q(
        o_data_bus[131]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_130_ ( .D(N649), .CP(CLK), .Q(
        o_data_bus[130]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_129_ ( .D(N648), .CP(CLK), .Q(
        o_data_bus[129]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_128_ ( .D(N647), .CP(CLK), .Q(
        o_data_bus[128]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_127_ ( .D(N646), .CP(CLK), .Q(
        o_data_bus[127]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_126_ ( .D(N645), .CP(CLK), .Q(
        o_data_bus[126]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_125_ ( .D(N644), .CP(CLK), .Q(
        o_data_bus[125]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_124_ ( .D(N560), .CP(CLK), .Q(
        o_data_bus[124]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_123_ ( .D(N559), .CP(CLK), .Q(
        o_data_bus[123]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_122_ ( .D(N558), .CP(CLK), .Q(
        o_data_bus[122]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_121_ ( .D(N557), .CP(CLK), .Q(
        o_data_bus[121]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_120_ ( .D(N556), .CP(CLK), .Q(
        o_data_bus[120]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_119_ ( .D(N555), .CP(CLK), .Q(
        o_data_bus[119]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_118_ ( .D(N554), .CP(CLK), .Q(
        o_data_bus[118]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_117_ ( .D(N553), .CP(CLK), .Q(
        o_data_bus[117]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_116_ ( .D(N552), .CP(CLK), .Q(
        o_data_bus[116]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_115_ ( .D(N551), .CP(CLK), .Q(
        o_data_bus[115]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_114_ ( .D(N550), .CP(CLK), .Q(
        o_data_bus[114]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_113_ ( .D(N549), .CP(CLK), .Q(
        o_data_bus[113]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_112_ ( .D(N548), .CP(CLK), .Q(
        o_data_bus[112]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_111_ ( .D(N547), .CP(CLK), .Q(
        o_data_bus[111]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_110_ ( .D(N546), .CP(CLK), .Q(
        o_data_bus[110]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_109_ ( .D(N545), .CP(CLK), .Q(
        o_data_bus[109]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_108_ ( .D(N544), .CP(CLK), .Q(
        o_data_bus[108]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_107_ ( .D(N543), .CP(CLK), .Q(
        o_data_bus[107]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_106_ ( .D(N542), .CP(CLK), .Q(
        o_data_bus[106]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_105_ ( .D(N541), .CP(CLK), .Q(
        o_data_bus[105]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_104_ ( .D(N540), .CP(CLK), .Q(
        o_data_bus[104]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_103_ ( .D(N539), .CP(CLK), .Q(
        o_data_bus[103]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_102_ ( .D(N538), .CP(CLK), .Q(
        o_data_bus[102]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_101_ ( .D(N537), .CP(CLK), .Q(
        o_data_bus[101]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_100_ ( .D(N536), .CP(CLK), .Q(
        o_data_bus[100]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_99_ ( .D(n65), .CP(CLK), .Q(
        o_data_bus[99]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_98_ ( .D(n64), .CP(CLK), .Q(
        o_data_bus[98]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_97_ ( .D(n63), .CP(CLK), .Q(
        o_data_bus[97]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_96_ ( .D(n62), .CP(CLK), .Q(
        o_data_bus[96]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_95_ ( .D(n61), .CP(CLK), .Q(
        o_data_bus[95]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_94_ ( .D(n60), .CP(CLK), .Q(
        o_data_bus[94]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_93_ ( .D(n59), .CP(CLK), .Q(
        o_data_bus[93]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_92_ ( .D(n58), .CP(CLK), .Q(
        o_data_bus[92]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_91_ ( .D(n57), .CP(CLK), .Q(
        o_data_bus[91]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_90_ ( .D(n56), .CP(CLK), .Q(
        o_data_bus[90]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_89_ ( .D(n55), .CP(CLK), .Q(
        o_data_bus[89]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_88_ ( .D(n54), .CP(CLK), .Q(
        o_data_bus[88]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_87_ ( .D(n126), .CP(CLK), .Q(
        o_data_bus[87]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_86_ ( .D(n125), .CP(CLK), .Q(
        o_data_bus[86]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_85_ ( .D(n124), .CP(CLK), .Q(
        o_data_bus[85]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_84_ ( .D(n123), .CP(CLK), .Q(
        o_data_bus[84]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_83_ ( .D(n122), .CP(CLK), .Q(
        o_data_bus[83]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_82_ ( .D(n121), .CP(CLK), .Q(
        o_data_bus[82]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_81_ ( .D(n120), .CP(CLK), .Q(
        o_data_bus[81]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_80_ ( .D(n119), .CP(CLK), .Q(
        o_data_bus[80]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_79_ ( .D(n118), .CP(CLK), .Q(
        o_data_bus[79]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_78_ ( .D(n117), .CP(CLK), .Q(
        o_data_bus[78]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_77_ ( .D(n116), .CP(CLK), .Q(
        o_data_bus[77]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_76_ ( .D(n115), .CP(CLK), .Q(
        o_data_bus[76]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_75_ ( .D(n114), .CP(CLK), .Q(
        o_data_bus[75]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_74_ ( .D(N344), .CP(CLK), .Q(
        o_data_bus[74]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_73_ ( .D(N343), .CP(CLK), .Q(
        o_data_bus[73]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_72_ ( .D(N342), .CP(CLK), .Q(
        o_data_bus[72]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_71_ ( .D(N341), .CP(CLK), .Q(
        o_data_bus[71]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_70_ ( .D(N340), .CP(CLK), .Q(
        o_data_bus[70]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_69_ ( .D(N339), .CP(CLK), .Q(
        o_data_bus[69]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_68_ ( .D(N338), .CP(CLK), .Q(
        o_data_bus[68]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_67_ ( .D(N337), .CP(CLK), .Q(
        o_data_bus[67]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_66_ ( .D(N336), .CP(CLK), .Q(
        o_data_bus[66]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_65_ ( .D(N335), .CP(CLK), .Q(
        o_data_bus[65]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_64_ ( .D(N334), .CP(CLK), .Q(
        o_data_bus[64]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_63_ ( .D(N333), .CP(CLK), .Q(
        o_data_bus[63]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_62_ ( .D(N332), .CP(CLK), .Q(
        o_data_bus[62]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_61_ ( .D(N331), .CP(CLK), .Q(
        o_data_bus[61]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_60_ ( .D(N330), .CP(CLK), .Q(
        o_data_bus[60]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_59_ ( .D(N329), .CP(CLK), .Q(
        o_data_bus[59]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_58_ ( .D(N328), .CP(CLK), .Q(
        o_data_bus[58]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_57_ ( .D(N327), .CP(CLK), .Q(
        o_data_bus[57]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_56_ ( .D(N326), .CP(CLK), .Q(
        o_data_bus[56]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_55_ ( .D(N325), .CP(CLK), .Q(
        o_data_bus[55]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_54_ ( .D(N324), .CP(CLK), .Q(
        o_data_bus[54]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_53_ ( .D(N323), .CP(CLK), .Q(
        o_data_bus[53]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_52_ ( .D(N322), .CP(CLK), .Q(
        o_data_bus[52]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_51_ ( .D(N321), .CP(CLK), .Q(
        o_data_bus[51]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_50_ ( .D(N320), .CP(CLK), .Q(
        o_data_bus[50]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_49_ ( .D(N236), .CP(CLK), .Q(
        o_data_bus[49]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_48_ ( .D(N235), .CP(CLK), .Q(
        o_data_bus[48]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_47_ ( .D(N234), .CP(CLK), .Q(
        o_data_bus[47]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_46_ ( .D(N233), .CP(CLK), .Q(
        o_data_bus[46]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_45_ ( .D(N232), .CP(CLK), .Q(
        o_data_bus[45]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_44_ ( .D(N231), .CP(CLK), .Q(
        o_data_bus[44]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_43_ ( .D(N230), .CP(CLK), .Q(
        o_data_bus[43]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_42_ ( .D(N229), .CP(CLK), .Q(
        o_data_bus[42]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_41_ ( .D(N228), .CP(CLK), .Q(
        o_data_bus[41]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_40_ ( .D(N227), .CP(CLK), .Q(
        o_data_bus[40]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_39_ ( .D(N226), .CP(CLK), .Q(
        o_data_bus[39]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_38_ ( .D(N225), .CP(CLK), .Q(
        o_data_bus[38]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_37_ ( .D(N224), .CP(CLK), .Q(
        o_data_bus[37]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_36_ ( .D(N223), .CP(CLK), .Q(
        o_data_bus[36]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_35_ ( .D(N222), .CP(CLK), .Q(
        o_data_bus[35]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_34_ ( .D(N221), .CP(CLK), .Q(
        o_data_bus[34]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_33_ ( .D(N220), .CP(CLK), .Q(
        o_data_bus[33]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_32_ ( .D(N219), .CP(CLK), .Q(
        o_data_bus[32]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_31_ ( .D(N218), .CP(CLK), .Q(
        o_data_bus[31]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_30_ ( .D(N217), .CP(CLK), .Q(
        o_data_bus[30]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_29_ ( .D(N216), .CP(CLK), .Q(
        o_data_bus[29]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_28_ ( .D(N215), .CP(CLK), .Q(
        o_data_bus[28]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_27_ ( .D(N214), .CP(CLK), .Q(
        o_data_bus[27]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_26_ ( .D(N213), .CP(CLK), .Q(
        o_data_bus[26]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_25_ ( .D(N212), .CP(CLK), .Q(
        o_data_bus[25]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_24_ ( .D(n177), .CP(CLK), .Q(
        o_data_bus[24]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_23_ ( .D(n176), .CP(CLK), .Q(
        o_data_bus[23]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_22_ ( .D(n175), .CP(CLK), .Q(
        o_data_bus[22]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_21_ ( .D(n174), .CP(CLK), .Q(
        o_data_bus[21]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_20_ ( .D(n173), .CP(CLK), .Q(
        o_data_bus[20]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_19_ ( .D(n172), .CP(CLK), .Q(
        o_data_bus[19]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_18_ ( .D(n171), .CP(CLK), .Q(
        o_data_bus[18]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_17_ ( .D(n170), .CP(CLK), .Q(
        o_data_bus[17]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_16_ ( .D(n169), .CP(CLK), .Q(
        o_data_bus[16]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_15_ ( .D(n168), .CP(CLK), .Q(
        o_data_bus[15]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_14_ ( .D(n167), .CP(CLK), .Q(
        o_data_bus[14]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_13_ ( .D(n166), .CP(CLK), .Q(
        o_data_bus[13]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_12_ ( .D(n228), .CP(CLK), .Q(
        o_data_bus[12]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_11_ ( .D(n227), .CP(CLK), .Q(
        o_data_bus[11]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_10_ ( .D(n226), .CP(CLK), .Q(
        o_data_bus[10]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_9_ ( .D(n225), .CP(CLK), .Q(
        o_data_bus[9]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_8_ ( .D(n224), .CP(CLK), .Q(
        o_data_bus[8]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_7_ ( .D(n223), .CP(CLK), .Q(
        o_data_bus[7]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_6_ ( .D(n222), .CP(CLK), .Q(
        o_data_bus[6]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_5_ ( .D(n221), .CP(CLK), .Q(
        o_data_bus[5]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_4_ ( .D(n220), .CP(CLK), .Q(
        o_data_bus[4]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_3_ ( .D(n219), .CP(CLK), .Q(
        o_data_bus[3]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_2_ ( .D(n218), .CP(CLK), .Q(
        o_data_bus[2]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_1_ ( .D(n217), .CP(CLK), .Q(
        o_data_bus[1]) );
  DFQD4BWP30P140LVT o_data_bus_reg_reg_0_ ( .D(n216), .CP(CLK), .Q(
        o_data_bus[0]) );
  NR3D1P5BWP30P140LVT U886 ( .A1(n38), .A2(o_cmd_forward_reg[36]), .A3(n37), 
        .ZN(n231) );
  NR3D1P5BWP30P140LVT U887 ( .A1(n29), .A2(o_cmd_forward_reg[20]), .A3(n28), 
        .ZN(n232) );
  NR3D1P5BWP30P140LVT U888 ( .A1(n32), .A2(o_cmd_forward_reg[50]), .A3(n31), 
        .ZN(n230) );
  NR3D1P5BWP30P140LVT U889 ( .A1(n26), .A2(n25), .A3(n24), .ZN(n234) );
  NR3D1P5BWP30P140LVT U890 ( .A1(n35), .A2(o_cmd_forward_reg[12]), .A3(n34), 
        .ZN(n233) );
  INVD2BWP30P140LVT U891 ( .I(n52), .ZN(n18) );
  CKAN2D1BWP30P140LVT U892 ( .A1(o_cmd_forward_reg[31]), .A2(n52), .Z(n245) );
  BUFFD2BWP30P140LVT U893 ( .I(n236), .Z(n20) );
  ND2D1BWP30P140LVT U894 ( .A1(n23), .A2(i_en), .ZN(n53) );
  NR2D1BWP30P140LVT U895 ( .A1(i_cmd[0]), .A2(i_cmd[1]), .ZN(n44) );
  ND2D1BWP30P140LVT U896 ( .A1(n250), .A2(n42), .ZN(n43) );
  NR2D1BWP30P140LVT U897 ( .A1(i_cmd[2]), .A2(i_cmd[3]), .ZN(n42) );
  INVD1BWP30P140LVT U898 ( .I(o_valid_forward_reg[2]), .ZN(n31) );
  ND2D1BWP30P140LVT U899 ( .A1(n30), .A2(n252), .ZN(n32) );
  AN4D1BWP30P140LVT U900 ( .A1(n253), .A2(n50), .A3(o_cmd_forward_reg[42]), 
        .A4(o_valid_forward_reg[4]), .Z(n238) );
  NR2D1BWP30P140LVT U901 ( .A1(o_cmd_forward_reg[41]), .A2(
        o_cmd_forward_reg[43]), .ZN(n50) );
  INVD1BWP30P140LVT U902 ( .I(o_cmd_forward_reg[38]), .ZN(n37) );
  ND2D1BWP30P140LVT U903 ( .A1(n36), .A2(n247), .ZN(n38) );
  CKBD1BWP30P140LVT U904 ( .I(n239), .Z(n19) );
  AN4D1BWP30P140LVT U905 ( .A1(n254), .A2(n51), .A3(o_cmd_forward_reg[27]), 
        .A4(o_valid_forward_reg[8]), .Z(n240) );
  NR2D1BWP30P140LVT U906 ( .A1(o_cmd_forward_reg[25]), .A2(
        o_cmd_forward_reg[26]), .ZN(n51) );
  INVD1BWP30P140LVT U907 ( .I(o_valid_forward_reg[9]), .ZN(n28) );
  ND2D1BWP30P140LVT U908 ( .A1(n27), .A2(n255), .ZN(n29) );
  AN4D1BWP30P140LVT U909 ( .A1(n47), .A2(n257), .A3(o_cmd_forward_reg[19]), 
        .A4(o_valid_forward_reg[10]), .Z(n241) );
  INVD1BWP30P140LVT U910 ( .I(o_valid_forward_reg[11]), .ZN(n34) );
  ND2D1BWP30P140LVT U911 ( .A1(n33), .A2(n259), .ZN(n35) );
  AN4D1BWP30P140LVT U912 ( .A1(n49), .A2(n258), .A3(o_cmd_forward_reg[10]), 
        .A4(o_valid_forward_reg[12]), .Z(n242) );
  AN4D1BWP30P140LVT U913 ( .A1(n48), .A2(n244), .A3(o_cmd_forward_reg[7]), 
        .A4(o_valid_forward_reg[13]), .Z(n243) );
  ND2D1BWP30P140LVT U914 ( .A1(o_cmd_forward_reg[2]), .A2(o_cmd_forward_reg[1]), .ZN(n26) );
  ND2D1BWP30P140LVT U915 ( .A1(o_valid_forward_reg[14]), .A2(
        o_cmd_forward_reg[3]), .ZN(n25) );
  ND2D1BWP30P140LVT U916 ( .A1(o_cmd_forward_reg[0]), .A2(n52), .ZN(n24) );
  INR2D1BWP30P140LVT U917 ( .A1(o_cmd_forward_reg[6]), .B1(n53), .ZN(n244) );
  INR2D1BWP30P140LVT U918 ( .A1(o_cmd_forward_reg[11]), .B1(n53), .ZN(n258) );
  INR2D1BWP30P140LVT U919 ( .A1(o_cmd_forward_reg[17]), .B1(n53), .ZN(n257) );
  INR2D1BWP30P140LVT U920 ( .A1(o_cmd_forward_reg[53]), .B1(n18), .ZN(n249) );
  INR4D0BWP30P140LVT U921 ( .A1(n245), .B1(o_cmd_forward_reg[29]), .B2(
        o_cmd_forward_reg[30]), .B3(n46), .ZN(n239) );
  INR4D0BWP30P140LVT U922 ( .A1(n249), .B1(o_cmd_forward_reg[54]), .B2(
        o_cmd_forward_reg[55]), .B3(n41), .ZN(n236) );
  CKAN2D1BWP30P140LVT U923 ( .A1(i_valid), .A2(n52), .Z(n250) );
  INR4D1BWP30P140LVT U924 ( .A1(n248), .B1(o_cmd_forward_reg[45]), .B2(
        o_cmd_forward_reg[47]), .B3(n40), .ZN(n21) );
  INR2D1BWP30P140LVT U925 ( .A1(o_cmd_forward_reg[46]), .B1(n53), .ZN(n248) );
  INR4D1BWP30P140LVT U926 ( .A1(n251), .B1(o_cmd_forward_reg[58]), .B2(
        o_cmd_forward_reg[59]), .B3(n45), .ZN(n22) );
  INR2D1BWP30P140LVT U927 ( .A1(o_cmd_forward_reg[56]), .B1(n53), .ZN(n251) );
  INVD1BWP30P140LVT U928 ( .I(n53), .ZN(n52) );
  INVD1BWP30P140LVT U929 ( .I(rst), .ZN(n23) );
  CKAN2D1BWP30P140LVT U930 ( .A1(i_data_bus[10]), .A2(n52), .Z(n188) );
  CKAN2D1BWP30P140LVT U931 ( .A1(i_data_bus[14]), .A2(n52), .Z(n192) );
  CKAN2D1BWP30P140LVT U932 ( .A1(i_data_bus[20]), .A2(n52), .Z(n198) );
  CKAN2D1BWP30P140LVT U933 ( .A1(i_data_bus[16]), .A2(n52), .Z(n194) );
  CKAN2D1BWP30P140LVT U934 ( .A1(i_data_bus[15]), .A2(n52), .Z(n193) );
  CKAN2D1BWP30P140LVT U935 ( .A1(i_data_bus[17]), .A2(n52), .Z(n195) );
  CKAN2D1BWP30P140LVT U936 ( .A1(i_data_bus[21]), .A2(n52), .Z(n199) );
  CKAN2D1BWP30P140LVT U937 ( .A1(i_data_bus[22]), .A2(n52), .Z(n200) );
  CKAN2D1BWP30P140LVT U938 ( .A1(i_data_bus[19]), .A2(n52), .Z(n197) );
  CKAN2D1BWP30P140LVT U939 ( .A1(i_data_bus[13]), .A2(n52), .Z(n191) );
  CKAN2D1BWP30P140LVT U940 ( .A1(i_data_bus[23]), .A2(n52), .Z(n201) );
  CKAN2D1BWP30P140LVT U941 ( .A1(i_data_bus[18]), .A2(n52), .Z(n196) );
  CKAN2D1BWP30P140LVT U942 ( .A1(i_data_bus[12]), .A2(n52), .Z(n190) );
  CKAN2D1BWP30P140LVT U943 ( .A1(i_data_bus[11]), .A2(n52), .Z(n189) );
  CKAN2D1BWP30P140LVT U944 ( .A1(i_data_bus[1]), .A2(n52), .Z(n179) );
  CKAN2D1BWP30P140LVT U945 ( .A1(i_data_bus[2]), .A2(n52), .Z(n180) );
  CKAN2D1BWP30P140LVT U946 ( .A1(i_data_bus[0]), .A2(n52), .Z(n178) );
  CKAN2D1BWP30P140LVT U947 ( .A1(i_data_bus[24]), .A2(n52), .Z(n202) );
  CKAN2D1BWP30P140LVT U948 ( .A1(i_data_bus[5]), .A2(n52), .Z(n183) );
  CKAN2D1BWP30P140LVT U949 ( .A1(i_data_bus[8]), .A2(n52), .Z(n186) );
  CKAN2D1BWP30P140LVT U950 ( .A1(i_data_bus[7]), .A2(n52), .Z(n185) );
  CKAN2D1BWP30P140LVT U951 ( .A1(i_data_bus[4]), .A2(n52), .Z(n182) );
  CKAN2D1BWP30P140LVT U952 ( .A1(i_data_bus[3]), .A2(n52), .Z(n181) );
  CKAN2D1BWP30P140LVT U953 ( .A1(i_data_bus[6]), .A2(n52), .Z(n184) );
  CKAN2D1BWP30P140LVT U954 ( .A1(i_data_bus[9]), .A2(n52), .Z(n187) );
  INR2D1BWP30P140LVT U955 ( .A1(o_cmd_forward_reg[21]), .B1(
        o_cmd_forward_reg[22]), .ZN(n27) );
  INR2D1BWP30P140LVT U956 ( .A1(o_cmd_forward_reg[23]), .B1(n18), .ZN(n255) );
  INR2D1BWP30P140LVT U957 ( .A1(o_cmd_forward_reg[48]), .B1(
        o_cmd_forward_reg[51]), .ZN(n30) );
  INR2D1BWP30P140LVT U958 ( .A1(o_cmd_forward_reg[49]), .B1(n18), .ZN(n252) );
  INR2D1BWP30P140LVT U959 ( .A1(o_cmd_forward_reg[14]), .B1(
        o_cmd_forward_reg[13]), .ZN(n33) );
  INR2D1BWP30P140LVT U960 ( .A1(o_cmd_forward_reg[15]), .B1(n53), .ZN(n259) );
  INR2D1BWP30P140LVT U961 ( .A1(o_valid_forward_reg[5]), .B1(
        o_cmd_forward_reg[39]), .ZN(n36) );
  INR2D1BWP30P140LVT U962 ( .A1(o_cmd_forward_reg[37]), .B1(n18), .ZN(n247) );
  INR2D1BWP30P140LVT U963 ( .A1(o_cmd_forward_reg[34]), .B1(n53), .ZN(n256) );
  ND3D1BWP30P140LVT U964 ( .A1(n256), .A2(o_cmd_forward_reg[33]), .A3(
        o_cmd_forward_reg[32]), .ZN(n39) );
  INR3D2BWP30P140LVT U965 ( .A1(o_valid_forward_reg[6]), .B1(
        o_cmd_forward_reg[35]), .B2(n39), .ZN(n246) );
  IND2D1BWP30P140LVT U966 ( .A1(o_cmd_forward_reg[44]), .B1(
        o_valid_forward_reg[3]), .ZN(n40) );
  INR4D1BWP30P140LVT U967 ( .A1(n248), .B1(o_cmd_forward_reg[45]), .B2(
        o_cmd_forward_reg[47]), .B3(n40), .ZN(n237) );
  IND2D1BWP30P140LVT U968 ( .A1(o_cmd_forward_reg[52]), .B1(
        o_valid_forward_reg[1]), .ZN(n41) );
  INR2D2BWP30P140LVT U969 ( .A1(n44), .B1(n43), .ZN(n229) );
  IND2D1BWP30P140LVT U970 ( .A1(o_cmd_forward_reg[57]), .B1(
        o_valid_forward_reg[0]), .ZN(n45) );
  INR4D1BWP30P140LVT U971 ( .A1(n251), .B1(o_cmd_forward_reg[58]), .B2(
        o_cmd_forward_reg[59]), .B3(n45), .ZN(n235) );
  IND2D1BWP30P140LVT U972 ( .A1(o_cmd_forward_reg[28]), .B1(
        o_valid_forward_reg[7]), .ZN(n46) );
  INR2D1BWP30P140LVT U973 ( .A1(o_cmd_forward_reg[16]), .B1(
        o_cmd_forward_reg[18]), .ZN(n47) );
  INR2D1BWP30P140LVT U974 ( .A1(o_cmd_forward_reg[5]), .B1(
        o_cmd_forward_reg[4]), .ZN(n48) );
  INR2D1BWP30P140LVT U975 ( .A1(o_cmd_forward_reg[8]), .B1(
        o_cmd_forward_reg[9]), .ZN(n49) );
  INR2D1BWP30P140LVT U976 ( .A1(o_cmd_forward_reg[40]), .B1(n53), .ZN(n253) );
  INR2D1BWP30P140LVT U977 ( .A1(o_cmd_forward_reg[24]), .B1(n53), .ZN(n254) );
  INR2D1BWP30P140LVT U978 ( .A1(o_data_forward_reg[374]), .B1(n53), .ZN(N261)
         );
  INR2D1BWP30P140LVT U979 ( .A1(o_data_forward_reg[302]), .B1(n53), .ZN(N455)
         );
  INR2D1BWP30P140LVT U980 ( .A1(o_data_forward_reg[371]), .B1(n18), .ZN(N258)
         );
  INR2D1BWP30P140LVT U981 ( .A1(o_data_forward_reg[370]), .B1(n18), .ZN(N257)
         );
  INR2D1BWP30P140LVT U982 ( .A1(o_data_forward_reg[369]), .B1(n53), .ZN(N256)
         );
  INR2D1BWP30P140LVT U983 ( .A1(o_data_forward_reg[368]), .B1(n18), .ZN(N255)
         );
  INR2D1BWP30P140LVT U984 ( .A1(o_data_forward_reg[367]), .B1(n53), .ZN(N254)
         );
  INR2D1BWP30P140LVT U985 ( .A1(o_data_forward_reg[366]), .B1(n18), .ZN(N253)
         );
  INR2D1BWP30P140LVT U986 ( .A1(o_data_forward_reg[365]), .B1(n18), .ZN(N252)
         );
  INR2D1BWP30P140LVT U987 ( .A1(o_data_forward_reg[364]), .B1(n53), .ZN(N251)
         );
  INR2D1BWP30P140LVT U988 ( .A1(o_data_forward_reg[363]), .B1(n53), .ZN(N250)
         );
  INR2D1BWP30P140LVT U989 ( .A1(o_data_forward_reg[362]), .B1(n53), .ZN(N249)
         );
  INR2D1BWP30P140LVT U990 ( .A1(o_data_forward_reg[361]), .B1(n18), .ZN(N248)
         );
  INR2D1BWP30P140LVT U991 ( .A1(o_data_forward_reg[360]), .B1(n18), .ZN(N247)
         );
  INR2D1BWP30P140LVT U992 ( .A1(o_data_forward_reg[359]), .B1(n18), .ZN(N246)
         );
  INR2D1BWP30P140LVT U993 ( .A1(o_data_forward_reg[358]), .B1(n18), .ZN(N245)
         );
  INR2D1BWP30P140LVT U994 ( .A1(o_data_forward_reg[357]), .B1(n18), .ZN(N244)
         );
  INR2D1BWP30P140LVT U995 ( .A1(o_data_forward_reg[356]), .B1(n18), .ZN(N243)
         );
  INR2D1BWP30P140LVT U996 ( .A1(o_data_forward_reg[355]), .B1(n18), .ZN(N242)
         );
  INR2D1BWP30P140LVT U997 ( .A1(o_data_forward_reg[372]), .B1(n18), .ZN(N259)
         );
  INR2D1BWP30P140LVT U998 ( .A1(o_data_forward_reg[303]), .B1(n18), .ZN(N456)
         );
  INR2D1BWP30P140LVT U999 ( .A1(o_data_forward_reg[348]), .B1(n18), .ZN(N368)
         );
  INR2D1BWP30P140LVT U1000 ( .A1(o_data_forward_reg[373]), .B1(n18), .ZN(N260)
         );
  INR2D1BWP30P140LVT U1001 ( .A1(o_data_forward_reg[346]), .B1(n53), .ZN(N366)
         );
  INR2D1BWP30P140LVT U1002 ( .A1(o_data_forward_reg[345]), .B1(n53), .ZN(N365)
         );
  INR2D1BWP30P140LVT U1003 ( .A1(o_data_forward_reg[344]), .B1(n53), .ZN(N364)
         );
  INR2D1BWP30P140LVT U1004 ( .A1(o_data_forward_reg[325]), .B1(n18), .ZN(N345)
         );
  INR2D1BWP30P140LVT U1005 ( .A1(o_data_forward_reg[326]), .B1(n53), .ZN(N346)
         );
  INR2D1BWP30P140LVT U1006 ( .A1(o_data_forward_reg[349]), .B1(n53), .ZN(N369)
         );
  INR2D1BWP30P140LVT U1007 ( .A1(o_data_forward_reg[300]), .B1(n18), .ZN(N453)
         );
  INR2D1BWP30P140LVT U1008 ( .A1(o_data_forward_reg[347]), .B1(n18), .ZN(N367)
         );
  INR2D1BWP30P140LVT U1009 ( .A1(o_data_forward_reg[330]), .B1(n53), .ZN(N350)
         );
  INR2D1BWP30P140LVT U1010 ( .A1(o_data_forward_reg[329]), .B1(n18), .ZN(N349)
         );
  INR2D1BWP30P140LVT U1011 ( .A1(o_data_forward_reg[328]), .B1(n18), .ZN(N348)
         );
  INR2D1BWP30P140LVT U1012 ( .A1(o_data_forward_reg[327]), .B1(n18), .ZN(N347)
         );
  INR2D1BWP30P140LVT U1013 ( .A1(o_data_forward_reg[305]), .B1(n18), .ZN(N458)
         );
  INR2D1BWP30P140LVT U1014 ( .A1(o_data_forward_reg[301]), .B1(n53), .ZN(N454)
         );
  INR2D1BWP30P140LVT U1015 ( .A1(o_data_forward_reg[304]), .B1(n18), .ZN(N457)
         );
  INR2D1BWP30P140LVT U1016 ( .A1(o_data_forward_reg[144]), .B1(n18), .ZN(N1228) );
  INR2D1BWP30P140LVT U1017 ( .A1(o_data_forward_reg[138]), .B1(n18), .ZN(N1222) );
  INR2D1BWP30P140LVT U1018 ( .A1(o_data_forward_reg[141]), .B1(n53), .ZN(N1225) );
  INR2D1BWP30P140LVT U1019 ( .A1(o_data_forward_reg[140]), .B1(n53), .ZN(N1224) );
  INR2D1BWP30P140LVT U1020 ( .A1(o_data_forward_reg[139]), .B1(n53), .ZN(N1223) );
  INR2D1BWP30P140LVT U1021 ( .A1(o_data_forward_reg[149]), .B1(n18), .ZN(N1233) );
  INR2D1BWP30P140LVT U1022 ( .A1(o_data_forward_reg[118]), .B1(n53), .ZN(N1335) );
  INR2D1BWP30P140LVT U1023 ( .A1(o_data_forward_reg[117]), .B1(n18), .ZN(N1334) );
  INR2D1BWP30P140LVT U1024 ( .A1(o_data_forward_reg[145]), .B1(n18), .ZN(N1229) );
  INR2D1BWP30P140LVT U1025 ( .A1(o_data_forward_reg[142]), .B1(n18), .ZN(N1226) );
  INR2D1BWP30P140LVT U1026 ( .A1(o_data_forward_reg[143]), .B1(n18), .ZN(N1227) );
  INR2D1BWP30P140LVT U1027 ( .A1(o_data_forward_reg[121]), .B1(n18), .ZN(N1338) );
  INR2D1BWP30P140LVT U1028 ( .A1(o_data_forward_reg[120]), .B1(n53), .ZN(N1337) );
  INR2D1BWP30P140LVT U1029 ( .A1(o_data_forward_reg[119]), .B1(n18), .ZN(N1336) );
  INR2D1BWP30P140LVT U1030 ( .A1(o_data_forward_reg[147]), .B1(n18), .ZN(N1231) );
  INR2D1BWP30P140LVT U1031 ( .A1(o_data_forward_reg[115]), .B1(n53), .ZN(N1332) );
  INR2D1BWP30P140LVT U1032 ( .A1(o_data_forward_reg[116]), .B1(n18), .ZN(N1333) );
  INR2D1BWP30P140LVT U1033 ( .A1(o_data_forward_reg[123]), .B1(n53), .ZN(N1340) );
  INR2D1BWP30P140LVT U1034 ( .A1(o_data_forward_reg[124]), .B1(n18), .ZN(N1341) );
  INR2D1BWP30P140LVT U1035 ( .A1(o_data_forward_reg[111]), .B1(n18), .ZN(N1328) );
  INR2D1BWP30P140LVT U1036 ( .A1(o_data_forward_reg[110]), .B1(n18), .ZN(N1327) );
  INR2D1BWP30P140LVT U1037 ( .A1(o_data_forward_reg[146]), .B1(n18), .ZN(N1230) );
  INR2D1BWP30P140LVT U1038 ( .A1(o_data_forward_reg[109]), .B1(n18), .ZN(N1326) );
  INR2D1BWP30P140LVT U1039 ( .A1(o_data_forward_reg[108]), .B1(n53), .ZN(N1325) );
  INR2D1BWP30P140LVT U1040 ( .A1(o_data_forward_reg[107]), .B1(n18), .ZN(N1324) );
  INR2D1BWP30P140LVT U1041 ( .A1(o_data_forward_reg[106]), .B1(n18), .ZN(N1323) );
  INR2D1BWP30P140LVT U1042 ( .A1(o_data_forward_reg[105]), .B1(n18), .ZN(N1322) );
  INR2D1BWP30P140LVT U1043 ( .A1(o_data_forward_reg[104]), .B1(n18), .ZN(N1321) );
  INR2D1BWP30P140LVT U1044 ( .A1(o_data_forward_reg[103]), .B1(n18), .ZN(N1320) );
  INR2D1BWP30P140LVT U1045 ( .A1(o_data_forward_reg[102]), .B1(n18), .ZN(N1319) );
  INR2D1BWP30P140LVT U1046 ( .A1(o_data_forward_reg[101]), .B1(n18), .ZN(N1318) );
  INR2D1BWP30P140LVT U1047 ( .A1(o_data_forward_reg[100]), .B1(n18), .ZN(N1317) );
  INR2D1BWP30P140LVT U1048 ( .A1(o_data_forward_reg[99]), .B1(n18), .ZN(N1449)
         );
  INR2D1BWP30P140LVT U1049 ( .A1(o_data_forward_reg[98]), .B1(n53), .ZN(N1448)
         );
  INR2D1BWP30P140LVT U1050 ( .A1(o_data_forward_reg[114]), .B1(n53), .ZN(N1331) );
  INR2D1BWP30P140LVT U1051 ( .A1(o_data_forward_reg[113]), .B1(n18), .ZN(N1330) );
  INR2D1BWP30P140LVT U1052 ( .A1(o_data_forward_reg[112]), .B1(n18), .ZN(N1329) );
  INR2D1BWP30P140LVT U1053 ( .A1(o_data_forward_reg[137]), .B1(n18), .ZN(N1221) );
  INR2D1BWP30P140LVT U1054 ( .A1(o_data_forward_reg[136]), .B1(n18), .ZN(N1220) );
  INR2D1BWP30P140LVT U1055 ( .A1(o_data_forward_reg[148]), .B1(n18), .ZN(N1232) );
  INR2D1BWP30P140LVT U1056 ( .A1(o_data_forward_reg[97]), .B1(n53), .ZN(N1447)
         );
  INR2D1BWP30P140LVT U1057 ( .A1(o_data_forward_reg[96]), .B1(n53), .ZN(N1446)
         );
  INR2D1BWP30P140LVT U1058 ( .A1(o_data_forward_reg[122]), .B1(n53), .ZN(N1339) );
  INR2D1BWP30P140LVT U1059 ( .A1(o_data_forward_reg[95]), .B1(n53), .ZN(N1445)
         );
  INR2D1BWP30P140LVT U1060 ( .A1(o_data_forward_reg[94]), .B1(n18), .ZN(N1444)
         );
  INR2D1BWP30P140LVT U1061 ( .A1(o_data_forward_reg[93]), .B1(n53), .ZN(N1443)
         );
  INR2D1BWP30P140LVT U1062 ( .A1(o_data_forward_reg[92]), .B1(n18), .ZN(N1442)
         );
  INR2D1BWP30P140LVT U1063 ( .A1(o_data_forward_reg[80]), .B1(n53), .ZN(N1430)
         );
  INR2D1BWP30P140LVT U1064 ( .A1(o_data_forward_reg[91]), .B1(n18), .ZN(N1441)
         );
  INR2D1BWP30P140LVT U1065 ( .A1(o_data_forward_reg[90]), .B1(n53), .ZN(N1440)
         );
  INR2D1BWP30P140LVT U1066 ( .A1(o_data_forward_reg[89]), .B1(n18), .ZN(N1439)
         );
  INR2D1BWP30P140LVT U1067 ( .A1(o_data_forward_reg[88]), .B1(n18), .ZN(N1438)
         );
  INR2D1BWP30P140LVT U1068 ( .A1(o_data_forward_reg[87]), .B1(n18), .ZN(N1437)
         );
  INR2D1BWP30P140LVT U1069 ( .A1(o_data_forward_reg[86]), .B1(n18), .ZN(N1436)
         );
  INR2D1BWP30P140LVT U1070 ( .A1(o_data_forward_reg[85]), .B1(n18), .ZN(N1435)
         );
  INR2D1BWP30P140LVT U1071 ( .A1(o_data_forward_reg[84]), .B1(n18), .ZN(N1434)
         );
  INR2D1BWP30P140LVT U1072 ( .A1(o_data_forward_reg[83]), .B1(n53), .ZN(N1433)
         );
  INR2D1BWP30P140LVT U1073 ( .A1(o_data_forward_reg[82]), .B1(n18), .ZN(N1432)
         );
  INR2D1BWP30P140LVT U1074 ( .A1(o_data_forward_reg[81]), .B1(n53), .ZN(N1431)
         );
  INR2D1BWP30P140LVT U1075 ( .A1(o_data_forward_reg[60]), .B1(n18), .ZN(N1543)
         );
  INR2D1BWP30P140LVT U1076 ( .A1(o_data_forward_reg[59]), .B1(n53), .ZN(N1542)
         );
  INR2D1BWP30P140LVT U1077 ( .A1(o_data_forward_reg[79]), .B1(n53), .ZN(N1429)
         );
  INR2D1BWP30P140LVT U1078 ( .A1(o_data_forward_reg[78]), .B1(n18), .ZN(N1428)
         );
  INR2D1BWP30P140LVT U1079 ( .A1(o_data_forward_reg[77]), .B1(n18), .ZN(N1427)
         );
  INR2D1BWP30P140LVT U1080 ( .A1(o_data_forward_reg[76]), .B1(n53), .ZN(N1426)
         );
  INR2D1BWP30P140LVT U1081 ( .A1(o_data_forward_reg[75]), .B1(n18), .ZN(N1425)
         );
  INR2D1BWP30P140LVT U1082 ( .A1(o_data_forward_reg[54]), .B1(n18), .ZN(N1537)
         );
  INR2D1BWP30P140LVT U1083 ( .A1(o_data_forward_reg[51]), .B1(n53), .ZN(N1534)
         );
  INR2D1BWP30P140LVT U1084 ( .A1(o_data_forward_reg[53]), .B1(n18), .ZN(N1536)
         );
  INR2D1BWP30P140LVT U1085 ( .A1(o_data_forward_reg[52]), .B1(n53), .ZN(N1535)
         );
  INR2D1BWP30P140LVT U1086 ( .A1(o_data_forward_reg[58]), .B1(n18), .ZN(N1541)
         );
  INR2D1BWP30P140LVT U1087 ( .A1(o_data_forward_reg[57]), .B1(n18), .ZN(N1540)
         );
  INR2D1BWP30P140LVT U1088 ( .A1(o_data_forward_reg[56]), .B1(n18), .ZN(N1539)
         );
  INR2D1BWP30P140LVT U1089 ( .A1(o_data_forward_reg[50]), .B1(n18), .ZN(N1533)
         );
  INR2D1BWP30P140LVT U1090 ( .A1(o_data_forward_reg[55]), .B1(n18), .ZN(N1538)
         );
  INR2D1BWP30P140LVT U1091 ( .A1(o_data_forward_reg[62]), .B1(n18), .ZN(N1545)
         );
  INR2D1BWP30P140LVT U1092 ( .A1(o_data_forward_reg[61]), .B1(n18), .ZN(N1544)
         );
  INR2D1BWP30P140LVT U1093 ( .A1(o_data_forward_reg[350]), .B1(n18), .ZN(N237)
         );
  INR2D1BWP30P140LVT U1094 ( .A1(o_data_forward_reg[353]), .B1(n18), .ZN(N240)
         );
  INR2D1BWP30P140LVT U1095 ( .A1(o_cmd_forward_reg[16]), .B1(n18), .ZN(N1343)
         );
  INR2D1BWP30P140LVT U1096 ( .A1(o_cmd_forward_reg[8]), .B1(n18), .ZN(N1559)
         );
  INR2D1BWP30P140LVT U1097 ( .A1(o_data_forward_reg[67]), .B1(n53), .ZN(N1550)
         );
  INR2D1BWP30P140LVT U1098 ( .A1(o_data_forward_reg[65]), .B1(n53), .ZN(N1548)
         );
  INR2D1BWP30P140LVT U1099 ( .A1(o_data_forward_reg[64]), .B1(n18), .ZN(N1547)
         );
  INR2D1BWP30P140LVT U1100 ( .A1(o_data_forward_reg[63]), .B1(n53), .ZN(N1546)
         );
  INR2D1BWP30P140LVT U1101 ( .A1(o_data_forward_reg[66]), .B1(n53), .ZN(N1549)
         );
  INR2D1BWP30P140LVT U1102 ( .A1(o_data_forward_reg[74]), .B1(n18), .ZN(N1557)
         );
  INR2D1BWP30P140LVT U1103 ( .A1(o_data_forward_reg[73]), .B1(n53), .ZN(N1556)
         );
  INR2D1BWP30P140LVT U1104 ( .A1(o_data_forward_reg[72]), .B1(n18), .ZN(N1555)
         );
  INR2D1BWP30P140LVT U1105 ( .A1(o_data_forward_reg[71]), .B1(n18), .ZN(N1554)
         );
  INR2D1BWP30P140LVT U1106 ( .A1(o_data_forward_reg[70]), .B1(n18), .ZN(N1553)
         );
  INR2D1BWP30P140LVT U1107 ( .A1(o_data_forward_reg[69]), .B1(n53), .ZN(N1552)
         );
  INR2D1BWP30P140LVT U1108 ( .A1(o_data_forward_reg[68]), .B1(n53), .ZN(N1551)
         );
  INR2D1BWP30P140LVT U1109 ( .A1(o_data_forward_reg[25]), .B1(n18), .ZN(N1641)
         );
  INR2D1BWP30P140LVT U1110 ( .A1(o_data_forward_reg[341]), .B1(n18), .ZN(N361)
         );
  INR2D1BWP30P140LVT U1111 ( .A1(o_data_forward_reg[340]), .B1(n18), .ZN(N360)
         );
  INR2D1BWP30P140LVT U1112 ( .A1(o_data_forward_reg[339]), .B1(n18), .ZN(N359)
         );
  INR2D1BWP30P140LVT U1113 ( .A1(o_data_forward_reg[338]), .B1(n53), .ZN(N358)
         );
  INR2D1BWP30P140LVT U1114 ( .A1(o_data_forward_reg[337]), .B1(n18), .ZN(N357)
         );
  INR2D1BWP30P140LVT U1115 ( .A1(o_data_forward_reg[336]), .B1(n53), .ZN(N356)
         );
  INR2D1BWP30P140LVT U1116 ( .A1(o_data_forward_reg[335]), .B1(n18), .ZN(N355)
         );
  INR2D1BWP30P140LVT U1117 ( .A1(o_data_forward_reg[334]), .B1(n18), .ZN(N354)
         );
  INR2D1BWP30P140LVT U1118 ( .A1(o_data_forward_reg[333]), .B1(n53), .ZN(N353)
         );
  INR2D1BWP30P140LVT U1119 ( .A1(o_data_forward_reg[343]), .B1(n18), .ZN(N363)
         );
  INR2D1BWP30P140LVT U1120 ( .A1(o_data_forward_reg[342]), .B1(n18), .ZN(N362)
         );
  INR2D1BWP30P140LVT U1121 ( .A1(o_data_forward_reg[331]), .B1(n18), .ZN(N351)
         );
  INR2D1BWP30P140LVT U1122 ( .A1(o_data_forward_reg[332]), .B1(n18), .ZN(N352)
         );
  INR2D1BWP30P140LVT U1123 ( .A1(o_data_forward_reg[26]), .B1(n18), .ZN(N1642)
         );
  INR2D1BWP30P140LVT U1124 ( .A1(o_data_forward_reg[27]), .B1(n18), .ZN(N1643)
         );
  INR2D1BWP30P140LVT U1125 ( .A1(o_data_forward_reg[33]), .B1(n18), .ZN(N1649)
         );
  INR2D1BWP30P140LVT U1126 ( .A1(o_data_forward_reg[29]), .B1(n53), .ZN(N1645)
         );
  INR2D1BWP30P140LVT U1127 ( .A1(o_data_forward_reg[30]), .B1(n53), .ZN(N1646)
         );
  INR2D1BWP30P140LVT U1128 ( .A1(o_data_forward_reg[31]), .B1(n18), .ZN(N1647)
         );
  INR2D1BWP30P140LVT U1129 ( .A1(o_data_forward_reg[28]), .B1(n18), .ZN(N1644)
         );
  INR2D1BWP30P140LVT U1130 ( .A1(o_data_forward_reg[352]), .B1(n18), .ZN(N239)
         );
  INR2D1BWP30P140LVT U1131 ( .A1(o_data_forward_reg[34]), .B1(n53), .ZN(N1650)
         );
  INR2D1BWP30P140LVT U1132 ( .A1(o_data_forward_reg[35]), .B1(n18), .ZN(N1651)
         );
  INR2D1BWP30P140LVT U1133 ( .A1(o_data_forward_reg[32]), .B1(n18), .ZN(N1648)
         );
  INR2D1BWP30P140LVT U1134 ( .A1(o_data_forward_reg[37]), .B1(n18), .ZN(N1653)
         );
  INR2D1BWP30P140LVT U1135 ( .A1(o_data_forward_reg[38]), .B1(n18), .ZN(N1654)
         );
  INR2D1BWP30P140LVT U1136 ( .A1(o_data_forward_reg[36]), .B1(n18), .ZN(N1652)
         );
  INR2D1BWP30P140LVT U1137 ( .A1(o_data_forward_reg[45]), .B1(n53), .ZN(N1661)
         );
  INR2D1BWP30P140LVT U1138 ( .A1(o_data_forward_reg[41]), .B1(n53), .ZN(N1657)
         );
  INR2D1BWP30P140LVT U1139 ( .A1(o_data_forward_reg[47]), .B1(n18), .ZN(N1663)
         );
  INR2D1BWP30P140LVT U1140 ( .A1(o_data_forward_reg[43]), .B1(n53), .ZN(N1659)
         );
  INR2D1BWP30P140LVT U1141 ( .A1(o_data_forward_reg[351]), .B1(n53), .ZN(N238)
         );
  INR2D1BWP30P140LVT U1142 ( .A1(o_data_forward_reg[48]), .B1(n18), .ZN(N1664)
         );
  INR2D1BWP30P140LVT U1143 ( .A1(o_data_forward_reg[46]), .B1(n18), .ZN(N1662)
         );
  INR2D1BWP30P140LVT U1144 ( .A1(o_data_forward_reg[44]), .B1(n18), .ZN(N1660)
         );
  INR2D1BWP30P140LVT U1145 ( .A1(o_data_forward_reg[39]), .B1(n53), .ZN(N1655)
         );
  INR2D1BWP30P140LVT U1146 ( .A1(o_data_forward_reg[49]), .B1(n53), .ZN(N1665)
         );
  INR2D1BWP30P140LVT U1147 ( .A1(o_data_forward_reg[354]), .B1(n18), .ZN(N241)
         );
  INR2D1BWP30P140LVT U1148 ( .A1(o_data_forward_reg[40]), .B1(n18), .ZN(N1656)
         );
  INR2D1BWP30P140LVT U1149 ( .A1(o_data_forward_reg[42]), .B1(n18), .ZN(N1658)
         );
  INR2D1BWP30P140LVT U1150 ( .A1(o_data_forward_reg[249]), .B1(n18), .ZN(N801)
         );
  INR2D1BWP30P140LVT U1151 ( .A1(o_data_forward_reg[248]), .B1(n18), .ZN(N800)
         );
  INR2D1BWP30P140LVT U1152 ( .A1(o_data_forward_reg[247]), .B1(n18), .ZN(N799)
         );
  INR2D1BWP30P140LVT U1153 ( .A1(o_data_forward_reg[246]), .B1(n18), .ZN(N798)
         );
  INR2D1BWP30P140LVT U1154 ( .A1(o_data_forward_reg[224]), .B1(n18), .ZN(N909)
         );
  INR2D1BWP30P140LVT U1155 ( .A1(o_data_forward_reg[222]), .B1(n18), .ZN(N907)
         );
  INR2D1BWP30P140LVT U1156 ( .A1(o_data_forward_reg[200]), .B1(n18), .ZN(N885)
         );
  INR2D1BWP30P140LVT U1157 ( .A1(o_data_forward_reg[205]), .B1(n18), .ZN(N890)
         );
  INR2D1BWP30P140LVT U1158 ( .A1(o_data_forward_reg[180]), .B1(n18), .ZN(N998)
         );
  INR2D1BWP30P140LVT U1159 ( .A1(o_data_forward_reg[202]), .B1(n18), .ZN(N887)
         );
  INR2D1BWP30P140LVT U1160 ( .A1(o_data_forward_reg[178]), .B1(n18), .ZN(N996)
         );
  INR2D1BWP30P140LVT U1161 ( .A1(o_data_forward_reg[201]), .B1(n18), .ZN(N886)
         );
  INR2D1BWP30P140LVT U1162 ( .A1(o_data_forward_reg[175]), .B1(n18), .ZN(N993)
         );
  INR2D1BWP30P140LVT U1163 ( .A1(o_data_forward_reg[192]), .B1(n18), .ZN(N1010) );
  INR2D1BWP30P140LVT U1164 ( .A1(o_data_forward_reg[203]), .B1(n18), .ZN(N888)
         );
  INR2D1BWP30P140LVT U1165 ( .A1(o_data_forward_reg[164]), .B1(n18), .ZN(N1115) );
  INR2D1BWP30P140LVT U1166 ( .A1(o_data_forward_reg[161]), .B1(n18), .ZN(N1112) );
  INR2D1BWP30P140LVT U1167 ( .A1(o_data_forward_reg[170]), .B1(n18), .ZN(N1121) );
  INR2D1BWP30P140LVT U1168 ( .A1(o_data_forward_reg[206]), .B1(n18), .ZN(N891)
         );
  INR2D1BWP30P140LVT U1169 ( .A1(o_data_forward_reg[207]), .B1(n18), .ZN(N892)
         );
  INR2D1BWP30P140LVT U1170 ( .A1(o_data_forward_reg[204]), .B1(n18), .ZN(N889)
         );
  INR2D1BWP30P140LVT U1171 ( .A1(o_data_forward_reg[167]), .B1(n18), .ZN(N1118) );
  INR2D1BWP30P140LVT U1172 ( .A1(o_data_forward_reg[194]), .B1(n18), .ZN(N1012) );
  INR2D1BWP30P140LVT U1173 ( .A1(o_data_forward_reg[193]), .B1(n18), .ZN(N1011) );
  INR2D1BWP30P140LVT U1174 ( .A1(o_data_forward_reg[158]), .B1(n18), .ZN(N1109) );
  INR2D1BWP30P140LVT U1175 ( .A1(o_data_forward_reg[154]), .B1(n18), .ZN(N1105) );
  INR2D1BWP30P140LVT U1176 ( .A1(o_data_forward_reg[150]), .B1(n18), .ZN(N1101) );
  INR2D1BWP30P140LVT U1177 ( .A1(o_data_forward_reg[155]), .B1(n18), .ZN(N1106) );
  INR2D1BWP30P140LVT U1178 ( .A1(o_data_forward_reg[187]), .B1(n18), .ZN(N1005) );
  INR2D1BWP30P140LVT U1179 ( .A1(o_data_forward_reg[131]), .B1(n18), .ZN(N1215) );
  INR2D1BWP30P140LVT U1180 ( .A1(o_data_forward_reg[128]), .B1(n53), .ZN(N1212) );
  INR2D1BWP30P140LVT U1181 ( .A1(o_data_forward_reg[132]), .B1(n18), .ZN(N1216) );
  INR2D1BWP30P140LVT U1182 ( .A1(o_data_forward_reg[126]), .B1(n18), .ZN(N1210) );
  INR2D1BWP30P140LVT U1183 ( .A1(o_data_forward_reg[191]), .B1(n18), .ZN(N1009) );
  INR2D1BWP30P140LVT U1184 ( .A1(o_data_forward_reg[221]), .B1(n53), .ZN(N906)
         );
  INR2D1BWP30P140LVT U1185 ( .A1(o_data_forward_reg[183]), .B1(n53), .ZN(N1001) );
  INR2D1BWP30P140LVT U1186 ( .A1(o_data_forward_reg[127]), .B1(n18), .ZN(N1211) );
  INR2D1BWP30P140LVT U1187 ( .A1(o_data_forward_reg[133]), .B1(n18), .ZN(N1217) );
  INR2D1BWP30P140LVT U1188 ( .A1(o_data_forward_reg[130]), .B1(n53), .ZN(N1214) );
  INR2D1BWP30P140LVT U1189 ( .A1(o_data_forward_reg[189]), .B1(n18), .ZN(N1007) );
  INR2D1BWP30P140LVT U1190 ( .A1(o_data_forward_reg[134]), .B1(n18), .ZN(N1218) );
  INR2D1BWP30P140LVT U1191 ( .A1(o_data_forward_reg[179]), .B1(n18), .ZN(N997)
         );
  INR2D1BWP30P140LVT U1192 ( .A1(o_data_forward_reg[174]), .B1(n53), .ZN(N1125) );
  INR2D1BWP30P140LVT U1193 ( .A1(o_data_forward_reg[166]), .B1(n18), .ZN(N1117) );
  INR2D1BWP30P140LVT U1194 ( .A1(o_data_forward_reg[172]), .B1(n18), .ZN(N1123) );
  INR2D1BWP30P140LVT U1195 ( .A1(o_data_forward_reg[129]), .B1(n18), .ZN(N1213) );
  INR2D1BWP30P140LVT U1196 ( .A1(o_data_forward_reg[186]), .B1(n53), .ZN(N1004) );
  INR2D1BWP30P140LVT U1197 ( .A1(o_data_forward_reg[157]), .B1(n53), .ZN(N1108) );
  INR2D1BWP30P140LVT U1198 ( .A1(o_data_forward_reg[173]), .B1(n18), .ZN(N1124) );
  INR2D1BWP30P140LVT U1199 ( .A1(o_data_forward_reg[196]), .B1(n18), .ZN(N1014) );
  INR2D1BWP30P140LVT U1200 ( .A1(o_data_forward_reg[153]), .B1(n53), .ZN(N1104) );
  INR2D1BWP30P140LVT U1201 ( .A1(o_data_forward_reg[135]), .B1(n18), .ZN(N1219) );
  INR2D1BWP30P140LVT U1202 ( .A1(o_data_forward_reg[199]), .B1(n18), .ZN(N1017) );
  INR2D1BWP30P140LVT U1203 ( .A1(o_data_forward_reg[151]), .B1(n18), .ZN(N1102) );
  INR2D1BWP30P140LVT U1204 ( .A1(o_data_forward_reg[188]), .B1(n53), .ZN(N1006) );
  INR2D1BWP30P140LVT U1205 ( .A1(o_data_forward_reg[163]), .B1(n18), .ZN(N1114) );
  INR2D1BWP30P140LVT U1206 ( .A1(o_data_forward_reg[169]), .B1(n18), .ZN(N1120) );
  INR2D1BWP30P140LVT U1207 ( .A1(o_data_forward_reg[160]), .B1(n18), .ZN(N1111) );
  INR2D1BWP30P140LVT U1208 ( .A1(o_data_forward_reg[177]), .B1(n53), .ZN(N995)
         );
  INR2D1BWP30P140LVT U1209 ( .A1(o_data_forward_reg[125]), .B1(n53), .ZN(N1209) );
  INR2D1BWP30P140LVT U1210 ( .A1(o_cmd_forward_reg[21]), .B1(n18), .ZN(N1236)
         );
  INR2D1BWP30P140LVT U1211 ( .A1(o_valid_forward_reg[5]), .B1(n18), .ZN(N802)
         );
  INR2D1BWP30P140LVT U1212 ( .A1(o_cmd_forward_reg[5]), .B1(n18), .ZN(N1668)
         );
  INR2D1BWP30P140LVT U1213 ( .A1(o_cmd_forward_reg[48]), .B1(n18), .ZN(N479)
         );
  INR2D1BWP30P140LVT U1214 ( .A1(o_cmd_forward_reg[14]), .B1(n18), .ZN(N1453)
         );
  INR2D1BWP30P140LVT U1215 ( .A1(o_cmd_forward_reg[13]), .B1(n53), .ZN(N1452)
         );
  INR2D1BWP30P140LVT U1216 ( .A1(o_cmd_forward_reg[30]), .B1(n18), .ZN(N1021)
         );
  INR2D1BWP30P140LVT U1217 ( .A1(o_cmd_forward_reg[33]), .B1(n18), .ZN(N912)
         );
  INR2D1BWP30P140LVT U1218 ( .A1(o_cmd_forward_reg[59]), .B1(n53), .ZN(N266)
         );
  INR2D1BWP30P140LVT U1219 ( .A1(o_cmd_forward_reg[47]), .B1(n18), .ZN(N590)
         );
  INR2D1BWP30P140LVT U1220 ( .A1(o_cmd_forward_reg[55]), .B1(n53), .ZN(N374)
         );
  INR2D1BWP30P140LVT U1221 ( .A1(o_cmd_forward_reg[58]), .B1(n18), .ZN(N265)
         );
  INR2D1BWP30P140LVT U1222 ( .A1(o_cmd_forward_reg[32]), .B1(n18), .ZN(N911)
         );
  INR2D1BWP30P140LVT U1223 ( .A1(o_cmd_forward_reg[29]), .B1(n53), .ZN(N1020)
         );
  INR2D1BWP30P140LVT U1224 ( .A1(o_cmd_forward_reg[45]), .B1(n18), .ZN(N588)
         );
  INR2D1BWP30P140LVT U1225 ( .A1(o_data_forward_reg[309]), .B1(n18), .ZN(N462)
         );
  INR2D1BWP30P140LVT U1226 ( .A1(o_data_forward_reg[321]), .B1(n18), .ZN(N474)
         );
  INR2D1BWP30P140LVT U1227 ( .A1(o_data_forward_reg[320]), .B1(n18), .ZN(N473)
         );
  INR2D1BWP30P140LVT U1228 ( .A1(o_data_forward_reg[308]), .B1(n18), .ZN(N461)
         );
  INR2D1BWP30P140LVT U1229 ( .A1(o_data_forward_reg[297]), .B1(n18), .ZN(N583)
         );
  INR2D1BWP30P140LVT U1230 ( .A1(o_data_forward_reg[295]), .B1(n18), .ZN(N581)
         );
  INR2D1BWP30P140LVT U1231 ( .A1(o_data_forward_reg[285]), .B1(n18), .ZN(N571)
         );
  INR2D1BWP30P140LVT U1232 ( .A1(o_data_forward_reg[323]), .B1(n18), .ZN(N476)
         );
  INR2D1BWP30P140LVT U1233 ( .A1(o_data_forward_reg[324]), .B1(n18), .ZN(N477)
         );
  INR2D1BWP30P140LVT U1234 ( .A1(o_data_forward_reg[306]), .B1(n18), .ZN(N459)
         );
  INR2D1BWP30P140LVT U1235 ( .A1(o_data_forward_reg[287]), .B1(n18), .ZN(N573)
         );
  INR2D1BWP30P140LVT U1236 ( .A1(o_data_forward_reg[299]), .B1(n18), .ZN(N585)
         );
  INR2D1BWP30P140LVT U1237 ( .A1(o_data_forward_reg[311]), .B1(n18), .ZN(N464)
         );
  INR2D1BWP30P140LVT U1238 ( .A1(o_data_forward_reg[317]), .B1(n18), .ZN(N470)
         );
  INR2D1BWP30P140LVT U1239 ( .A1(o_data_forward_reg[307]), .B1(n18), .ZN(N460)
         );
  INR2D1BWP30P140LVT U1240 ( .A1(o_data_forward_reg[318]), .B1(n18), .ZN(N471)
         );
  INR2D1BWP30P140LVT U1241 ( .A1(o_data_forward_reg[290]), .B1(n18), .ZN(N576)
         );
  INR2D1BWP30P140LVT U1242 ( .A1(o_data_forward_reg[316]), .B1(n18), .ZN(N469)
         );
  INR2D1BWP30P140LVT U1243 ( .A1(o_data_forward_reg[271]), .B1(n18), .ZN(N690)
         );
  INR2D1BWP30P140LVT U1244 ( .A1(o_data_forward_reg[269]), .B1(n18), .ZN(N688)
         );
  INR2D1BWP30P140LVT U1245 ( .A1(o_data_forward_reg[268]), .B1(n18), .ZN(N687)
         );
  INR2D1BWP30P140LVT U1246 ( .A1(o_data_forward_reg[265]), .B1(n18), .ZN(N684)
         );
  INR2D1BWP30P140LVT U1247 ( .A1(o_data_forward_reg[274]), .B1(n18), .ZN(N693)
         );
  INR2D1BWP30P140LVT U1248 ( .A1(o_data_forward_reg[314]), .B1(n18), .ZN(N467)
         );
  INR2D1BWP30P140LVT U1249 ( .A1(o_data_forward_reg[264]), .B1(n18), .ZN(N683)
         );
  INR2D1BWP30P140LVT U1250 ( .A1(o_data_forward_reg[262]), .B1(n18), .ZN(N681)
         );
  INR2D1BWP30P140LVT U1251 ( .A1(o_data_forward_reg[260]), .B1(n18), .ZN(N679)
         );
  INR2D1BWP30P140LVT U1252 ( .A1(o_data_forward_reg[257]), .B1(n18), .ZN(N676)
         );
  INR2D1BWP30P140LVT U1253 ( .A1(o_data_forward_reg[255]), .B1(n18), .ZN(N674)
         );
  INR2D1BWP30P140LVT U1254 ( .A1(o_data_forward_reg[253]), .B1(n18), .ZN(N672)
         );
  INR2D1BWP30P140LVT U1255 ( .A1(o_data_forward_reg[251]), .B1(n18), .ZN(N670)
         );
  INR2D1BWP30P140LVT U1256 ( .A1(o_data_forward_reg[293]), .B1(n18), .ZN(N579)
         );
  INR2D1BWP30P140LVT U1257 ( .A1(o_data_forward_reg[291]), .B1(n18), .ZN(N577)
         );
  INR2D1BWP30P140LVT U1258 ( .A1(o_data_forward_reg[231]), .B1(n18), .ZN(N783)
         );
  INR2D1BWP30P140LVT U1259 ( .A1(o_data_forward_reg[230]), .B1(n18), .ZN(N782)
         );
  INR2D1BWP30P140LVT U1260 ( .A1(o_data_forward_reg[227]), .B1(n18), .ZN(N779)
         );
  INR2D1BWP30P140LVT U1261 ( .A1(o_data_forward_reg[225]), .B1(n18), .ZN(N777)
         );
  INR2D1BWP30P140LVT U1262 ( .A1(o_data_forward_reg[280]), .B1(n18), .ZN(N566)
         );
  INR2D1BWP30P140LVT U1263 ( .A1(o_data_forward_reg[312]), .B1(n18), .ZN(N465)
         );
  INR2D1BWP30P140LVT U1264 ( .A1(o_data_forward_reg[313]), .B1(n18), .ZN(N466)
         );
  INR2D1BWP30P140LVT U1265 ( .A1(o_data_forward_reg[278]), .B1(n18), .ZN(N564)
         );
  INR2D1BWP30P140LVT U1266 ( .A1(o_data_forward_reg[315]), .B1(n18), .ZN(N468)
         );
  INR2D1BWP30P140LVT U1267 ( .A1(o_data_forward_reg[276]), .B1(n18), .ZN(N562)
         );
  INR2D1BWP30P140LVT U1268 ( .A1(o_data_forward_reg[310]), .B1(n18), .ZN(N463)
         );
  INR2D1BWP30P140LVT U1269 ( .A1(o_data_forward_reg[242]), .B1(n18), .ZN(N794)
         );
  INR2D1BWP30P140LVT U1270 ( .A1(o_data_forward_reg[252]), .B1(n18), .ZN(N671)
         );
  INR2D1BWP30P140LVT U1271 ( .A1(o_data_forward_reg[256]), .B1(n18), .ZN(N675)
         );
  INR2D1BWP30P140LVT U1272 ( .A1(o_data_forward_reg[250]), .B1(n18), .ZN(N669)
         );
  INR2D1BWP30P140LVT U1273 ( .A1(o_data_forward_reg[258]), .B1(n18), .ZN(N677)
         );
  INR2D1BWP30P140LVT U1274 ( .A1(o_data_forward_reg[237]), .B1(n18), .ZN(N789)
         );
  INR2D1BWP30P140LVT U1275 ( .A1(o_data_forward_reg[259]), .B1(n18), .ZN(N678)
         );
  INR2D1BWP30P140LVT U1276 ( .A1(o_data_forward_reg[275]), .B1(n18), .ZN(N561)
         );
  INR2D1BWP30P140LVT U1277 ( .A1(o_data_forward_reg[322]), .B1(n18), .ZN(N475)
         );
  INR2D1BWP30P140LVT U1278 ( .A1(o_data_forward_reg[261]), .B1(n18), .ZN(N680)
         );
  INR2D1BWP30P140LVT U1279 ( .A1(o_data_forward_reg[263]), .B1(n18), .ZN(N682)
         );
  INR2D1BWP30P140LVT U1280 ( .A1(o_data_forward_reg[266]), .B1(n18), .ZN(N685)
         );
  INR2D1BWP30P140LVT U1281 ( .A1(o_data_forward_reg[267]), .B1(n18), .ZN(N686)
         );
  INR2D1BWP30P140LVT U1282 ( .A1(o_data_forward_reg[245]), .B1(n18), .ZN(N797)
         );
  INR2D1BWP30P140LVT U1283 ( .A1(o_data_forward_reg[244]), .B1(n18), .ZN(N796)
         );
  INR2D1BWP30P140LVT U1284 ( .A1(o_data_forward_reg[243]), .B1(n18), .ZN(N795)
         );
  INR2D1BWP30P140LVT U1285 ( .A1(o_data_forward_reg[226]), .B1(n18), .ZN(N778)
         );
  INR2D1BWP30P140LVT U1286 ( .A1(o_data_forward_reg[241]), .B1(n18), .ZN(N793)
         );
  INR2D1BWP30P140LVT U1287 ( .A1(o_data_forward_reg[240]), .B1(n18), .ZN(N792)
         );
  INR2D1BWP30P140LVT U1288 ( .A1(o_data_forward_reg[239]), .B1(n18), .ZN(N791)
         );
  INR2D1BWP30P140LVT U1289 ( .A1(o_data_forward_reg[238]), .B1(n18), .ZN(N790)
         );
  INR2D1BWP30P140LVT U1290 ( .A1(o_data_forward_reg[279]), .B1(n18), .ZN(N565)
         );
  INR2D1BWP30P140LVT U1291 ( .A1(o_data_forward_reg[236]), .B1(n18), .ZN(N788)
         );
  INR2D1BWP30P140LVT U1292 ( .A1(o_data_forward_reg[235]), .B1(n18), .ZN(N787)
         );
  INR2D1BWP30P140LVT U1293 ( .A1(o_data_forward_reg[234]), .B1(n18), .ZN(N786)
         );
  INR2D1BWP30P140LVT U1294 ( .A1(o_data_forward_reg[233]), .B1(n18), .ZN(N785)
         );
  INR2D1BWP30P140LVT U1295 ( .A1(o_data_forward_reg[232]), .B1(n18), .ZN(N784)
         );
  INR2D1BWP30P140LVT U1296 ( .A1(o_data_forward_reg[270]), .B1(n18), .ZN(N689)
         );
  INR2D1BWP30P140LVT U1297 ( .A1(o_data_forward_reg[272]), .B1(n18), .ZN(N691)
         );
  INR2D1BWP30P140LVT U1298 ( .A1(o_data_forward_reg[229]), .B1(n18), .ZN(N781)
         );
  INR2D1BWP30P140LVT U1299 ( .A1(o_data_forward_reg[228]), .B1(n18), .ZN(N780)
         );
  INR2D1BWP30P140LVT U1300 ( .A1(o_data_forward_reg[273]), .B1(n18), .ZN(N692)
         );
  INR2D1BWP30P140LVT U1301 ( .A1(o_data_forward_reg[294]), .B1(n18), .ZN(N580)
         );
  INR2D1BWP30P140LVT U1302 ( .A1(o_data_forward_reg[254]), .B1(n18), .ZN(N673)
         );
  INR2D1BWP30P140LVT U1303 ( .A1(o_data_forward_reg[292]), .B1(n18), .ZN(N578)
         );
  INR2D1BWP30P140LVT U1304 ( .A1(o_data_forward_reg[298]), .B1(n18), .ZN(N584)
         );
  INR2D1BWP30P140LVT U1305 ( .A1(o_data_forward_reg[288]), .B1(n18), .ZN(N574)
         );
  INR2D1BWP30P140LVT U1306 ( .A1(o_data_forward_reg[296]), .B1(n18), .ZN(N582)
         );
  INR2D1BWP30P140LVT U1307 ( .A1(o_data_forward_reg[319]), .B1(n18), .ZN(N472)
         );
  INR2D1BWP30P140LVT U1308 ( .A1(o_data_forward_reg[284]), .B1(n18), .ZN(N570)
         );
  INR2D1BWP30P140LVT U1309 ( .A1(o_data_forward_reg[283]), .B1(n18), .ZN(N569)
         );
  INR2D1BWP30P140LVT U1310 ( .A1(o_data_forward_reg[286]), .B1(n18), .ZN(N572)
         );
  INR2D1BWP30P140LVT U1311 ( .A1(o_data_forward_reg[289]), .B1(n18), .ZN(N575)
         );
  INR2D1BWP30P140LVT U1312 ( .A1(o_data_forward_reg[281]), .B1(n18), .ZN(N567)
         );
  INR2D1BWP30P140LVT U1313 ( .A1(o_cmd_forward_reg[54]), .B1(n18), .ZN(N373)
         );
  INR2D1BWP30P140LVT U1314 ( .A1(o_data_forward_reg[220]), .B1(n53), .ZN(N905)
         );
  INR2D1BWP30P140LVT U1315 ( .A1(o_data_forward_reg[218]), .B1(n53), .ZN(N903)
         );
  INR2D1BWP30P140LVT U1316 ( .A1(o_data_forward_reg[223]), .B1(n53), .ZN(N908)
         );
  INR2D1BWP30P140LVT U1317 ( .A1(o_data_forward_reg[216]), .B1(n53), .ZN(N901)
         );
  INR2D1BWP30P140LVT U1318 ( .A1(o_data_forward_reg[159]), .B1(n53), .ZN(N1110) );
  INR2D1BWP30P140LVT U1319 ( .A1(o_data_forward_reg[162]), .B1(n53), .ZN(N1113) );
  INR2D1BWP30P140LVT U1320 ( .A1(o_data_forward_reg[156]), .B1(n53), .ZN(N1107) );
  INR2D1BWP30P140LVT U1321 ( .A1(o_data_forward_reg[165]), .B1(n53), .ZN(N1116) );
  INR2D1BWP30P140LVT U1322 ( .A1(o_data_forward_reg[213]), .B1(n53), .ZN(N898)
         );
  INR2D1BWP30P140LVT U1323 ( .A1(o_data_forward_reg[168]), .B1(n53), .ZN(N1119) );
  INR2D1BWP30P140LVT U1324 ( .A1(o_data_forward_reg[215]), .B1(n53), .ZN(N900)
         );
  INR2D1BWP30P140LVT U1325 ( .A1(o_data_forward_reg[171]), .B1(n53), .ZN(N1122) );
  INR2D1BWP30P140LVT U1326 ( .A1(o_data_forward_reg[190]), .B1(n53), .ZN(N1008) );
  INR2D1BWP30P140LVT U1327 ( .A1(o_data_forward_reg[212]), .B1(n53), .ZN(N897)
         );
  INR2D1BWP30P140LVT U1328 ( .A1(o_data_forward_reg[211]), .B1(n53), .ZN(N896)
         );
  INR2D1BWP30P140LVT U1329 ( .A1(o_data_forward_reg[210]), .B1(n53), .ZN(N895)
         );
  INR2D1BWP30P140LVT U1330 ( .A1(o_data_forward_reg[176]), .B1(n53), .ZN(N994)
         );
  INR2D1BWP30P140LVT U1331 ( .A1(o_data_forward_reg[195]), .B1(n53), .ZN(N1013) );
  INR2D1BWP30P140LVT U1332 ( .A1(o_data_forward_reg[152]), .B1(n53), .ZN(N1103) );
  INR2D1BWP30P140LVT U1333 ( .A1(o_data_forward_reg[282]), .B1(n53), .ZN(N568)
         );
  INR2D1BWP30P140LVT U1334 ( .A1(o_data_forward_reg[181]), .B1(n53), .ZN(N999)
         );
  INR2D1BWP30P140LVT U1335 ( .A1(o_data_forward_reg[182]), .B1(n53), .ZN(N1000) );
  INR2D1BWP30P140LVT U1336 ( .A1(o_data_forward_reg[219]), .B1(n53), .ZN(N904)
         );
  INR2D1BWP30P140LVT U1337 ( .A1(o_data_forward_reg[184]), .B1(n53), .ZN(N1002) );
  INR2D1BWP30P140LVT U1338 ( .A1(o_data_forward_reg[185]), .B1(n53), .ZN(N1003) );
  INR2D1BWP30P140LVT U1339 ( .A1(o_data_forward_reg[209]), .B1(n53), .ZN(N894)
         );
  INR2D1BWP30P140LVT U1340 ( .A1(o_data_forward_reg[208]), .B1(n53), .ZN(N893)
         );
  INR2D1BWP30P140LVT U1341 ( .A1(o_data_forward_reg[198]), .B1(n53), .ZN(N1016) );
  INR2D1BWP30P140LVT U1342 ( .A1(o_data_forward_reg[217]), .B1(n53), .ZN(N902)
         );
  INR2D1BWP30P140LVT U1343 ( .A1(o_data_forward_reg[197]), .B1(n53), .ZN(N1015) );
  INR2D1BWP30P140LVT U1344 ( .A1(o_data_forward_reg[277]), .B1(n53), .ZN(N563)
         );
  INR2D1BWP30P140LVT U1345 ( .A1(o_data_forward_reg[214]), .B1(n53), .ZN(N899)
         );
  INR2D1BWP30P140LVT U1346 ( .A1(o_cmd_forward_reg[26]), .B1(n18), .ZN(N1129)
         );
  INR2D1BWP30P140LVT U1347 ( .A1(o_cmd_forward_reg[43]), .B1(n18), .ZN(N698)
         );
  INR2D1BWP30P140LVT U1348 ( .A1(o_cmd_forward_reg[22]), .B1(n18), .ZN(N1237)
         );
  INR2D1BWP30P140LVT U1349 ( .A1(o_cmd_forward_reg[51]), .B1(n18), .ZN(N482)
         );
  INR2D1BWP30P140LVT U1350 ( .A1(o_cmd_forward_reg[39]), .B1(n18), .ZN(N806)
         );
  INR2D1BWP30P140LVT U1351 ( .A1(i_cmd[2]), .B1(n18), .ZN(N157) );
  INR2D1BWP30P140LVT U1352 ( .A1(i_cmd[3]), .B1(n18), .ZN(N158) );
  INR2D1BWP30P140LVT U1353 ( .A1(i_cmd[1]), .B1(n18), .ZN(N156) );
  CKAN2D1BWP30P140LVT U1354 ( .A1(n230), .A2(o_data_forward_reg[313]), .Z(n54)
         );
  CKAN2D1BWP30P140LVT U1355 ( .A1(n230), .A2(o_data_forward_reg[314]), .Z(n55)
         );
  CKAN2D1BWP30P140LVT U1356 ( .A1(n230), .A2(o_data_forward_reg[315]), .Z(n56)
         );
  CKAN2D1BWP30P140LVT U1357 ( .A1(n230), .A2(o_data_forward_reg[316]), .Z(n57)
         );
  CKAN2D1BWP30P140LVT U1358 ( .A1(n230), .A2(o_data_forward_reg[317]), .Z(n58)
         );
  CKAN2D1BWP30P140LVT U1359 ( .A1(n230), .A2(o_data_forward_reg[318]), .Z(n59)
         );
  CKAN2D1BWP30P140LVT U1360 ( .A1(n230), .A2(o_data_forward_reg[319]), .Z(n60)
         );
  CKAN2D1BWP30P140LVT U1361 ( .A1(n230), .A2(o_data_forward_reg[320]), .Z(n61)
         );
  CKAN2D1BWP30P140LVT U1362 ( .A1(n230), .A2(o_data_forward_reg[321]), .Z(n62)
         );
  CKAN2D1BWP30P140LVT U1363 ( .A1(n230), .A2(o_data_forward_reg[322]), .Z(n63)
         );
  CKAN2D1BWP30P140LVT U1364 ( .A1(n230), .A2(o_data_forward_reg[323]), .Z(n64)
         );
  CKAN2D1BWP30P140LVT U1365 ( .A1(n230), .A2(o_data_forward_reg[324]), .Z(n65)
         );
  CKAN2D1BWP30P140LVT U1366 ( .A1(n231), .A2(o_data_forward_reg[238]), .Z(n66)
         );
  CKAN2D1BWP30P140LVT U1367 ( .A1(n231), .A2(o_data_forward_reg[239]), .Z(n67)
         );
  CKAN2D1BWP30P140LVT U1368 ( .A1(n231), .A2(o_data_forward_reg[240]), .Z(n68)
         );
  CKAN2D1BWP30P140LVT U1369 ( .A1(n231), .A2(o_data_forward_reg[241]), .Z(n69)
         );
  CKAN2D1BWP30P140LVT U1370 ( .A1(n231), .A2(o_data_forward_reg[242]), .Z(n70)
         );
  CKAN2D1BWP30P140LVT U1371 ( .A1(n231), .A2(o_data_forward_reg[243]), .Z(n71)
         );
  CKAN2D1BWP30P140LVT U1372 ( .A1(n231), .A2(o_data_forward_reg[244]), .Z(n72)
         );
  CKAN2D1BWP30P140LVT U1373 ( .A1(n231), .A2(o_data_forward_reg[245]), .Z(n73)
         );
  CKAN2D1BWP30P140LVT U1374 ( .A1(n231), .A2(o_data_forward_reg[246]), .Z(n74)
         );
  CKAN2D1BWP30P140LVT U1375 ( .A1(n231), .A2(o_data_forward_reg[247]), .Z(n75)
         );
  CKAN2D1BWP30P140LVT U1376 ( .A1(n231), .A2(o_data_forward_reg[248]), .Z(n76)
         );
  CKAN2D1BWP30P140LVT U1377 ( .A1(n231), .A2(o_data_forward_reg[249]), .Z(n77)
         );
  CKAN2D1BWP30P140LVT U1378 ( .A1(n232), .A2(o_data_forward_reg[138]), .Z(n78)
         );
  CKAN2D1BWP30P140LVT U1379 ( .A1(n232), .A2(o_data_forward_reg[139]), .Z(n79)
         );
  CKAN2D1BWP30P140LVT U1380 ( .A1(n232), .A2(o_data_forward_reg[140]), .Z(n80)
         );
  CKAN2D1BWP30P140LVT U1381 ( .A1(n232), .A2(o_data_forward_reg[141]), .Z(n81)
         );
  CKAN2D1BWP30P140LVT U1382 ( .A1(n232), .A2(o_data_forward_reg[142]), .Z(n82)
         );
  CKAN2D1BWP30P140LVT U1383 ( .A1(n232), .A2(o_data_forward_reg[143]), .Z(n83)
         );
  CKAN2D1BWP30P140LVT U1384 ( .A1(n232), .A2(o_data_forward_reg[144]), .Z(n84)
         );
  CKAN2D1BWP30P140LVT U1385 ( .A1(n232), .A2(o_data_forward_reg[145]), .Z(n85)
         );
  CKAN2D1BWP30P140LVT U1386 ( .A1(n232), .A2(o_data_forward_reg[146]), .Z(n86)
         );
  CKAN2D1BWP30P140LVT U1387 ( .A1(n232), .A2(o_data_forward_reg[147]), .Z(n87)
         );
  CKAN2D1BWP30P140LVT U1388 ( .A1(n232), .A2(o_data_forward_reg[148]), .Z(n88)
         );
  CKAN2D1BWP30P140LVT U1389 ( .A1(n232), .A2(o_data_forward_reg[149]), .Z(n89)
         );
  CKAN2D1BWP30P140LVT U1390 ( .A1(n233), .A2(o_data_forward_reg[88]), .Z(n90)
         );
  CKAN2D1BWP30P140LVT U1391 ( .A1(n233), .A2(o_data_forward_reg[89]), .Z(n91)
         );
  CKAN2D1BWP30P140LVT U1392 ( .A1(n233), .A2(o_data_forward_reg[90]), .Z(n92)
         );
  CKAN2D1BWP30P140LVT U1393 ( .A1(n233), .A2(o_data_forward_reg[91]), .Z(n93)
         );
  CKAN2D1BWP30P140LVT U1394 ( .A1(n233), .A2(o_data_forward_reg[92]), .Z(n94)
         );
  CKAN2D1BWP30P140LVT U1395 ( .A1(n233), .A2(o_data_forward_reg[93]), .Z(n95)
         );
  CKAN2D1BWP30P140LVT U1396 ( .A1(n233), .A2(o_data_forward_reg[94]), .Z(n96)
         );
  CKAN2D1BWP30P140LVT U1397 ( .A1(n233), .A2(o_data_forward_reg[95]), .Z(n97)
         );
  CKAN2D1BWP30P140LVT U1398 ( .A1(n233), .A2(o_data_forward_reg[96]), .Z(n98)
         );
  CKAN2D1BWP30P140LVT U1399 ( .A1(n233), .A2(o_data_forward_reg[97]), .Z(n99)
         );
  CKAN2D1BWP30P140LVT U1400 ( .A1(n233), .A2(o_data_forward_reg[98]), .Z(n100)
         );
  CKAN2D1BWP30P140LVT U1401 ( .A1(n233), .A2(o_data_forward_reg[99]), .Z(n101)
         );
  CKAN2D1BWP30P140LVT U1402 ( .A1(n234), .A2(o_data_forward_reg[13]), .Z(n102)
         );
  CKAN2D1BWP30P140LVT U1403 ( .A1(n234), .A2(o_data_forward_reg[14]), .Z(n103)
         );
  CKAN2D1BWP30P140LVT U1404 ( .A1(n234), .A2(o_data_forward_reg[15]), .Z(n104)
         );
  CKAN2D1BWP30P140LVT U1405 ( .A1(n234), .A2(o_data_forward_reg[16]), .Z(n105)
         );
  CKAN2D1BWP30P140LVT U1406 ( .A1(n234), .A2(o_data_forward_reg[17]), .Z(n106)
         );
  CKAN2D1BWP30P140LVT U1407 ( .A1(n234), .A2(o_data_forward_reg[18]), .Z(n107)
         );
  CKAN2D1BWP30P140LVT U1408 ( .A1(n234), .A2(o_data_forward_reg[19]), .Z(n108)
         );
  CKAN2D1BWP30P140LVT U1409 ( .A1(n234), .A2(o_data_forward_reg[20]), .Z(n109)
         );
  CKAN2D1BWP30P140LVT U1410 ( .A1(n234), .A2(o_data_forward_reg[21]), .Z(n110)
         );
  CKAN2D1BWP30P140LVT U1411 ( .A1(n234), .A2(o_data_forward_reg[22]), .Z(n111)
         );
  CKAN2D1BWP30P140LVT U1412 ( .A1(n234), .A2(o_data_forward_reg[23]), .Z(n112)
         );
  CKAN2D1BWP30P140LVT U1413 ( .A1(n234), .A2(o_data_forward_reg[24]), .Z(n113)
         );
  CKAN2D1BWP30P140LVT U1414 ( .A1(n230), .A2(o_data_forward_reg[300]), .Z(n114) );
  CKAN2D1BWP30P140LVT U1415 ( .A1(n230), .A2(o_data_forward_reg[301]), .Z(n115) );
  CKAN2D1BWP30P140LVT U1416 ( .A1(n230), .A2(o_data_forward_reg[302]), .Z(n116) );
  CKAN2D1BWP30P140LVT U1417 ( .A1(n230), .A2(o_data_forward_reg[303]), .Z(n117) );
  CKAN2D1BWP30P140LVT U1418 ( .A1(n230), .A2(o_data_forward_reg[304]), .Z(n118) );
  CKAN2D1BWP30P140LVT U1419 ( .A1(n230), .A2(o_data_forward_reg[305]), .Z(n119) );
  CKAN2D1BWP30P140LVT U1420 ( .A1(n230), .A2(o_data_forward_reg[306]), .Z(n120) );
  CKAN2D1BWP30P140LVT U1421 ( .A1(n230), .A2(o_data_forward_reg[307]), .Z(n121) );
  CKAN2D1BWP30P140LVT U1422 ( .A1(n230), .A2(o_data_forward_reg[308]), .Z(n122) );
  CKAN2D1BWP30P140LVT U1423 ( .A1(n230), .A2(o_data_forward_reg[309]), .Z(n123) );
  CKAN2D1BWP30P140LVT U1424 ( .A1(n230), .A2(o_data_forward_reg[310]), .Z(n124) );
  CKAN2D1BWP30P140LVT U1425 ( .A1(n230), .A2(o_data_forward_reg[311]), .Z(n125) );
  CKAN2D1BWP30P140LVT U1426 ( .A1(n230), .A2(o_data_forward_reg[312]), .Z(n126) );
  CKAN2D1BWP30P140LVT U1427 ( .A1(n231), .A2(o_data_forward_reg[225]), .Z(n127) );
  CKAN2D1BWP30P140LVT U1428 ( .A1(n231), .A2(o_data_forward_reg[226]), .Z(n128) );
  CKAN2D1BWP30P140LVT U1429 ( .A1(n231), .A2(o_data_forward_reg[227]), .Z(n129) );
  CKAN2D1BWP30P140LVT U1430 ( .A1(n231), .A2(o_data_forward_reg[228]), .Z(n130) );
  CKAN2D1BWP30P140LVT U1431 ( .A1(n231), .A2(o_data_forward_reg[229]), .Z(n131) );
  CKAN2D1BWP30P140LVT U1432 ( .A1(n231), .A2(o_data_forward_reg[230]), .Z(n132) );
  CKAN2D1BWP30P140LVT U1433 ( .A1(n231), .A2(o_data_forward_reg[231]), .Z(n133) );
  CKAN2D1BWP30P140LVT U1434 ( .A1(n231), .A2(o_data_forward_reg[232]), .Z(n134) );
  CKAN2D1BWP30P140LVT U1435 ( .A1(n231), .A2(o_data_forward_reg[233]), .Z(n135) );
  CKAN2D1BWP30P140LVT U1436 ( .A1(n231), .A2(o_data_forward_reg[234]), .Z(n136) );
  CKAN2D1BWP30P140LVT U1437 ( .A1(n231), .A2(o_data_forward_reg[235]), .Z(n137) );
  CKAN2D1BWP30P140LVT U1438 ( .A1(n231), .A2(o_data_forward_reg[236]), .Z(n138) );
  CKAN2D1BWP30P140LVT U1439 ( .A1(n231), .A2(o_data_forward_reg[237]), .Z(n139) );
  CKAN2D1BWP30P140LVT U1440 ( .A1(n232), .A2(o_data_forward_reg[125]), .Z(n140) );
  CKAN2D1BWP30P140LVT U1441 ( .A1(n232), .A2(o_data_forward_reg[126]), .Z(n141) );
  CKAN2D1BWP30P140LVT U1442 ( .A1(n232), .A2(o_data_forward_reg[127]), .Z(n142) );
  CKAN2D1BWP30P140LVT U1443 ( .A1(n232), .A2(o_data_forward_reg[128]), .Z(n143) );
  CKAN2D1BWP30P140LVT U1444 ( .A1(n232), .A2(o_data_forward_reg[129]), .Z(n144) );
  CKAN2D1BWP30P140LVT U1445 ( .A1(n232), .A2(o_data_forward_reg[130]), .Z(n145) );
  CKAN2D1BWP30P140LVT U1446 ( .A1(n232), .A2(o_data_forward_reg[131]), .Z(n146) );
  CKAN2D1BWP30P140LVT U1447 ( .A1(n232), .A2(o_data_forward_reg[132]), .Z(n147) );
  CKAN2D1BWP30P140LVT U1448 ( .A1(n232), .A2(o_data_forward_reg[133]), .Z(n148) );
  CKAN2D1BWP30P140LVT U1449 ( .A1(n232), .A2(o_data_forward_reg[134]), .Z(n149) );
  CKAN2D1BWP30P140LVT U1450 ( .A1(n232), .A2(o_data_forward_reg[135]), .Z(n150) );
  CKAN2D1BWP30P140LVT U1451 ( .A1(n232), .A2(o_data_forward_reg[136]), .Z(n151) );
  CKAN2D1BWP30P140LVT U1452 ( .A1(n232), .A2(o_data_forward_reg[137]), .Z(n152) );
  CKAN2D1BWP30P140LVT U1453 ( .A1(n233), .A2(o_data_forward_reg[75]), .Z(n153)
         );
  CKAN2D1BWP30P140LVT U1454 ( .A1(n233), .A2(o_data_forward_reg[76]), .Z(n154)
         );
  CKAN2D1BWP30P140LVT U1455 ( .A1(n233), .A2(o_data_forward_reg[77]), .Z(n155)
         );
  CKAN2D1BWP30P140LVT U1456 ( .A1(n233), .A2(o_data_forward_reg[78]), .Z(n156)
         );
  CKAN2D1BWP30P140LVT U1457 ( .A1(n233), .A2(o_data_forward_reg[79]), .Z(n157)
         );
  CKAN2D1BWP30P140LVT U1458 ( .A1(n233), .A2(o_data_forward_reg[80]), .Z(n158)
         );
  CKAN2D1BWP30P140LVT U1459 ( .A1(n233), .A2(o_data_forward_reg[81]), .Z(n159)
         );
  CKAN2D1BWP30P140LVT U1460 ( .A1(n233), .A2(o_data_forward_reg[82]), .Z(n160)
         );
  CKAN2D1BWP30P140LVT U1461 ( .A1(n233), .A2(o_data_forward_reg[83]), .Z(n161)
         );
  CKAN2D1BWP30P140LVT U1462 ( .A1(n233), .A2(o_data_forward_reg[84]), .Z(n162)
         );
  CKAN2D1BWP30P140LVT U1463 ( .A1(n233), .A2(o_data_forward_reg[85]), .Z(n163)
         );
  CKAN2D1BWP30P140LVT U1464 ( .A1(n233), .A2(o_data_forward_reg[86]), .Z(n164)
         );
  CKAN2D1BWP30P140LVT U1465 ( .A1(n233), .A2(o_data_forward_reg[87]), .Z(n165)
         );
  CKAN2D1BWP30P140LVT U1466 ( .A1(n229), .A2(i_data_bus[13]), .Z(n166) );
  CKAN2D1BWP30P140LVT U1467 ( .A1(n229), .A2(i_data_bus[14]), .Z(n167) );
  CKAN2D1BWP30P140LVT U1468 ( .A1(n229), .A2(i_data_bus[15]), .Z(n168) );
  CKAN2D1BWP30P140LVT U1469 ( .A1(n229), .A2(i_data_bus[16]), .Z(n169) );
  CKAN2D1BWP30P140LVT U1470 ( .A1(n229), .A2(i_data_bus[17]), .Z(n170) );
  CKAN2D1BWP30P140LVT U1471 ( .A1(n229), .A2(i_data_bus[18]), .Z(n171) );
  CKAN2D1BWP30P140LVT U1472 ( .A1(n229), .A2(i_data_bus[19]), .Z(n172) );
  CKAN2D1BWP30P140LVT U1473 ( .A1(n229), .A2(i_data_bus[20]), .Z(n173) );
  CKAN2D1BWP30P140LVT U1474 ( .A1(n229), .A2(i_data_bus[21]), .Z(n174) );
  CKAN2D1BWP30P140LVT U1475 ( .A1(n229), .A2(i_data_bus[22]), .Z(n175) );
  CKAN2D1BWP30P140LVT U1476 ( .A1(n229), .A2(i_data_bus[23]), .Z(n176) );
  CKAN2D1BWP30P140LVT U1477 ( .A1(n229), .A2(i_data_bus[24]), .Z(n177) );
  CKAN2D1BWP30P140LVT U1478 ( .A1(n234), .A2(o_data_forward_reg[0]), .Z(n203)
         );
  CKAN2D1BWP30P140LVT U1479 ( .A1(n234), .A2(o_data_forward_reg[1]), .Z(n204)
         );
  CKAN2D1BWP30P140LVT U1480 ( .A1(n234), .A2(o_data_forward_reg[2]), .Z(n205)
         );
  CKAN2D1BWP30P140LVT U1481 ( .A1(n234), .A2(o_data_forward_reg[3]), .Z(n206)
         );
  CKAN2D1BWP30P140LVT U1482 ( .A1(n234), .A2(o_data_forward_reg[4]), .Z(n207)
         );
  CKAN2D1BWP30P140LVT U1483 ( .A1(n234), .A2(o_data_forward_reg[5]), .Z(n208)
         );
  CKAN2D1BWP30P140LVT U1484 ( .A1(n234), .A2(o_data_forward_reg[6]), .Z(n209)
         );
  CKAN2D1BWP30P140LVT U1485 ( .A1(n234), .A2(o_data_forward_reg[7]), .Z(n210)
         );
  CKAN2D1BWP30P140LVT U1486 ( .A1(n234), .A2(o_data_forward_reg[8]), .Z(n211)
         );
  CKAN2D1BWP30P140LVT U1487 ( .A1(n234), .A2(o_data_forward_reg[9]), .Z(n212)
         );
  CKAN2D1BWP30P140LVT U1488 ( .A1(n234), .A2(o_data_forward_reg[10]), .Z(n213)
         );
  CKAN2D1BWP30P140LVT U1489 ( .A1(n234), .A2(o_data_forward_reg[11]), .Z(n214)
         );
  CKAN2D1BWP30P140LVT U1490 ( .A1(n234), .A2(o_data_forward_reg[12]), .Z(n215)
         );
  CKAN2D1BWP30P140LVT U1491 ( .A1(n229), .A2(i_data_bus[0]), .Z(n216) );
  CKAN2D1BWP30P140LVT U1492 ( .A1(n229), .A2(i_data_bus[1]), .Z(n217) );
  CKAN2D1BWP30P140LVT U1493 ( .A1(n229), .A2(i_data_bus[2]), .Z(n218) );
  CKAN2D1BWP30P140LVT U1494 ( .A1(n229), .A2(i_data_bus[3]), .Z(n219) );
  CKAN2D1BWP30P140LVT U1495 ( .A1(n229), .A2(i_data_bus[4]), .Z(n220) );
  CKAN2D1BWP30P140LVT U1496 ( .A1(n229), .A2(i_data_bus[5]), .Z(n221) );
  CKAN2D1BWP30P140LVT U1497 ( .A1(n229), .A2(i_data_bus[6]), .Z(n222) );
  CKAN2D1BWP30P140LVT U1498 ( .A1(n229), .A2(i_data_bus[7]), .Z(n223) );
  CKAN2D1BWP30P140LVT U1499 ( .A1(n229), .A2(i_data_bus[8]), .Z(n224) );
  CKAN2D1BWP30P140LVT U1500 ( .A1(n229), .A2(i_data_bus[9]), .Z(n225) );
  CKAN2D1BWP30P140LVT U1501 ( .A1(n229), .A2(i_data_bus[10]), .Z(n226) );
  CKAN2D1BWP30P140LVT U1502 ( .A1(n229), .A2(i_data_bus[11]), .Z(n227) );
  CKAN2D1BWP30P140LVT U1503 ( .A1(n229), .A2(i_data_bus[12]), .Z(n228) );
  CKAN2D1BWP30P140LVT U1504 ( .A1(n235), .A2(o_data_forward_reg[350]), .Z(N212) );
  CKAN2D1BWP30P140LVT U1505 ( .A1(n235), .A2(o_data_forward_reg[351]), .Z(N213) );
  CKAN2D1BWP30P140LVT U1506 ( .A1(n235), .A2(o_data_forward_reg[352]), .Z(N214) );
  CKAN2D1BWP30P140LVT U1507 ( .A1(n235), .A2(o_data_forward_reg[353]), .Z(N215) );
  CKAN2D1BWP30P140LVT U1508 ( .A1(n235), .A2(o_data_forward_reg[354]), .Z(N216) );
  CKAN2D1BWP30P140LVT U1509 ( .A1(n235), .A2(o_data_forward_reg[355]), .Z(N217) );
  CKAN2D1BWP30P140LVT U1510 ( .A1(n235), .A2(o_data_forward_reg[356]), .Z(N218) );
  CKAN2D1BWP30P140LVT U1511 ( .A1(n235), .A2(o_data_forward_reg[357]), .Z(N219) );
  CKAN2D1BWP30P140LVT U1512 ( .A1(n235), .A2(o_data_forward_reg[358]), .Z(N220) );
  CKAN2D1BWP30P140LVT U1513 ( .A1(n235), .A2(o_data_forward_reg[359]), .Z(N221) );
  CKAN2D1BWP30P140LVT U1514 ( .A1(n235), .A2(o_data_forward_reg[360]), .Z(N222) );
  CKAN2D1BWP30P140LVT U1515 ( .A1(n235), .A2(o_data_forward_reg[361]), .Z(N223) );
  CKAN2D1BWP30P140LVT U1516 ( .A1(n235), .A2(o_data_forward_reg[362]), .Z(N224) );
  CKAN2D1BWP30P140LVT U1517 ( .A1(n22), .A2(o_data_forward_reg[363]), .Z(N225)
         );
  CKAN2D1BWP30P140LVT U1518 ( .A1(n22), .A2(o_data_forward_reg[364]), .Z(N226)
         );
  CKAN2D1BWP30P140LVT U1519 ( .A1(n22), .A2(o_data_forward_reg[365]), .Z(N227)
         );
  CKAN2D1BWP30P140LVT U1520 ( .A1(n22), .A2(o_data_forward_reg[366]), .Z(N228)
         );
  CKAN2D1BWP30P140LVT U1521 ( .A1(n22), .A2(o_data_forward_reg[367]), .Z(N229)
         );
  CKAN2D1BWP30P140LVT U1522 ( .A1(n22), .A2(o_data_forward_reg[368]), .Z(N230)
         );
  CKAN2D1BWP30P140LVT U1523 ( .A1(n22), .A2(o_data_forward_reg[369]), .Z(N231)
         );
  CKAN2D1BWP30P140LVT U1524 ( .A1(n22), .A2(o_data_forward_reg[370]), .Z(N232)
         );
  CKAN2D1BWP30P140LVT U1525 ( .A1(n22), .A2(o_data_forward_reg[371]), .Z(N233)
         );
  CKAN2D1BWP30P140LVT U1526 ( .A1(n22), .A2(o_data_forward_reg[372]), .Z(N234)
         );
  CKAN2D1BWP30P140LVT U1527 ( .A1(n22), .A2(o_data_forward_reg[373]), .Z(N235)
         );
  CKAN2D1BWP30P140LVT U1528 ( .A1(n22), .A2(o_data_forward_reg[374]), .Z(N236)
         );
  CKAN2D1BWP30P140LVT U1529 ( .A1(n20), .A2(o_data_forward_reg[325]), .Z(N320)
         );
  CKAN2D1BWP30P140LVT U1530 ( .A1(n20), .A2(o_data_forward_reg[326]), .Z(N321)
         );
  CKAN2D1BWP30P140LVT U1531 ( .A1(n20), .A2(o_data_forward_reg[327]), .Z(N322)
         );
  CKAN2D1BWP30P140LVT U1532 ( .A1(n20), .A2(o_data_forward_reg[328]), .Z(N323)
         );
  CKAN2D1BWP30P140LVT U1533 ( .A1(n20), .A2(o_data_forward_reg[329]), .Z(N324)
         );
  CKAN2D1BWP30P140LVT U1534 ( .A1(n20), .A2(o_data_forward_reg[330]), .Z(N325)
         );
  CKAN2D1BWP30P140LVT U1535 ( .A1(n20), .A2(o_data_forward_reg[331]), .Z(N326)
         );
  CKAN2D1BWP30P140LVT U1536 ( .A1(n20), .A2(o_data_forward_reg[332]), .Z(N327)
         );
  CKAN2D1BWP30P140LVT U1537 ( .A1(n20), .A2(o_data_forward_reg[333]), .Z(N328)
         );
  CKAN2D1BWP30P140LVT U1538 ( .A1(n20), .A2(o_data_forward_reg[334]), .Z(N329)
         );
  CKAN2D1BWP30P140LVT U1539 ( .A1(n20), .A2(o_data_forward_reg[335]), .Z(N330)
         );
  CKAN2D1BWP30P140LVT U1540 ( .A1(n20), .A2(o_data_forward_reg[336]), .Z(N331)
         );
  CKAN2D1BWP30P140LVT U1541 ( .A1(n20), .A2(o_data_forward_reg[337]), .Z(N332)
         );
  CKAN2D1BWP30P140LVT U1542 ( .A1(n20), .A2(o_data_forward_reg[338]), .Z(N333)
         );
  CKAN2D1BWP30P140LVT U1543 ( .A1(n20), .A2(o_data_forward_reg[339]), .Z(N334)
         );
  CKAN2D1BWP30P140LVT U1544 ( .A1(n20), .A2(o_data_forward_reg[340]), .Z(N335)
         );
  CKAN2D1BWP30P140LVT U1545 ( .A1(n20), .A2(o_data_forward_reg[341]), .Z(N336)
         );
  CKAN2D1BWP30P140LVT U1546 ( .A1(n20), .A2(o_data_forward_reg[342]), .Z(N337)
         );
  CKAN2D1BWP30P140LVT U1547 ( .A1(n20), .A2(o_data_forward_reg[343]), .Z(N338)
         );
  CKAN2D1BWP30P140LVT U1548 ( .A1(n20), .A2(o_data_forward_reg[344]), .Z(N339)
         );
  CKAN2D1BWP30P140LVT U1549 ( .A1(n20), .A2(o_data_forward_reg[345]), .Z(N340)
         );
  CKAN2D1BWP30P140LVT U1550 ( .A1(n20), .A2(o_data_forward_reg[346]), .Z(N341)
         );
  CKAN2D1BWP30P140LVT U1551 ( .A1(n20), .A2(o_data_forward_reg[347]), .Z(N342)
         );
  CKAN2D1BWP30P140LVT U1552 ( .A1(n20), .A2(o_data_forward_reg[348]), .Z(N343)
         );
  CKAN2D1BWP30P140LVT U1553 ( .A1(n20), .A2(o_data_forward_reg[349]), .Z(N344)
         );
  CKAN2D1BWP30P140LVT U1554 ( .A1(n237), .A2(o_data_forward_reg[275]), .Z(N536) );
  CKAN2D1BWP30P140LVT U1555 ( .A1(n237), .A2(o_data_forward_reg[276]), .Z(N537) );
  CKAN2D1BWP30P140LVT U1556 ( .A1(n237), .A2(o_data_forward_reg[277]), .Z(N538) );
  CKAN2D1BWP30P140LVT U1557 ( .A1(n237), .A2(o_data_forward_reg[278]), .Z(N539) );
  CKAN2D1BWP30P140LVT U1558 ( .A1(n237), .A2(o_data_forward_reg[279]), .Z(N540) );
  CKAN2D1BWP30P140LVT U1559 ( .A1(n237), .A2(o_data_forward_reg[280]), .Z(N541) );
  CKAN2D1BWP30P140LVT U1560 ( .A1(n237), .A2(o_data_forward_reg[281]), .Z(N542) );
  CKAN2D1BWP30P140LVT U1561 ( .A1(n237), .A2(o_data_forward_reg[282]), .Z(N543) );
  CKAN2D1BWP30P140LVT U1562 ( .A1(n237), .A2(o_data_forward_reg[283]), .Z(N544) );
  CKAN2D1BWP30P140LVT U1563 ( .A1(n237), .A2(o_data_forward_reg[284]), .Z(N545) );
  CKAN2D1BWP30P140LVT U1564 ( .A1(n237), .A2(o_data_forward_reg[285]), .Z(N546) );
  CKAN2D1BWP30P140LVT U1565 ( .A1(n237), .A2(o_data_forward_reg[286]), .Z(N547) );
  CKAN2D1BWP30P140LVT U1566 ( .A1(n237), .A2(o_data_forward_reg[287]), .Z(N548) );
  CKAN2D1BWP30P140LVT U1567 ( .A1(n21), .A2(o_data_forward_reg[288]), .Z(N549)
         );
  CKAN2D1BWP30P140LVT U1568 ( .A1(n21), .A2(o_data_forward_reg[289]), .Z(N550)
         );
  CKAN2D1BWP30P140LVT U1569 ( .A1(n21), .A2(o_data_forward_reg[290]), .Z(N551)
         );
  CKAN2D1BWP30P140LVT U1570 ( .A1(n21), .A2(o_data_forward_reg[291]), .Z(N552)
         );
  CKAN2D1BWP30P140LVT U1571 ( .A1(n21), .A2(o_data_forward_reg[292]), .Z(N553)
         );
  CKAN2D1BWP30P140LVT U1572 ( .A1(n21), .A2(o_data_forward_reg[293]), .Z(N554)
         );
  CKAN2D1BWP30P140LVT U1573 ( .A1(n21), .A2(o_data_forward_reg[294]), .Z(N555)
         );
  CKAN2D1BWP30P140LVT U1574 ( .A1(n21), .A2(o_data_forward_reg[295]), .Z(N556)
         );
  CKAN2D1BWP30P140LVT U1575 ( .A1(n21), .A2(o_data_forward_reg[296]), .Z(N557)
         );
  CKAN2D1BWP30P140LVT U1576 ( .A1(n21), .A2(o_data_forward_reg[297]), .Z(N558)
         );
  CKAN2D1BWP30P140LVT U1577 ( .A1(n21), .A2(o_data_forward_reg[298]), .Z(N559)
         );
  CKAN2D1BWP30P140LVT U1578 ( .A1(n21), .A2(o_data_forward_reg[299]), .Z(N560)
         );
  CKAN2D1BWP30P140LVT U1579 ( .A1(n238), .A2(o_data_forward_reg[250]), .Z(N644) );
  CKAN2D1BWP30P140LVT U1580 ( .A1(n238), .A2(o_data_forward_reg[251]), .Z(N645) );
  CKAN2D1BWP30P140LVT U1581 ( .A1(n238), .A2(o_data_forward_reg[252]), .Z(N646) );
  CKAN2D1BWP30P140LVT U1582 ( .A1(n238), .A2(o_data_forward_reg[253]), .Z(N647) );
  CKAN2D1BWP30P140LVT U1583 ( .A1(n238), .A2(o_data_forward_reg[254]), .Z(N648) );
  CKAN2D1BWP30P140LVT U1584 ( .A1(n238), .A2(o_data_forward_reg[255]), .Z(N649) );
  CKAN2D1BWP30P140LVT U1585 ( .A1(n238), .A2(o_data_forward_reg[256]), .Z(N650) );
  CKAN2D1BWP30P140LVT U1586 ( .A1(n238), .A2(o_data_forward_reg[257]), .Z(N651) );
  CKAN2D1BWP30P140LVT U1587 ( .A1(n238), .A2(o_data_forward_reg[258]), .Z(N652) );
  CKAN2D1BWP30P140LVT U1588 ( .A1(n238), .A2(o_data_forward_reg[259]), .Z(N653) );
  CKAN2D1BWP30P140LVT U1589 ( .A1(n238), .A2(o_data_forward_reg[260]), .Z(N654) );
  CKAN2D1BWP30P140LVT U1590 ( .A1(n238), .A2(o_data_forward_reg[261]), .Z(N655) );
  CKAN2D1BWP30P140LVT U1591 ( .A1(n238), .A2(o_data_forward_reg[262]), .Z(N656) );
  CKAN2D1BWP30P140LVT U1592 ( .A1(n238), .A2(o_data_forward_reg[263]), .Z(N657) );
  CKAN2D1BWP30P140LVT U1593 ( .A1(n238), .A2(o_data_forward_reg[264]), .Z(N658) );
  CKAN2D1BWP30P140LVT U1594 ( .A1(n238), .A2(o_data_forward_reg[265]), .Z(N659) );
  CKAN2D1BWP30P140LVT U1595 ( .A1(n238), .A2(o_data_forward_reg[266]), .Z(N660) );
  CKAN2D1BWP30P140LVT U1596 ( .A1(n238), .A2(o_data_forward_reg[267]), .Z(N661) );
  CKAN2D1BWP30P140LVT U1597 ( .A1(n238), .A2(o_data_forward_reg[268]), .Z(N662) );
  CKAN2D1BWP30P140LVT U1598 ( .A1(n238), .A2(o_data_forward_reg[269]), .Z(N663) );
  CKAN2D1BWP30P140LVT U1599 ( .A1(n238), .A2(o_data_forward_reg[270]), .Z(N664) );
  CKAN2D1BWP30P140LVT U1600 ( .A1(n238), .A2(o_data_forward_reg[271]), .Z(N665) );
  CKAN2D1BWP30P140LVT U1601 ( .A1(n238), .A2(o_data_forward_reg[272]), .Z(N666) );
  CKAN2D1BWP30P140LVT U1602 ( .A1(n238), .A2(o_data_forward_reg[273]), .Z(N667) );
  CKAN2D1BWP30P140LVT U1603 ( .A1(n238), .A2(o_data_forward_reg[274]), .Z(N668) );
  CKAN2D1BWP30P140LVT U1604 ( .A1(n246), .A2(o_data_forward_reg[200]), .Z(N860) );
  CKAN2D1BWP30P140LVT U1605 ( .A1(n246), .A2(o_data_forward_reg[201]), .Z(N861) );
  CKAN2D1BWP30P140LVT U1606 ( .A1(n246), .A2(o_data_forward_reg[202]), .Z(N862) );
  CKAN2D1BWP30P140LVT U1607 ( .A1(n246), .A2(o_data_forward_reg[203]), .Z(N863) );
  CKAN2D1BWP30P140LVT U1608 ( .A1(n246), .A2(o_data_forward_reg[204]), .Z(N864) );
  CKAN2D1BWP30P140LVT U1609 ( .A1(n246), .A2(o_data_forward_reg[205]), .Z(N865) );
  CKAN2D1BWP30P140LVT U1610 ( .A1(n246), .A2(o_data_forward_reg[206]), .Z(N866) );
  CKAN2D1BWP30P140LVT U1611 ( .A1(n246), .A2(o_data_forward_reg[207]), .Z(N867) );
  CKAN2D1BWP30P140LVT U1612 ( .A1(n246), .A2(o_data_forward_reg[208]), .Z(N868) );
  CKAN2D1BWP30P140LVT U1613 ( .A1(n246), .A2(o_data_forward_reg[209]), .Z(N869) );
  CKAN2D1BWP30P140LVT U1614 ( .A1(n246), .A2(o_data_forward_reg[210]), .Z(N870) );
  CKAN2D1BWP30P140LVT U1615 ( .A1(n246), .A2(o_data_forward_reg[211]), .Z(N871) );
  CKAN2D1BWP30P140LVT U1616 ( .A1(n246), .A2(o_data_forward_reg[212]), .Z(N872) );
  CKAN2D1BWP30P140LVT U1617 ( .A1(n246), .A2(o_data_forward_reg[213]), .Z(N873) );
  CKAN2D1BWP30P140LVT U1618 ( .A1(n246), .A2(o_data_forward_reg[214]), .Z(N874) );
  CKAN2D1BWP30P140LVT U1619 ( .A1(n246), .A2(o_data_forward_reg[215]), .Z(N875) );
  CKAN2D1BWP30P140LVT U1620 ( .A1(n246), .A2(o_data_forward_reg[216]), .Z(N876) );
  CKAN2D1BWP30P140LVT U1621 ( .A1(n246), .A2(o_data_forward_reg[217]), .Z(N877) );
  CKAN2D1BWP30P140LVT U1622 ( .A1(n246), .A2(o_data_forward_reg[218]), .Z(N878) );
  CKAN2D1BWP30P140LVT U1623 ( .A1(n246), .A2(o_data_forward_reg[219]), .Z(N879) );
  CKAN2D1BWP30P140LVT U1624 ( .A1(n246), .A2(o_data_forward_reg[220]), .Z(N880) );
  CKAN2D1BWP30P140LVT U1625 ( .A1(n246), .A2(o_data_forward_reg[221]), .Z(N881) );
  CKAN2D1BWP30P140LVT U1626 ( .A1(n246), .A2(o_data_forward_reg[222]), .Z(N882) );
  CKAN2D1BWP30P140LVT U1627 ( .A1(n246), .A2(o_data_forward_reg[223]), .Z(N883) );
  CKAN2D1BWP30P140LVT U1628 ( .A1(n246), .A2(o_data_forward_reg[224]), .Z(N884) );
  CKAN2D1BWP30P140LVT U1629 ( .A1(n19), .A2(o_data_forward_reg[175]), .Z(N968)
         );
  CKAN2D1BWP30P140LVT U1630 ( .A1(n19), .A2(o_data_forward_reg[176]), .Z(N969)
         );
  CKAN2D1BWP30P140LVT U1631 ( .A1(n19), .A2(o_data_forward_reg[177]), .Z(N970)
         );
  CKAN2D1BWP30P140LVT U1632 ( .A1(n19), .A2(o_data_forward_reg[178]), .Z(N971)
         );
  CKAN2D1BWP30P140LVT U1633 ( .A1(n19), .A2(o_data_forward_reg[179]), .Z(N972)
         );
  CKAN2D1BWP30P140LVT U1634 ( .A1(n19), .A2(o_data_forward_reg[180]), .Z(N973)
         );
  CKAN2D1BWP30P140LVT U1635 ( .A1(n19), .A2(o_data_forward_reg[181]), .Z(N974)
         );
  CKAN2D1BWP30P140LVT U1636 ( .A1(n19), .A2(o_data_forward_reg[182]), .Z(N975)
         );
  CKAN2D1BWP30P140LVT U1637 ( .A1(n19), .A2(o_data_forward_reg[183]), .Z(N976)
         );
  CKAN2D1BWP30P140LVT U1638 ( .A1(n19), .A2(o_data_forward_reg[184]), .Z(N977)
         );
  CKAN2D1BWP30P140LVT U1639 ( .A1(n19), .A2(o_data_forward_reg[185]), .Z(N978)
         );
  CKAN2D1BWP30P140LVT U1640 ( .A1(n19), .A2(o_data_forward_reg[186]), .Z(N979)
         );
  CKAN2D1BWP30P140LVT U1641 ( .A1(n19), .A2(o_data_forward_reg[187]), .Z(N980)
         );
  CKAN2D1BWP30P140LVT U1642 ( .A1(n19), .A2(o_data_forward_reg[188]), .Z(N981)
         );
  CKAN2D1BWP30P140LVT U1643 ( .A1(n19), .A2(o_data_forward_reg[189]), .Z(N982)
         );
  CKAN2D1BWP30P140LVT U1644 ( .A1(n19), .A2(o_data_forward_reg[190]), .Z(N983)
         );
  CKAN2D1BWP30P140LVT U1645 ( .A1(n19), .A2(o_data_forward_reg[191]), .Z(N984)
         );
  CKAN2D1BWP30P140LVT U1646 ( .A1(n19), .A2(o_data_forward_reg[192]), .Z(N985)
         );
  CKAN2D1BWP30P140LVT U1647 ( .A1(n19), .A2(o_data_forward_reg[193]), .Z(N986)
         );
  CKAN2D1BWP30P140LVT U1648 ( .A1(n19), .A2(o_data_forward_reg[194]), .Z(N987)
         );
  CKAN2D1BWP30P140LVT U1649 ( .A1(n19), .A2(o_data_forward_reg[195]), .Z(N988)
         );
  CKAN2D1BWP30P140LVT U1650 ( .A1(n19), .A2(o_data_forward_reg[196]), .Z(N989)
         );
  CKAN2D1BWP30P140LVT U1651 ( .A1(n19), .A2(o_data_forward_reg[197]), .Z(N990)
         );
  CKAN2D1BWP30P140LVT U1652 ( .A1(n19), .A2(o_data_forward_reg[198]), .Z(N991)
         );
  CKAN2D1BWP30P140LVT U1653 ( .A1(n19), .A2(o_data_forward_reg[199]), .Z(N992)
         );
  CKAN2D1BWP30P140LVT U1654 ( .A1(n240), .A2(o_data_forward_reg[150]), .Z(
        N1076) );
  CKAN2D1BWP30P140LVT U1655 ( .A1(n240), .A2(o_data_forward_reg[151]), .Z(
        N1077) );
  CKAN2D1BWP30P140LVT U1656 ( .A1(n240), .A2(o_data_forward_reg[152]), .Z(
        N1078) );
  CKAN2D1BWP30P140LVT U1657 ( .A1(n240), .A2(o_data_forward_reg[153]), .Z(
        N1079) );
  CKAN2D1BWP30P140LVT U1658 ( .A1(n240), .A2(o_data_forward_reg[154]), .Z(
        N1080) );
  CKAN2D1BWP30P140LVT U1659 ( .A1(n240), .A2(o_data_forward_reg[155]), .Z(
        N1081) );
  CKAN2D1BWP30P140LVT U1660 ( .A1(n240), .A2(o_data_forward_reg[156]), .Z(
        N1082) );
  CKAN2D1BWP30P140LVT U1661 ( .A1(n240), .A2(o_data_forward_reg[157]), .Z(
        N1083) );
  CKAN2D1BWP30P140LVT U1662 ( .A1(n240), .A2(o_data_forward_reg[158]), .Z(
        N1084) );
  CKAN2D1BWP30P140LVT U1663 ( .A1(n240), .A2(o_data_forward_reg[159]), .Z(
        N1085) );
  CKAN2D1BWP30P140LVT U1664 ( .A1(n240), .A2(o_data_forward_reg[160]), .Z(
        N1086) );
  CKAN2D1BWP30P140LVT U1665 ( .A1(n240), .A2(o_data_forward_reg[161]), .Z(
        N1087) );
  CKAN2D1BWP30P140LVT U1666 ( .A1(n240), .A2(o_data_forward_reg[162]), .Z(
        N1088) );
  CKAN2D1BWP30P140LVT U1667 ( .A1(n240), .A2(o_data_forward_reg[163]), .Z(
        N1089) );
  CKAN2D1BWP30P140LVT U1668 ( .A1(n240), .A2(o_data_forward_reg[164]), .Z(
        N1090) );
  CKAN2D1BWP30P140LVT U1669 ( .A1(n240), .A2(o_data_forward_reg[165]), .Z(
        N1091) );
  CKAN2D1BWP30P140LVT U1670 ( .A1(n240), .A2(o_data_forward_reg[166]), .Z(
        N1092) );
  CKAN2D1BWP30P140LVT U1671 ( .A1(n240), .A2(o_data_forward_reg[167]), .Z(
        N1093) );
  CKAN2D1BWP30P140LVT U1672 ( .A1(n240), .A2(o_data_forward_reg[168]), .Z(
        N1094) );
  CKAN2D1BWP30P140LVT U1673 ( .A1(n240), .A2(o_data_forward_reg[169]), .Z(
        N1095) );
  CKAN2D1BWP30P140LVT U1674 ( .A1(n240), .A2(o_data_forward_reg[170]), .Z(
        N1096) );
  CKAN2D1BWP30P140LVT U1675 ( .A1(n240), .A2(o_data_forward_reg[171]), .Z(
        N1097) );
  CKAN2D1BWP30P140LVT U1676 ( .A1(n240), .A2(o_data_forward_reg[172]), .Z(
        N1098) );
  CKAN2D1BWP30P140LVT U1677 ( .A1(n240), .A2(o_data_forward_reg[173]), .Z(
        N1099) );
  CKAN2D1BWP30P140LVT U1678 ( .A1(n240), .A2(o_data_forward_reg[174]), .Z(
        N1100) );
  CKAN2D1BWP30P140LVT U1679 ( .A1(n241), .A2(o_data_forward_reg[100]), .Z(
        N1292) );
  CKAN2D1BWP30P140LVT U1680 ( .A1(n241), .A2(o_data_forward_reg[101]), .Z(
        N1293) );
  CKAN2D1BWP30P140LVT U1681 ( .A1(n241), .A2(o_data_forward_reg[102]), .Z(
        N1294) );
  CKAN2D1BWP30P140LVT U1682 ( .A1(n241), .A2(o_data_forward_reg[103]), .Z(
        N1295) );
  CKAN2D1BWP30P140LVT U1683 ( .A1(n241), .A2(o_data_forward_reg[104]), .Z(
        N1296) );
  CKAN2D1BWP30P140LVT U1684 ( .A1(n241), .A2(o_data_forward_reg[105]), .Z(
        N1297) );
  CKAN2D1BWP30P140LVT U1685 ( .A1(n241), .A2(o_data_forward_reg[106]), .Z(
        N1298) );
  CKAN2D1BWP30P140LVT U1686 ( .A1(n241), .A2(o_data_forward_reg[107]), .Z(
        N1299) );
  CKAN2D1BWP30P140LVT U1687 ( .A1(n241), .A2(o_data_forward_reg[108]), .Z(
        N1300) );
  CKAN2D1BWP30P140LVT U1688 ( .A1(n241), .A2(o_data_forward_reg[109]), .Z(
        N1301) );
  CKAN2D1BWP30P140LVT U1689 ( .A1(n241), .A2(o_data_forward_reg[110]), .Z(
        N1302) );
  CKAN2D1BWP30P140LVT U1690 ( .A1(n241), .A2(o_data_forward_reg[111]), .Z(
        N1303) );
  CKAN2D1BWP30P140LVT U1691 ( .A1(n241), .A2(o_data_forward_reg[112]), .Z(
        N1304) );
  CKAN2D1BWP30P140LVT U1692 ( .A1(n241), .A2(o_data_forward_reg[113]), .Z(
        N1305) );
  CKAN2D1BWP30P140LVT U1693 ( .A1(n241), .A2(o_data_forward_reg[114]), .Z(
        N1306) );
  CKAN2D1BWP30P140LVT U1694 ( .A1(n241), .A2(o_data_forward_reg[115]), .Z(
        N1307) );
  CKAN2D1BWP30P140LVT U1695 ( .A1(n241), .A2(o_data_forward_reg[116]), .Z(
        N1308) );
  CKAN2D1BWP30P140LVT U1696 ( .A1(n241), .A2(o_data_forward_reg[117]), .Z(
        N1309) );
  CKAN2D1BWP30P140LVT U1697 ( .A1(n241), .A2(o_data_forward_reg[118]), .Z(
        N1310) );
  CKAN2D1BWP30P140LVT U1698 ( .A1(n241), .A2(o_data_forward_reg[119]), .Z(
        N1311) );
  CKAN2D1BWP30P140LVT U1699 ( .A1(n241), .A2(o_data_forward_reg[120]), .Z(
        N1312) );
  CKAN2D1BWP30P140LVT U1700 ( .A1(n241), .A2(o_data_forward_reg[121]), .Z(
        N1313) );
  CKAN2D1BWP30P140LVT U1701 ( .A1(n241), .A2(o_data_forward_reg[122]), .Z(
        N1314) );
  CKAN2D1BWP30P140LVT U1702 ( .A1(n241), .A2(o_data_forward_reg[123]), .Z(
        N1315) );
  CKAN2D1BWP30P140LVT U1703 ( .A1(n241), .A2(o_data_forward_reg[124]), .Z(
        N1316) );
  CKAN2D1BWP30P140LVT U1704 ( .A1(n242), .A2(o_data_forward_reg[50]), .Z(N1508) );
  CKAN2D1BWP30P140LVT U1705 ( .A1(n242), .A2(o_data_forward_reg[51]), .Z(N1509) );
  CKAN2D1BWP30P140LVT U1706 ( .A1(n242), .A2(o_data_forward_reg[52]), .Z(N1510) );
  CKAN2D1BWP30P140LVT U1707 ( .A1(n242), .A2(o_data_forward_reg[53]), .Z(N1511) );
  CKAN2D1BWP30P140LVT U1708 ( .A1(n242), .A2(o_data_forward_reg[54]), .Z(N1512) );
  CKAN2D1BWP30P140LVT U1709 ( .A1(n242), .A2(o_data_forward_reg[55]), .Z(N1513) );
  CKAN2D1BWP30P140LVT U1710 ( .A1(n242), .A2(o_data_forward_reg[56]), .Z(N1514) );
  CKAN2D1BWP30P140LVT U1711 ( .A1(n242), .A2(o_data_forward_reg[57]), .Z(N1515) );
  CKAN2D1BWP30P140LVT U1712 ( .A1(n242), .A2(o_data_forward_reg[58]), .Z(N1516) );
  CKAN2D1BWP30P140LVT U1713 ( .A1(n242), .A2(o_data_forward_reg[59]), .Z(N1517) );
  CKAN2D1BWP30P140LVT U1714 ( .A1(n242), .A2(o_data_forward_reg[60]), .Z(N1518) );
  CKAN2D1BWP30P140LVT U1715 ( .A1(n242), .A2(o_data_forward_reg[61]), .Z(N1519) );
  CKAN2D1BWP30P140LVT U1716 ( .A1(n242), .A2(o_data_forward_reg[62]), .Z(N1520) );
  CKAN2D1BWP30P140LVT U1717 ( .A1(n242), .A2(o_data_forward_reg[63]), .Z(N1521) );
  CKAN2D1BWP30P140LVT U1718 ( .A1(n242), .A2(o_data_forward_reg[64]), .Z(N1522) );
  CKAN2D1BWP30P140LVT U1719 ( .A1(n242), .A2(o_data_forward_reg[65]), .Z(N1523) );
  CKAN2D1BWP30P140LVT U1720 ( .A1(n242), .A2(o_data_forward_reg[66]), .Z(N1524) );
  CKAN2D1BWP30P140LVT U1721 ( .A1(n242), .A2(o_data_forward_reg[67]), .Z(N1525) );
  CKAN2D1BWP30P140LVT U1722 ( .A1(n242), .A2(o_data_forward_reg[68]), .Z(N1526) );
  CKAN2D1BWP30P140LVT U1723 ( .A1(n242), .A2(o_data_forward_reg[69]), .Z(N1527) );
  CKAN2D1BWP30P140LVT U1724 ( .A1(n242), .A2(o_data_forward_reg[70]), .Z(N1528) );
  CKAN2D1BWP30P140LVT U1725 ( .A1(n242), .A2(o_data_forward_reg[71]), .Z(N1529) );
  CKAN2D1BWP30P140LVT U1726 ( .A1(n242), .A2(o_data_forward_reg[72]), .Z(N1530) );
  CKAN2D1BWP30P140LVT U1727 ( .A1(n242), .A2(o_data_forward_reg[73]), .Z(N1531) );
  CKAN2D1BWP30P140LVT U1728 ( .A1(n242), .A2(o_data_forward_reg[74]), .Z(N1532) );
  CKAN2D1BWP30P140LVT U1729 ( .A1(n243), .A2(o_data_forward_reg[25]), .Z(N1616) );
  CKAN2D1BWP30P140LVT U1730 ( .A1(n243), .A2(o_data_forward_reg[26]), .Z(N1617) );
  CKAN2D1BWP30P140LVT U1731 ( .A1(n243), .A2(o_data_forward_reg[27]), .Z(N1618) );
  CKAN2D1BWP30P140LVT U1732 ( .A1(n243), .A2(o_data_forward_reg[28]), .Z(N1619) );
  CKAN2D1BWP30P140LVT U1733 ( .A1(n243), .A2(o_data_forward_reg[29]), .Z(N1620) );
  CKAN2D1BWP30P140LVT U1734 ( .A1(n243), .A2(o_data_forward_reg[30]), .Z(N1621) );
  CKAN2D1BWP30P140LVT U1735 ( .A1(n243), .A2(o_data_forward_reg[31]), .Z(N1622) );
  CKAN2D1BWP30P140LVT U1736 ( .A1(n243), .A2(o_data_forward_reg[32]), .Z(N1623) );
  CKAN2D1BWP30P140LVT U1737 ( .A1(n243), .A2(o_data_forward_reg[33]), .Z(N1624) );
  CKAN2D1BWP30P140LVT U1738 ( .A1(n243), .A2(o_data_forward_reg[34]), .Z(N1625) );
  CKAN2D1BWP30P140LVT U1739 ( .A1(n243), .A2(o_data_forward_reg[35]), .Z(N1626) );
  CKAN2D1BWP30P140LVT U1740 ( .A1(n243), .A2(o_data_forward_reg[36]), .Z(N1627) );
  CKAN2D1BWP30P140LVT U1741 ( .A1(n243), .A2(o_data_forward_reg[37]), .Z(N1628) );
  CKAN2D1BWP30P140LVT U1742 ( .A1(n243), .A2(o_data_forward_reg[38]), .Z(N1629) );
  CKAN2D1BWP30P140LVT U1743 ( .A1(n243), .A2(o_data_forward_reg[39]), .Z(N1630) );
  CKAN2D1BWP30P140LVT U1744 ( .A1(n243), .A2(o_data_forward_reg[40]), .Z(N1631) );
  CKAN2D1BWP30P140LVT U1745 ( .A1(n243), .A2(o_data_forward_reg[41]), .Z(N1632) );
  CKAN2D1BWP30P140LVT U1746 ( .A1(n243), .A2(o_data_forward_reg[42]), .Z(N1633) );
  CKAN2D1BWP30P140LVT U1747 ( .A1(n243), .A2(o_data_forward_reg[43]), .Z(N1634) );
  CKAN2D1BWP30P140LVT U1748 ( .A1(n243), .A2(o_data_forward_reg[44]), .Z(N1635) );
  CKAN2D1BWP30P140LVT U1749 ( .A1(n243), .A2(o_data_forward_reg[45]), .Z(N1636) );
  CKAN2D1BWP30P140LVT U1750 ( .A1(n243), .A2(o_data_forward_reg[46]), .Z(N1637) );
  CKAN2D1BWP30P140LVT U1751 ( .A1(n243), .A2(o_data_forward_reg[47]), .Z(N1638) );
  CKAN2D1BWP30P140LVT U1752 ( .A1(n243), .A2(o_data_forward_reg[48]), .Z(N1639) );
  CKAN2D1BWP30P140LVT U1753 ( .A1(n243), .A2(o_data_forward_reg[49]), .Z(N1640) );
  INR2D1BWP30P140LVT U1754 ( .A1(o_cmd_forward_reg[4]), .B1(n53), .ZN(N1667)
         );
  INR2D1BWP30P140LVT U1755 ( .A1(o_cmd_forward_reg[7]), .B1(n53), .ZN(N1670)
         );
  INR2D1BWP30P140LVT U1756 ( .A1(o_valid_forward_reg[13]), .B1(n18), .ZN(N1666) );
  INR2D1BWP30P140LVT U1757 ( .A1(o_cmd_forward_reg[9]), .B1(n53), .ZN(N1560)
         );
  INR2D1BWP30P140LVT U1758 ( .A1(o_cmd_forward_reg[10]), .B1(n18), .ZN(N1561)
         );
  INR2D1BWP30P140LVT U1759 ( .A1(o_valid_forward_reg[12]), .B1(n18), .ZN(N1558) );
  INR2D1BWP30P140LVT U1760 ( .A1(o_cmd_forward_reg[12]), .B1(n18), .ZN(N1451)
         );
  INR2D1BWP30P140LVT U1761 ( .A1(o_valid_forward_reg[11]), .B1(n53), .ZN(N1450) );
  INR2D1BWP30P140LVT U1762 ( .A1(o_cmd_forward_reg[18]), .B1(n18), .ZN(N1345)
         );
  INR2D1BWP30P140LVT U1763 ( .A1(o_cmd_forward_reg[19]), .B1(n53), .ZN(N1346)
         );
  INR2D1BWP30P140LVT U1764 ( .A1(o_valid_forward_reg[10]), .B1(n18), .ZN(N1342) );
  INR2D1BWP30P140LVT U1765 ( .A1(o_cmd_forward_reg[20]), .B1(n18), .ZN(N1235)
         );
  INR2D1BWP30P140LVT U1766 ( .A1(o_valid_forward_reg[9]), .B1(n18), .ZN(N1234)
         );
  INR2D1BWP30P140LVT U1767 ( .A1(o_cmd_forward_reg[25]), .B1(n18), .ZN(N1128)
         );
  INR2D1BWP30P140LVT U1768 ( .A1(o_cmd_forward_reg[27]), .B1(n53), .ZN(N1130)
         );
  INR2D1BWP30P140LVT U1769 ( .A1(o_valid_forward_reg[8]), .B1(n18), .ZN(N1126)
         );
  INR2D1BWP30P140LVT U1770 ( .A1(o_cmd_forward_reg[28]), .B1(n18), .ZN(N1019)
         );
  INR2D1BWP30P140LVT U1771 ( .A1(o_valid_forward_reg[7]), .B1(n18), .ZN(N1018)
         );
  INR2D1BWP30P140LVT U1772 ( .A1(o_cmd_forward_reg[35]), .B1(n18), .ZN(N914)
         );
  INR2D1BWP30P140LVT U1773 ( .A1(o_valid_forward_reg[6]), .B1(n18), .ZN(N910)
         );
  INR2D1BWP30P140LVT U1774 ( .A1(o_cmd_forward_reg[36]), .B1(n18), .ZN(N803)
         );
  INR2D1BWP30P140LVT U1775 ( .A1(o_cmd_forward_reg[38]), .B1(n53), .ZN(N805)
         );
  INR2D1BWP30P140LVT U1776 ( .A1(o_cmd_forward_reg[41]), .B1(n18), .ZN(N696)
         );
  INR2D1BWP30P140LVT U1777 ( .A1(o_cmd_forward_reg[42]), .B1(n53), .ZN(N697)
         );
  INR2D1BWP30P140LVT U1778 ( .A1(o_valid_forward_reg[4]), .B1(n53), .ZN(N694)
         );
  INR2D1BWP30P140LVT U1779 ( .A1(o_cmd_forward_reg[44]), .B1(n18), .ZN(N587)
         );
  INR2D1BWP30P140LVT U1780 ( .A1(o_valid_forward_reg[3]), .B1(n18), .ZN(N586)
         );
  INR2D1BWP30P140LVT U1781 ( .A1(o_cmd_forward_reg[50]), .B1(n53), .ZN(N481)
         );
  INR2D1BWP30P140LVT U1782 ( .A1(o_valid_forward_reg[2]), .B1(n53), .ZN(N478)
         );
  INR2D1BWP30P140LVT U1783 ( .A1(o_cmd_forward_reg[52]), .B1(n53), .ZN(N371)
         );
  INR2D1BWP30P140LVT U1784 ( .A1(o_valid_forward_reg[1]), .B1(n18), .ZN(N370)
         );
  INR2D1BWP30P140LVT U1785 ( .A1(o_cmd_forward_reg[57]), .B1(n18), .ZN(N264)
         );
  INR2D1BWP30P140LVT U1786 ( .A1(o_valid_forward_reg[0]), .B1(n18), .ZN(N262)
         );
  INR2D1BWP30P140LVT U1787 ( .A1(i_cmd[0]), .B1(n18), .ZN(N155) );
endmodule

